// Verilog netlist created by TD v5.0.38657
// Fri Feb 25 00:18:31 2022

`timescale 1ns / 1ps
module SOC_TOP  // ../RTL/soc_top/soc_top.v(5)
  (
  i_clk,
  i_io_rx,
  i_rstn,
  o_io_tx
  );

  input i_clk;  // ../RTL/soc_top/soc_top.v(6)
  input i_io_rx;  // ../RTL/soc_top/soc_top.v(9)
  input i_rstn;  // ../RTL/soc_top/soc_top.v(7)
  output o_io_tx;  // ../RTL/soc_top/soc_top.v(10)

  wire [31:0] periph_addr;  // ../RTL/soc_top/soc_top.v(40)
  wire [31:0] periph_rdata;  // ../RTL/soc_top/soc_top.v(44)
  wire [31:0] periph_wdata;  // ../RTL/soc_top/soc_top.v(43)
  wire [31:0] \u_PERIPH_TOP/timer_ribs_rdata ;  // ../RTL/periph/periph_top.v(65)
  wire [31:0] \u_PERIPH_TOP/u_SLAVE_SEL/n14 ;
  wire [1:0] \u_PERIPH_TOP/u_SLAVE_SEL/sel_tag ;  // ../RTL/core/rib.v(78)
  wire [7:0] \u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id ;  // ../RTL/core/rib.v(113)
  wire [63:0] \u_PERIPH_TOP/u_TIMER2RIB/n12 ;
  wire [63:0] \u_PERIPH_TOP/u_TIMER2RIB/n13 ;
  wire [63:0] \u_PERIPH_TOP/u_TIMER2RIB/n14 ;
  wire [63:0] \u_PERIPH_TOP/u_TIMER2RIB/n18 ;
  wire [31:0] \u_PERIPH_TOP/u_TIMER2RIB/n2 ;
  wire [31:0] \u_PERIPH_TOP/u_TIMER2RIB/n4 ;
  wire [31:0] \u_PERIPH_TOP/u_TIMER2RIB/n5 ;
  wire [63:0] \u_PERIPH_TOP/u_TIMER2RIB/timer_cnt ;  // ../RTL/periph/timer2rib.v(30)
  wire [31:0] \u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl ;  // ../RTL/periph/timer2rib.v(29)
  wire [31:0] \u_PERIPH_TOP/u_USART2RIB/n2 ;
  wire [31:0] \u_PERIPH_TOP/u_USART2RIB/n5 ;
  wire [31:0] \u_PERIPH_TOP/u_USART2RIB/n6 ;
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/rx_data ;  // ../RTL/periph/usart2rib.v(34)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/tx_buffer ;  // ../RTL/periph/usart2rib.v(30)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 ;  // al_ip/usart_gate.v(45)
  wire [5:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 ;  // al_ip/usart_gate.v(46)
  wire [5:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 ;  // al_ip/usart_gate.v(49)
  wire [5:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 ;  // al_ip/usart_gate.v(48)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 ;  // al_ip/usart_gate.v(47)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 ;  // al_ip/usart_gate.v(50)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 ;  // al_ip/usart_gate.v(52)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 ;  // al_ip/usart_gate.v(51)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 ;  // al_ip/usart_gate.v(55)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 ;  // al_ip/usart_gate.v(56)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 ;  // al_ip/usart_gate.v(57)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 ;  // al_ip/usart_gate.v(60)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 ;  // al_ip/usart_gate.v(59)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 ;  // al_ip/usart_gate.v(58)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 ;  // al_ip/usart_gate.v(61)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 ;  // al_ip/usart_gate.v(67)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A68B0 ;  // al_ip/usart_gate.v(69)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A7020 ;  // al_ip/usart_gate.v(68)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 ;  // al_ip/usart_gate.v(70)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 ;  // al_ip/usart_gate.v(71)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 ;  // al_ip/usart_gate.v(72)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 ;  // al_ip/usart_gate.v(73)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 ;  // al_ip/usart_gate.v(74)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 ;  // al_ip/usart_gate.v(75)
  wire [31:0] \u_PERIPH_TOP/usart_rib_rdata ;  // ../RTL/periph/periph_top.v(35)
  wire [4:0] \u_internal_reset/synch_regs_q ;  // ../RTL/core/reset.v(13)
  wire clk_84mhz;  // ../RTL/soc_top/soc_top.v(16)
  wire extlock;  // ../RTL/soc_top/soc_top.v(15)
  wire n0;
  wire n1;
  wire \periph_addr[10]_neg ;
  wire \periph_addr[11]_neg ;
  wire \periph_addr[12]_neg ;
  wire \periph_addr[13]_neg ;
  wire \periph_addr[14]_neg ;
  wire \periph_addr[15]_neg ;
  wire \periph_addr[4]_neg ;
  wire \periph_addr[5]_neg ;
  wire \periph_addr[6]_neg ;
  wire \periph_addr[7]_neg ;
  wire \periph_addr[8]_neg ;
  wire \periph_addr[9]_neg ;
  wire periph_req;  // ../RTL/soc_top/soc_top.v(45)
  wire periph_wrcs;  // ../RTL/soc_top/soc_top.v(41)
  wire reset;  // ../RTL/soc_top/soc_top.v(31)
  wire \u_PERIPH_TOP/timer_ribs_req ;  // ../RTL/periph/periph_top.v(66)
  wire \u_PERIPH_TOP/timer_ribs_rsp ;  // ../RTL/periph/periph_top.v(68)
  wire \u_PERIPH_TOP/u_SLAVE_SEL/default_cs ;  // ../RTL/core/rib.v(112)
  wire \u_PERIPH_TOP/u_SLAVE_SEL/default_cs_neg ;
  wire \u_PERIPH_TOP/u_SLAVE_SEL/handshake_rdy ;  // ../RTL/core/rib.v(114)
  wire \u_PERIPH_TOP/u_SLAVE_SEL/handshake_rdy_last ;  // ../RTL/core/rib.v(117)
  wire \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_SLAVE_SEL/n0 ;
  wire \u_PERIPH_TOP/u_SLAVE_SEL/n1 ;
  wire \u_PERIPH_TOP/u_SLAVE_SEL/n2 ;
  wire \u_PERIPH_TOP/u_SLAVE_SEL/n3 ;
  wire \u_PERIPH_TOP/u_SLAVE_SEL/n5 ;
  wire \u_PERIPH_TOP/u_SLAVE_SEL/n6 ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/mux3_b0_sel_is_3_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/mux4_b0_sel_is_3_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/n6 ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/n7 ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/n8 ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel0_b0_sel_is_3_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_0_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_10_sel_is_0_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_1_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_2_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_3_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_4_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_5_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_6_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_7_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_8_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_9_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b10_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b11_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b12_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b13_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b14_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b15_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b16_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b17_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b18_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b19_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b1_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b20_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b21_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b22_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b23_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b24_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b25_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b26_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b27_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b28_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b29_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b2_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b30_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b31_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b3_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b4_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b5_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b6_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b7_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b8_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b9_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/mux1_b0_sel_is_3_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/mux2_b0_sel_is_3_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/n13 ;
  wire \u_PERIPH_TOP/u_USART2RIB/n16 ;
  wire \u_PERIPH_TOP/u_USART2RIB/rx_err ;  // ../RTL/periph/usart2rib.v(35)
  wire \u_PERIPH_TOP/u_USART2RIB/rx_vld ;  // ../RTL/periph/usart2rib.v(33)
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b0_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b1_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b2_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b3_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b4_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b5_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b6_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b7_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/tx_en ;  // ../RTL/periph/usart2rib.v(37)
  wire \u_PERIPH_TOP/u_USART2RIB/tx_rdy ;  // ../RTL/periph/usart2rib.v(36)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533120 ;  // al_ip/usart_gate.v(160)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533280 ;  // al_ip/usart_gate.v(157)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533330 ;  // al_ip/usart_gate.v(163)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5335F0 ;  // al_ip/usart_gate.v(158)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533B70 ;  // al_ip/usart_gate.v(161)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533CD0 ;  // al_ip/usart_gate.v(165)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533D80 ;  // al_ip/usart_gate.v(167)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533EE0 ;  // al_ip/usart_gate.v(168)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534040 ;  // al_ip/usart_gate.v(171)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5340F0 ;  // al_ip/usart_gate.v(173)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5341A0 ;  // al_ip/usart_gate.v(180)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534250 ;  // al_ip/usart_gate.v(181)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534300 ;  // al_ip/usart_gate.v(182)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534460 ;  // al_ip/usart_gate.v(169)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534510 ;  // al_ip/usart_gate.v(164)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5345C0 ;  // al_ip/usart_gate.v(176)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534880 ;  // al_ip/usart_gate.v(162)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534A90 ;  // al_ip/usart_gate.v(174)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534B40 ;  // al_ip/usart_gate.v(175)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534BF0 ;  // al_ip/usart_gate.v(177)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534D50 ;  // al_ip/usart_gate.v(178)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535380 ;  // al_ip/usart_gate.v(166)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535430 ;  // al_ip/usart_gate.v(170)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535590 ;  // al_ip/usart_gate.v(172)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535640 ;  // al_ip/usart_gate.v(179)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535BC0 ;  // al_ip/usart_gate.v(159)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A340 ;  // al_ip/usart_gate.v(200)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A550 ;  // al_ip/usart_gate.v(199)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A550340 ;  // al_ip/usart_gate.v(53)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ;  // al_ip/usart_gate.v(213)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ;  // al_ip/usart_gate.v(214)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E290 ;  // al_ip/usart_gate.v(143)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E3F0 ;  // al_ip/usart_gate.v(147)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E4A0 ;  // al_ip/usart_gate.v(144)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E600 ;  // al_ip/usart_gate.v(148)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E8C0 ;  // al_ip/usart_gate.v(149)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82ECE0 ;  // al_ip/usart_gate.v(142)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FB50 ;  // al_ip/usart_gate.v(146)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FCB0 ;  // al_ip/usart_gate.v(150)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FEC0 ;  // al_ip/usart_gate.v(151)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830020 ;  // al_ip/usart_gate.v(145)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830390 ;  // al_ip/usart_gate.v(152)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830B20 ;  // al_ip/usart_gate.v(141)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830C80 ;  // al_ip/usart_gate.v(156)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ;  // al_ip/usart_gate.v(154)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A831C50 ;  // al_ip/usart_gate.v(153)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A832AC0 ;  // al_ip/usart_gate.v(183)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A832EE0 ;  // al_ip/usart_gate.v(155)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ;  // al_ip/usart_gate.v(184)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ;  // al_ip/usart_gate.v(187)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C9110 ;  // al_ip/usart_gate.v(186)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C93D0 ;  // al_ip/usart_gate.v(188)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C95E0 ;  // al_ip/usart_gate.v(185)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB2C0 ;  // al_ip/usart_gate.v(189)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB420 ;  // al_ip/usart_gate.v(190)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB6E0 ;  // al_ip/usart_gate.v(192)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB790 ;  // al_ip/usart_gate.v(196)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB840 ;  // al_ip/usart_gate.v(191)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CBF20 ;  // al_ip/usart_gate.v(197)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CC810 ;  // al_ip/usart_gate.v(198)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCA20 ;  // al_ip/usart_gate.v(195)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCD90 ;  // al_ip/usart_gate.v(193)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD470 ;  // al_ip/usart_gate.v(194)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD890 ;  // al_ip/usart_gate.v(201)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ;  // al_ip/usart_gate.v(202)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2010 ;  // al_ip/usart_gate.v(204)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2F30 ;  // al_ip/usart_gate.v(203)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D3FB0 ;  // al_ip/usart_gate.v(211)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4320 ;  // al_ip/usart_gate.v(205)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4480 ;  // al_ip/usart_gate.v(209)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4C10 ;  // al_ip/usart_gate.v(207)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D50E0 ;  // al_ip/usart_gate.v(206)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5A80 ;  // al_ip/usart_gate.v(210)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5B30 ;  // al_ip/usart_gate.v(212)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5BE0 ;  // al_ip/usart_gate.v(208)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5BBF0 ;  // al_ip/usart_gate.v(54)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5D780 ;  // al_ip/usart_gate.v(62)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5F070 ;  // al_ip/usart_gate.v(63)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA60730 ;  // al_ip/usart_gate.v(64)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA63600 ;  // al_ip/usart_gate.v(65)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9D8A0 ;  // al_ip/usart_gate.v(139)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9D950 ;  // al_ip/usart_gate.v(80)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DA00 ;  // al_ip/usart_gate.v(135)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DAB0 ;  // al_ip/usart_gate.v(118)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DB60 ;  // al_ip/usart_gate.v(119)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DC10 ;  // al_ip/usart_gate.v(126)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DCC0 ;  // al_ip/usart_gate.v(136)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ;  // al_ip/usart_gate.v(121)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DE20 ;  // al_ip/usart_gate.v(76)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DED0 ;  // al_ip/usart_gate.v(78)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DF80 ;  // al_ip/usart_gate.v(92)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ;  // al_ip/usart_gate.v(96)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E0E0 ;  // al_ip/usart_gate.v(97)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E190 ;  // al_ip/usart_gate.v(101)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E240 ;  // al_ip/usart_gate.v(87)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ;  // al_ip/usart_gate.v(127)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E500 ;  // al_ip/usart_gate.v(116)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ;  // al_ip/usart_gate.v(128)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E710 ;  // al_ip/usart_gate.v(138)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E7C0 ;  // al_ip/usart_gate.v(91)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ;  // al_ip/usart_gate.v(79)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E920 ;  // al_ip/usart_gate.v(93)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E9D0 ;  // al_ip/usart_gate.v(103)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EA80 ;  // al_ip/usart_gate.v(102)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EB30 ;  // al_ip/usart_gate.v(104)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EBE0 ;  // al_ip/usart_gate.v(105)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EC90 ;  // al_ip/usart_gate.v(106)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EDF0 ;  // al_ip/usart_gate.v(140)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EEA0 ;  // al_ip/usart_gate.v(107)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EF50 ;  // al_ip/usart_gate.v(108)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F000 ;  // al_ip/usart_gate.v(89)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ;  // al_ip/usart_gate.v(134)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F160 ;  // al_ip/usart_gate.v(125)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F210 ;  // al_ip/usart_gate.v(122)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ;  // al_ip/usart_gate.v(77)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F370 ;  // al_ip/usart_gate.v(81)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F420 ;  // al_ip/usart_gate.v(123)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F4D0 ;  // al_ip/usart_gate.v(84)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F580 ;  // al_ip/usart_gate.v(131)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F630 ;  // al_ip/usart_gate.v(85)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F6E0 ;  // al_ip/usart_gate.v(94)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F790 ;  // al_ip/usart_gate.v(98)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ;  // al_ip/usart_gate.v(124)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F8F0 ;  // al_ip/usart_gate.v(82)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F9A0 ;  // al_ip/usart_gate.v(88)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FA50 ;  // al_ip/usart_gate.v(83)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FB00 ;  // al_ip/usart_gate.v(90)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ;  // al_ip/usart_gate.v(117)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FC60 ;  // al_ip/usart_gate.v(95)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FD10 ;  // al_ip/usart_gate.v(99)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FDC0 ;  // al_ip/usart_gate.v(100)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FF20 ;  // al_ip/usart_gate.v(132)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FFD0 ;  // al_ip/usart_gate.v(129)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0080 ;  // al_ip/usart_gate.v(133)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA01E0 ;  // al_ip/usart_gate.v(137)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0290 ;  // al_ip/usart_gate.v(130)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0340 ;  // al_ip/usart_gate.v(86)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA03F0 ;  // al_ip/usart_gate.v(120)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0760 ;  // al_ip/usart_gate.v(115)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0A20 ;  // al_ip/usart_gate.v(114)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1100 ;  // al_ip/usart_gate.v(110)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1940 ;  // al_ip/usart_gate.v(112)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1AA0 ;  // al_ip/usart_gate.v(109)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1F70 ;  // al_ip/usart_gate.v(113)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA22E0 ;  // al_ip/usart_gate.v(111)
  wire \u_PERIPH_TOP/usart_rib_req ;  // ../RTL/periph/periph_top.v(36)
  wire \u_PERIPH_TOP/usart_rib_rsp ;  // ../RTL/periph/periph_top.v(38)
  wire \u_pll/clk0_buf ;  // al_ip/pll.v(32)

  not \periph_addr[10]_inv  (\periph_addr[10]_neg , periph_addr[10]);
  not \periph_addr[11]_inv  (\periph_addr[11]_neg , periph_addr[11]);
  not \periph_addr[12]_inv  (\periph_addr[12]_neg , periph_addr[12]);
  not \periph_addr[13]_inv  (\periph_addr[13]_neg , periph_addr[13]);
  not \periph_addr[14]_inv  (\periph_addr[14]_neg , periph_addr[14]);
  not \periph_addr[15]_inv  (\periph_addr[15]_neg , periph_addr[15]);
  not \periph_addr[4]_inv  (\periph_addr[4]_neg , periph_addr[4]);
  not \periph_addr[5]_inv  (\periph_addr[5]_neg , periph_addr[5]);
  not \periph_addr[6]_inv  (\periph_addr[6]_neg , periph_addr[6]);
  not \periph_addr[7]_inv  (\periph_addr[7]_neg , periph_addr[7]);
  not \periph_addr[8]_inv  (\periph_addr[8]_neg , periph_addr[8]);
  not \periph_addr[9]_inv  (\periph_addr[9]_neg , periph_addr[9]);
  not u1 (n0, i_rstn);  // ../RTL/soc_top/soc_top.v(19)
  and u2 (n1, i_rstn, extlock);  // ../RTL/soc_top/soc_top.v(34)
  CORE_TOP u_CORE_TOP (
    .i_clk(clk_84mhz),
    .i_ribp_gnt(\u_PERIPH_TOP/u_SLAVE_SEL/n0 ),
    .i_ribp_rdata(periph_rdata),
    .i_ribp_rsp(\u_PERIPH_TOP/u_SLAVE_SEL/n1 ),
    .i_ribx_gnt(1'b0),
    .i_ribx_rdata(32'b00000000000000000000000000000000),
    .i_ribx_rsp(1'b0),
    .i_rstn(reset),
    .o_ribp_addr({periph_addr[31:24],open_n0,open_n1,open_n2,open_n3,open_n4,open_n5,open_n6,open_n7,periph_addr[15:2],open_n8,open_n9}),
    .o_ribp_req(periph_req),
    .o_ribp_wdata(periph_wdata),
    .o_ribp_wrcs(periph_wrcs));  // ../RTL/soc_top/soc_top.v(51)
  not \u_PERIPH_TOP/u_SLAVE_SEL/default_cs_inv  (\u_PERIPH_TOP/u_SLAVE_SEL/default_cs_neg , \u_PERIPH_TOP/u_SLAVE_SEL/default_cs );
  AL_DFF_X \u_PERIPH_TOP/u_SLAVE_SEL/default_cs_reg  (
    .ar(1'b0),
    .as(~reset),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/n3 ),
    .en(\u_PERIPH_TOP/u_SLAVE_SEL/n6 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ));  // ../RTL/core/rib.v(121)
  eq_w8 \u_PERIPH_TOP/u_SLAVE_SEL/eq0  (
    .i0(periph_addr[31:24]),
    .i1(8'b11110001),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [0]));  // ../RTL/core/rib.v(83)
  eq_w8 \u_PERIPH_TOP/u_SLAVE_SEL/eq1  (
    .i0(periph_addr[31:24]),
    .i1(8'b11110010),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]));  // ../RTL/core/rib.v(83)
  AL_DFF_X \u_PERIPH_TOP/u_SLAVE_SEL/handshake_rdy_last_reg  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/handshake_rdy ),
    .en(\u_PERIPH_TOP/u_SLAVE_SEL/n6 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_SLAVE_SEL/handshake_rdy_last ));  // ../RTL/core/rib.v(121)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux2_b0  (
    .i0(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [0]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux2_b1  (
    .i0(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [1]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux2_b2  (
    .i0(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [2]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux2_b3  (
    .i0(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [3]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux2_b4  (
    .i0(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [4]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux2_b5  (
    .i0(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [5]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux2_b6  (
    .i0(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [6]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux2_b7  (
    .i0(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [7]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b0  (
    .i0(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [0]),
    .i1(1'b0),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .o(periph_rdata[0]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b1  (
    .i0(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [1]),
    .i1(1'b0),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .o(periph_rdata[1]));  // ../RTL/core/rib.v(146)
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[10]));
  and \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2  (\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o , \u_PERIPH_TOP/u_SLAVE_SEL/default_cs_neg , \u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]);
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b11  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[11]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b12  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[12]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b13  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[13]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b14  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[14]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b15  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[15]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b16  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[16]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b17  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[17]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b18  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[18]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b19  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[19]));
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b2  (
    .i0(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [2]),
    .i1(1'b0),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .o(periph_rdata[2]));  // ../RTL/core/rib.v(146)
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b20  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[20]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b21  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[21]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b22  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[22]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b23  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[23]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b24  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[24]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b25  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[25]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b26  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[26]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b27  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[27]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b28  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[28]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b29  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[29]));
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b3  (
    .i0(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [3]),
    .i1(1'b0),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .o(periph_rdata[3]));  // ../RTL/core/rib.v(146)
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b30  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[30]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b31  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[31]));
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b4  (
    .i0(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [4]),
    .i1(1'b0),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .o(periph_rdata[4]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b5  (
    .i0(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [5]),
    .i1(1'b0),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .o(periph_rdata[5]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b6  (
    .i0(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [6]),
    .i1(1'b0),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .o(periph_rdata[6]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b7  (
    .i0(\u_PERIPH_TOP/u_SLAVE_SEL/n14 [7]),
    .i1(1'b0),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .o(periph_rdata[7]));  // ../RTL/core/rib.v(146)
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b8  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[8]));
  AL_MUX \u_PERIPH_TOP/u_SLAVE_SEL/mux3_b9  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .sel(\u_PERIPH_TOP/u_SLAVE_SEL/mux3_b10_sel_is_2_o ),
    .o(periph_rdata[9]));
  AL_DFF_X \u_PERIPH_TOP/u_SLAVE_SEL/reg0_b0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .en(\u_PERIPH_TOP/u_SLAVE_SEL/n6 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]));  // ../RTL/core/rib.v(121)
  and \u_PERIPH_TOP/u_SLAVE_SEL/u14  (\u_PERIPH_TOP/usart_rib_req , periph_req, \u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [0]);  // ../RTL/core/rib.v(90)
  and \u_PERIPH_TOP/u_SLAVE_SEL/u159  (\u_PERIPH_TOP/timer_ribs_req , periph_req, \u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]);  // ../RTL/core/rib.v(90)
  or \u_PERIPH_TOP/u_SLAVE_SEL/u16  (\u_PERIPH_TOP/u_SLAVE_SEL/n0 , \u_PERIPH_TOP/usart_rib_req , \u_PERIPH_TOP/timer_ribs_req );  // ../RTL/core/rib.v(95)
  or \u_PERIPH_TOP/u_SLAVE_SEL/u18  (\u_PERIPH_TOP/u_SLAVE_SEL/n1 , \u_PERIPH_TOP/usart_rib_rsp , \u_PERIPH_TOP/timer_ribs_rsp );  // ../RTL/core/rib.v(97)
  not \u_PERIPH_TOP/u_SLAVE_SEL/u23  (\u_PERIPH_TOP/u_SLAVE_SEL/n3 , \u_PERIPH_TOP/u_SLAVE_SEL/n2 );  // ../RTL/core/rib.v(105)
  and \u_PERIPH_TOP/u_SLAVE_SEL/u25  (\u_PERIPH_TOP/u_SLAVE_SEL/handshake_rdy , periph_req, \u_PERIPH_TOP/u_SLAVE_SEL/n0 );  // ../RTL/core/rib.v(114)
  not \u_PERIPH_TOP/u_SLAVE_SEL/u31  (\u_PERIPH_TOP/u_SLAVE_SEL/n5 , \u_PERIPH_TOP/u_SLAVE_SEL/handshake_rdy_last );  // ../RTL/core/rib.v(128)
  or \u_PERIPH_TOP/u_SLAVE_SEL/u32  (\u_PERIPH_TOP/u_SLAVE_SEL/n6 , \u_PERIPH_TOP/u_SLAVE_SEL/n1 , \u_PERIPH_TOP/u_SLAVE_SEL/n5 );  // ../RTL/core/rib.v(128)
  or \u_PERIPH_TOP/u_SLAVE_SEL/u33  (\u_PERIPH_TOP/u_SLAVE_SEL/n2 , \u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [0], \u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]);  // ../RTL/core/rib.v(105)
  add_pu64_pu64_o64 \u_PERIPH_TOP/u_TIMER2RIB/add0  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt ),
    .i1(64'b0000000000000000000000000000000000000000000000000000000000000001),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n13 ));  // ../RTL/periph/timer2rib.v(73)
  eq_w16 \u_PERIPH_TOP/u_TIMER2RIB/eq0  (
    .i0({periph_addr[15:2],2'b00}),
    .i1(16'b0000000000000000),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n6 ));  // ../RTL/periph/timer2rib.v(42)
  eq_w16 \u_PERIPH_TOP/u_TIMER2RIB/eq1  (
    .i0({periph_addr[15:2],2'b00}),
    .i1(16'b0000000000000100),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n7 ));  // ../RTL/periph/timer2rib.v(52)
  eq_w16 \u_PERIPH_TOP/u_TIMER2RIB/eq2  (
    .i0({periph_addr[15:2],2'b00}),
    .i1(16'b0000000000001000),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n8 ));  // ../RTL/periph/timer2rib.v(60)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b0  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [0]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [0]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [0]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b1  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [1]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [1]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [1]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b10  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [10]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [10]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [10]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b11  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [11]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [11]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [11]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b12  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [12]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [12]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [12]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b13  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [13]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [13]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [13]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b14  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [14]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [14]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [14]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b15  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [15]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [15]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [15]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b16  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [16]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [16]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [16]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b17  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [17]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [17]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [17]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b18  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [18]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [18]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [18]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b19  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [19]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [19]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [19]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b2  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [2]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [2]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [2]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b20  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [20]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [20]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [20]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b21  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [21]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [21]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [21]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b22  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [22]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [22]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [22]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b23  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [23]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [23]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [23]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b24  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [24]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [24]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [24]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b25  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [25]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [25]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [25]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b26  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [26]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [26]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [26]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b27  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [27]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [27]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [27]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b28  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [28]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [28]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [28]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b29  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [29]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [29]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [29]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b3  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [3]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [3]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [3]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b30  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [30]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [30]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [30]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b31  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [31]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [31]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [31]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b32  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [32]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [32]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [32]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b33  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [33]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [33]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [33]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b34  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [34]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [34]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [34]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b35  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [35]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [35]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [35]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b36  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [36]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [36]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [36]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b37  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [37]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [37]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [37]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b38  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [38]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [38]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [38]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b39  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [39]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [39]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [39]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b4  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [4]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [4]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [4]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b40  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [40]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [40]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [40]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b41  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [41]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [41]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [41]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b42  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [42]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [42]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [42]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b43  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [43]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [43]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [43]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b44  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [44]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [44]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [44]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b45  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [45]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [45]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [45]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b46  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [46]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [46]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [46]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b47  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [47]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [47]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [47]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b48  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [48]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [48]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [48]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b49  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [49]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [49]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [49]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b5  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [5]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [5]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [5]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b50  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [50]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [50]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [50]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b51  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [51]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [51]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [51]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b52  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [52]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [52]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [52]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b53  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [53]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [53]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [53]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b54  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [54]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [54]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [54]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b55  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [55]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [55]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [55]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b56  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [56]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [56]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [56]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b57  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [57]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [57]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [57]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b58  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [58]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [58]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [58]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b59  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [59]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [59]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [59]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b6  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [6]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [6]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [6]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b60  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [60]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [60]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [60]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b61  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [61]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [61]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [61]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b62  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [62]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [62]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [62]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b63  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [63]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [63]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [63]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b7  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [7]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [7]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [7]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b8  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [8]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [8]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [8]));  // ../RTL/periph/timer2rib.v(72)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux2_b9  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [9]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n13 [9]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [9]));  // ../RTL/periph/timer2rib.v(72)
  and \u_PERIPH_TOP/u_TIMER2RIB/mux3_b0_sel_is_3  (\u_PERIPH_TOP/u_TIMER2RIB/mux3_b0_sel_is_3_o , \u_PERIPH_TOP/timer_ribs_req , \u_PERIPH_TOP/u_TIMER2RIB/sel0_b0_sel_is_3_o );
  and \u_PERIPH_TOP/u_TIMER2RIB/mux4_b0_sel_is_3  (\u_PERIPH_TOP/u_TIMER2RIB/mux4_b0_sel_is_3_o , \u_PERIPH_TOP/timer_ribs_req , \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_0_sel_is_2_o );
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b0  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [0]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [0]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [0]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b1  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [1]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [1]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [1]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b10  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [10]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [10]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [10]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b11  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [11]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [11]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [11]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b12  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [12]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [12]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [12]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b13  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [13]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [13]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [13]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b14  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [14]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [14]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [14]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b15  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [15]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [15]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [15]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b16  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [16]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [16]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [16]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b17  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [17]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [17]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [17]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b18  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [18]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [18]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [18]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b19  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [19]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [19]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [19]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b2  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [2]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [2]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [2]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b20  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [20]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [20]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [20]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b21  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [21]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [21]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [21]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b22  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [22]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [22]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [22]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b23  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [23]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [23]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [23]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b24  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [24]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [24]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [24]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b25  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [25]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [25]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [25]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b26  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [26]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [26]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [26]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b27  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [27]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [27]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [27]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b28  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [28]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [28]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [28]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b29  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [29]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [29]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [29]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b3  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [3]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [3]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [3]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b30  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [30]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [30]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [30]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b31  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [31]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [31]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [31]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b32  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [32]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [32]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [32]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b33  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [33]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [33]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [33]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b34  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [34]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [34]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [34]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b35  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [35]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [35]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [35]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b36  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [36]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [36]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [36]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b37  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [37]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [37]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [37]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b38  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [38]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [38]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [38]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b39  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [39]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [39]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [39]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b4  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [4]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [4]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [4]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b40  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [40]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [40]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [40]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b41  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [41]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [41]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [41]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b42  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [42]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [42]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [42]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b43  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [43]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [43]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [43]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b44  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [44]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [44]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [44]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b45  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [45]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [45]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [45]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b46  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [46]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [46]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [46]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b47  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [47]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [47]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [47]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b48  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [48]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [48]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [48]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b49  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [49]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [49]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [49]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b5  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [5]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [5]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [5]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b50  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [50]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [50]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [50]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b51  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [51]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [51]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [51]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b52  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [52]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [52]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [52]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b53  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [53]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [53]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [53]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b54  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [54]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [54]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [54]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b55  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [55]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [55]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [55]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b56  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [56]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [56]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [56]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b57  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [57]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [57]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [57]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b58  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [58]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [58]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [58]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b59  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [59]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [59]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [59]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b6  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [6]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [6]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [6]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b60  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [60]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [60]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [60]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b61  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [61]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [61]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [61]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b62  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [62]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [62]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [62]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b63  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [63]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [63]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [63]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b7  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [7]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [7]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [7]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b8  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [8]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [8]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [8]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux5_b9  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n14 [9]),
    .i1(\u_PERIPH_TOP/u_TIMER2RIB/n12 [9]),
    .sel(\u_PERIPH_TOP/timer_ribs_req ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [9]));  // ../RTL/periph/timer2rib.v(39)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b0  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [32]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [0]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b1  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [33]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [1]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b10  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [42]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [10]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b11  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [43]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [11]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b12  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [44]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [12]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b13  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [45]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [13]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b14  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [46]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [14]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b15  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [47]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [15]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b16  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [48]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [16]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b17  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [49]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [17]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b18  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [50]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [18]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b19  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [51]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [19]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b2  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [34]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [2]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b20  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [52]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [20]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b21  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [53]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [21]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b22  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [54]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [22]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b23  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [55]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [23]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b24  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [56]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [24]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b25  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [57]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [25]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b26  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [58]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [26]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b27  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [59]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [27]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b28  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [60]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [28]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b29  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [61]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [29]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b3  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [35]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [3]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b30  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [62]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [30]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b31  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [63]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [31]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b32  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [0]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [0]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b33  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [1]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [1]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b34  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [2]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [2]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b35  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [3]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [3]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b36  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [4]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [4]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b37  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [5]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [5]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b38  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [6]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [6]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b39  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [7]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [7]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b4  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [36]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [4]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b40  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [8]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [8]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b41  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [9]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [9]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b42  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [10]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [10]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b43  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [11]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [11]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b44  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [12]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [12]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b45  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [13]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [13]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b46  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [14]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [14]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b47  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [15]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [15]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b48  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [16]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [16]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b49  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [17]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [17]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b5  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [37]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [5]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b50  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [18]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [18]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b51  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [19]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [19]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b52  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [20]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [20]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b53  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [21]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [21]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b54  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [22]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [22]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b55  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [23]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [23]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b56  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [24]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [24]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b57  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [25]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [25]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b58  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [26]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [26]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b59  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [27]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [27]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b6  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [38]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [6]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b60  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [28]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [28]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b61  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [29]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [29]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b62  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [30]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [30]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b63  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [31]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n4 [31]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b64  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [0]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b65  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [1]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b66  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [2]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b67  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [3]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b68  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [4]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b69  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [5]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b7  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [39]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [7]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b70  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [6]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b71  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [7]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b72  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [8]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b73  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [9]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b74  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [10]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b75  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [11]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b76  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [12]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b77  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [13]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b78  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [14]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b79  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [15]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b8  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [40]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [8]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b80  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [16]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b81  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [17]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b82  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [18]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b83  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [19]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b84  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [20]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b85  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [21]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b86  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [22]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b87  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [23]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b88  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [24]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b89  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [25]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b9  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [41]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n5 [9]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b90  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [26]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b91  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [27]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b92  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [28]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b93  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [29]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b94  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [30]));  // ../RTL/periph/timer2rib.v(43)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_TIMER2RIB/mux6_b95  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n2 [31]));  // ../RTL/periph/timer2rib.v(43)
  and \u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2  (\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o , reset, \u_PERIPH_TOP/u_TIMER2RIB/mux4_b0_sel_is_3_o );
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/o_ribs_rsp_reg  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/timer_ribs_req ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rsp ));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [0]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b1  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [1]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b10  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [10]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b11  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [11]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b12  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [12]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b13  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [13]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b14  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [14]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b15  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [15]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b16  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [16]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b17  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [17]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b18  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [18]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b19  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [19]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b2  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [2]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b20  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [20]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b21  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [21]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b22  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [22]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b23  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [23]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b24  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [24]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b25  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [25]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b26  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [26]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b27  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [27]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b28  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [28]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b29  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [29]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b3  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [3]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b30  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [30]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b31  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [31]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b32  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [32]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b33  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [33]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b34  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [34]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b35  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [35]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b36  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [36]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b37  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [37]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b38  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [38]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b39  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [39]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b4  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [4]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b40  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [40]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b41  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [41]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b42  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [42]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b43  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [43]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b44  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [44]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b45  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [45]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b46  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [46]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b47  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [47]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b48  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [48]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b49  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [49]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b5  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [5]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b50  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [50]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b51  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [51]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b52  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [52]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b53  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [53]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b54  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [54]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b55  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [55]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b56  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [56]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b57  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [57]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b58  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [58]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b59  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [59]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b6  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [6]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b60  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [60]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b61  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [61]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b62  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [62]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [62]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b63  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [63]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [63]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b7  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [7]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b8  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [8]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg0_b9  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [9]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [0]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b1_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [1]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b10_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [10]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b11_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [11]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b12_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [12]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b13_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [13]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b14_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [14]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b15_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [15]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b16_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [16]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b17_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [17]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b18_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [18]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b19_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [19]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b2_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [2]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b20_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [20]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b21_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [21]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b22_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [22]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b23_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [23]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b24_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [24]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b25_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [25]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b26_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [26]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b27_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [27]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b28_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [28]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b29_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [29]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b3_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [3]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b30_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [30]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b31_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [31]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b4_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [4]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b5_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [5]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b6_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [6]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b7_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [7]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b8_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [8]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg1_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b9_var_o ),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [9]));  // ../RTL/periph/timer2rib.v(34)
  AL_DFF_X \u_PERIPH_TOP/u_TIMER2RIB/reg2_b0  (
    .ar(1'b0),
    .as(~reset),
    .clk(clk_84mhz),
    .d(periph_wdata[0]),
    .en(\u_PERIPH_TOP/u_TIMER2RIB/mux3_b0_sel_is_3_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]));  // ../RTL/periph/timer2rib.v(34)
  and \u_PERIPH_TOP/u_TIMER2RIB/sel0_b0_sel_is_3  (\u_PERIPH_TOP/u_TIMER2RIB/sel0_b0_sel_is_3_o , \u_PERIPH_TOP/u_TIMER2RIB/n6 , periph_wrcs);
  and \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_0_sel_is_2  (\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_0_sel_is_2_o , \periph_addr[15]_neg , \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_1_sel_is_2_o );
  and \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_10_sel_is_0  (\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_10_sel_is_0_o , \periph_addr[5]_neg , \periph_addr[4]_neg );
  and \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_1_sel_is_2  (\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_1_sel_is_2_o , \periph_addr[14]_neg , \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_2_sel_is_2_o );
  and \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_2_sel_is_2  (\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_2_sel_is_2_o , \periph_addr[13]_neg , \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_3_sel_is_2_o );
  and \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_3_sel_is_2  (\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_3_sel_is_2_o , \periph_addr[12]_neg , \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_4_sel_is_2_o );
  and \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_4_sel_is_2  (\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_4_sel_is_2_o , \periph_addr[11]_neg , \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_5_sel_is_2_o );
  and \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_5_sel_is_2  (\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_5_sel_is_2_o , \periph_addr[10]_neg , \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_6_sel_is_2_o );
  and \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_6_sel_is_2  (\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_6_sel_is_2_o , \periph_addr[9]_neg , \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_7_sel_is_2_o );
  and \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_7_sel_is_2  (\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_7_sel_is_2_o , \periph_addr[8]_neg , \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_8_sel_is_2_o );
  and \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_8_sel_is_2  (\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_8_sel_is_2_o , \periph_addr[7]_neg , \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_9_sel_is_2_o );
  and \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_9_sel_is_2  (\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_9_sel_is_2_o , \periph_addr[6]_neg , \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_10_sel_is_0_o );
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [0]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [0]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [0]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b10_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [10]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [10]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [10]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b10_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b11_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [11]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [11]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [11]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b11_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b12_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [12]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [12]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [12]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b12_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b13_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [13]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [13]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [13]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b13_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b14_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [14]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [14]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [14]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b14_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b15_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [15]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [15]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [15]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b15_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b16_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [16]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [16]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [16]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b16_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b17_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [17]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [17]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [17]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b17_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b18_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [18]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [18]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [18]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b18_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b19_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [19]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [19]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [19]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b19_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b1_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [1]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [1]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [1]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b1_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b20_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [20]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [20]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [20]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b20_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b21_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [21]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [21]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [21]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b21_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b22_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [22]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [22]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [22]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b22_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b23_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [23]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [23]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [23]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b23_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b24_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [24]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [24]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [24]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b24_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b25_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [25]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [25]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [25]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b25_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b26_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [26]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [26]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [26]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b26_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b27_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [27]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [27]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [27]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b27_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b28_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [28]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [28]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [28]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b28_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b29_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [29]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [29]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [29]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b29_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b2_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [2]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [2]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [2]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b2_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b30_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [30]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [30]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [30]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b30_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b31_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [31]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [31]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [31]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b31_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b3_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [3]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [3]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [3]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b3_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b4_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [4]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [4]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [4]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b4_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b5_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [5]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [5]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [5]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b5_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b6_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [6]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [6]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [6]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b6_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b7_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [7]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [7]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [7]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b7_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b8_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [8]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [8]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [8]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b8_var_o ));  // ../RTL/periph/timer2rib.v(41)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_TIMER2RIB/sel1_b9_var  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/n2 [9]),
    .i1(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .i10(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .i11(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .i12(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .i13(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .i14(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .i15(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .i2(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .i3(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .i4(\u_PERIPH_TOP/u_TIMER2RIB/n4 [9]),
    .i5(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .i6(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .i7(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .i8(\u_PERIPH_TOP/u_TIMER2RIB/n5 [9]),
    .i9(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b9_var_o ));  // ../RTL/periph/timer2rib.v(41)
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b0  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [0]),
    .i1(periph_wdata[0]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [0]));
  and \u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3  (\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o , \u_PERIPH_TOP/u_TIMER2RIB/n7 , periph_wrcs);
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b1  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [1]),
    .i1(periph_wdata[1]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [1]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b10  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [10]),
    .i1(periph_wdata[10]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [10]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b11  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [11]),
    .i1(periph_wdata[11]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [11]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b12  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [12]),
    .i1(periph_wdata[12]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [12]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b13  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [13]),
    .i1(periph_wdata[13]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [13]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b14  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [14]),
    .i1(periph_wdata[14]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [14]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b15  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [15]),
    .i1(periph_wdata[15]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [15]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b16  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [16]),
    .i1(periph_wdata[16]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [16]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b17  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [17]),
    .i1(periph_wdata[17]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [17]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b18  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [18]),
    .i1(periph_wdata[18]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [18]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b19  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [19]),
    .i1(periph_wdata[19]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [19]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b2  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [2]),
    .i1(periph_wdata[2]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [2]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b20  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [20]),
    .i1(periph_wdata[20]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [20]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b21  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [21]),
    .i1(periph_wdata[21]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [21]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b22  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [22]),
    .i1(periph_wdata[22]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [22]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b23  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [23]),
    .i1(periph_wdata[23]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [23]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b24  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [24]),
    .i1(periph_wdata[24]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [24]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b25  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [25]),
    .i1(periph_wdata[25]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [25]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b26  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [26]),
    .i1(periph_wdata[26]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [26]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b27  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [27]),
    .i1(periph_wdata[27]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [27]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b28  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [28]),
    .i1(periph_wdata[28]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [28]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b29  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [29]),
    .i1(periph_wdata[29]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [29]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b3  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [3]),
    .i1(periph_wdata[3]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [3]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b30  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [30]),
    .i1(periph_wdata[30]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [30]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b31  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [31]),
    .i1(periph_wdata[31]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [31]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b32  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [32]),
    .i1(periph_wdata[0]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [32]));
  and \u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3  (\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o , \u_PERIPH_TOP/u_TIMER2RIB/n8 , periph_wrcs);
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b33  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [33]),
    .i1(periph_wdata[1]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [33]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b34  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [34]),
    .i1(periph_wdata[2]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [34]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b35  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [35]),
    .i1(periph_wdata[3]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [35]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b36  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [36]),
    .i1(periph_wdata[4]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [36]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b37  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [37]),
    .i1(periph_wdata[5]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [37]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b38  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [38]),
    .i1(periph_wdata[6]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [38]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b39  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [39]),
    .i1(periph_wdata[7]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [39]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b4  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [4]),
    .i1(periph_wdata[4]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [4]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b40  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [40]),
    .i1(periph_wdata[8]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [40]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b41  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [41]),
    .i1(periph_wdata[9]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [41]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b42  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [42]),
    .i1(periph_wdata[10]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [42]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b43  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [43]),
    .i1(periph_wdata[11]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [43]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b44  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [44]),
    .i1(periph_wdata[12]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [44]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b45  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [45]),
    .i1(periph_wdata[13]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [45]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b46  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [46]),
    .i1(periph_wdata[14]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [46]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b47  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [47]),
    .i1(periph_wdata[15]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [47]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b48  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [48]),
    .i1(periph_wdata[16]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [48]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b49  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [49]),
    .i1(periph_wdata[17]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [49]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b5  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [5]),
    .i1(periph_wdata[5]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [5]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b50  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [50]),
    .i1(periph_wdata[18]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [50]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b51  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [51]),
    .i1(periph_wdata[19]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [51]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b52  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [52]),
    .i1(periph_wdata[20]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [52]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b53  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [53]),
    .i1(periph_wdata[21]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [53]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b54  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [54]),
    .i1(periph_wdata[22]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [54]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b55  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [55]),
    .i1(periph_wdata[23]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [55]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b56  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [56]),
    .i1(periph_wdata[24]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [56]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b57  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [57]),
    .i1(periph_wdata[25]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [57]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b58  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [58]),
    .i1(periph_wdata[26]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [58]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b59  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [59]),
    .i1(periph_wdata[27]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [59]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b6  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [6]),
    .i1(periph_wdata[6]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [6]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b60  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [60]),
    .i1(periph_wdata[28]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [60]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b61  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [61]),
    .i1(periph_wdata[29]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [61]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b62  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [62]),
    .i1(periph_wdata[30]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [62]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b63  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [63]),
    .i1(periph_wdata[31]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [63]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b7  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [7]),
    .i1(periph_wdata[7]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [7]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b8  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [8]),
    .i1(periph_wdata[8]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [8]));
  AL_MUX \u_PERIPH_TOP/u_TIMER2RIB/sel2_b9  (
    .i0(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [9]),
    .i1(periph_wdata[9]),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [9]));
  and \u_PERIPH_TOP/u_USART2RIB/mux1_b0_sel_is_3  (\u_PERIPH_TOP/u_USART2RIB/mux1_b0_sel_is_3_o , \u_PERIPH_TOP/usart_rib_req , \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_0_sel_is_2_o );
  and \u_PERIPH_TOP/u_USART2RIB/mux2_b0_sel_is_3  (\u_PERIPH_TOP/u_USART2RIB/mux2_b0_sel_is_3_o , \u_PERIPH_TOP/usart_rib_req , \u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o );
  and \u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2  (\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o , reset, \u_PERIPH_TOP/u_USART2RIB/mux1_b0_sel_is_3_o );
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b0  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/rx_data [0]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n6 [0]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b1  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/rx_data [1]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n6 [1]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b2  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/rx_data [2]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n6 [2]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b3  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/rx_data [3]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n6 [3]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b32  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [0]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n5 [0]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b33  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [1]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n5 [1]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b34  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [2]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n5 [2]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b35  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [3]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n5 [3]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b36  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [4]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n5 [4]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b37  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [5]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n5 [5]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b38  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [6]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n5 [6]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b39  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [7]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n5 [7]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b4  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/rx_data [4]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n6 [4]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b5  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/rx_data [5]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n6 [5]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b6  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/rx_data [6]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n6 [6]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b64  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/tx_rdy ),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n2 [0]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b65  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/rx_vld ),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n2 [1]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b66  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/rx_err ),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n2 [2]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b67  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n2 [3]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b68  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n2 [4]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b69  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n2 [5]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b7  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/rx_data [7]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n6 [7]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b70  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n2 [6]));  // ../RTL/periph/usart2rib.v(56)
  binary_mux_s1_w1 \u_PERIPH_TOP/u_USART2RIB/mux4_b71  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .sel(periph_wrcs),
    .o(\u_PERIPH_TOP/u_USART2RIB/n2 [7]));  // ../RTL/periph/usart2rib.v(56)
  and \u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2  (\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o , reset, \u_PERIPH_TOP/u_USART2RIB/mux2_b0_sel_is_3_o );
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/o_ribs_rsp_reg  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/usart_rib_req ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/usart_rib_rsp ));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg0_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b0_var_o ),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/usart_rib_rdata [0]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg0_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b1_var_o ),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/usart_rib_rdata [1]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg0_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b2_var_o ),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/usart_rib_rdata [2]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg0_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b3_var_o ),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/usart_rib_rdata [3]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg0_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b4_var_o ),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/usart_rib_rdata [4]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg0_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b5_var_o ),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/usart_rib_rdata [5]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg0_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b6_var_o ),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/usart_rib_rdata [6]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg0_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b7_var_o ),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/usart_rib_rdata [7]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg1_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(periph_wdata[0]),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [0]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg1_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(periph_wdata[1]),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [1]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg1_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(periph_wdata[2]),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [2]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg1_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(periph_wdata[3]),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [3]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg1_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(periph_wdata[4]),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [4]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg1_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(periph_wdata[5]),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [5]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg1_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(periph_wdata[6]),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [6]));  // ../RTL/periph/usart2rib.v(48)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/reg1_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(periph_wdata[7]),
    .en(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [7]));  // ../RTL/periph/usart2rib.v(48)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_USART2RIB/sel0_b0_var  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/n2 [0]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i10(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i11(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i12(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i13(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i14(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i15(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i2(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i3(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i4(\u_PERIPH_TOP/u_USART2RIB/n5 [0]),
    .i5(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i6(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i7(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .i8(\u_PERIPH_TOP/u_USART2RIB/n6 [0]),
    .i9(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b0_var_o ));  // ../RTL/periph/usart2rib.v(54)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_USART2RIB/sel0_b1_var  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/n2 [1]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i10(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i11(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i12(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i13(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i14(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i15(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i2(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i3(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i4(\u_PERIPH_TOP/u_USART2RIB/n5 [1]),
    .i5(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i6(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i7(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .i8(\u_PERIPH_TOP/u_USART2RIB/n6 [1]),
    .i9(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b1_var_o ));  // ../RTL/periph/usart2rib.v(54)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_USART2RIB/sel0_b2_var  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/n2 [2]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i10(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i11(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i12(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i13(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i14(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i15(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i2(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i3(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i4(\u_PERIPH_TOP/u_USART2RIB/n5 [2]),
    .i5(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i6(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i7(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .i8(\u_PERIPH_TOP/u_USART2RIB/n6 [2]),
    .i9(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b2_var_o ));  // ../RTL/periph/usart2rib.v(54)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_USART2RIB/sel0_b3_var  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/n2 [3]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i10(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i11(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i12(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i13(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i14(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i15(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i2(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i3(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i4(\u_PERIPH_TOP/u_USART2RIB/n5 [3]),
    .i5(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i6(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i7(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .i8(\u_PERIPH_TOP/u_USART2RIB/n6 [3]),
    .i9(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b3_var_o ));  // ../RTL/periph/usart2rib.v(54)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_USART2RIB/sel0_b4_var  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/n2 [4]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i10(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i11(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i12(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i13(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i14(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i15(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i2(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i3(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i4(\u_PERIPH_TOP/u_USART2RIB/n5 [4]),
    .i5(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i6(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i7(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .i8(\u_PERIPH_TOP/u_USART2RIB/n6 [4]),
    .i9(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b4_var_o ));  // ../RTL/periph/usart2rib.v(54)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_USART2RIB/sel0_b5_var  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/n2 [5]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i10(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i11(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i12(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i13(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i14(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i15(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i2(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i3(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i4(\u_PERIPH_TOP/u_USART2RIB/n5 [5]),
    .i5(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i6(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i7(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .i8(\u_PERIPH_TOP/u_USART2RIB/n6 [5]),
    .i9(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b5_var_o ));  // ../RTL/periph/usart2rib.v(54)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_USART2RIB/sel0_b6_var  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/n2 [6]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i10(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i11(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i12(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i13(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i14(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i15(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i2(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i3(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i4(\u_PERIPH_TOP/u_USART2RIB/n5 [6]),
    .i5(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i6(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i7(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .i8(\u_PERIPH_TOP/u_USART2RIB/n6 [6]),
    .i9(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b6_var_o ));  // ../RTL/periph/usart2rib.v(54)
  binary_mux_s4_w1 \u_PERIPH_TOP/u_USART2RIB/sel0_b7_var  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/n2 [7]),
    .i1(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i10(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i11(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i12(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i13(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i14(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i15(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i2(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i3(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i4(\u_PERIPH_TOP/u_USART2RIB/n5 [7]),
    .i5(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i6(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i7(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .i8(\u_PERIPH_TOP/u_USART2RIB/n6 [7]),
    .i9(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .sel({periph_addr[3:2],2'b00}),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b7_var_o ));  // ../RTL/periph/usart2rib.v(54)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/tx_en_reg  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/n16 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_en ));  // ../RTL/periph/usart2rib.v(48)
  AL_MUX \u_PERIPH_TOP/u_USART2RIB/u13  (
    .i0(\u_PERIPH_TOP/u_USART2RIB/tx_en ),
    .i1(1'b1),
    .sel(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b0_sel_is_3_o ),
    .o(\u_PERIPH_TOP/u_USART2RIB/n13 ));
  AL_MUX \u_PERIPH_TOP/u_USART2RIB/u14  (
    .i0(1'b0),
    .i1(\u_PERIPH_TOP/u_USART2RIB/n13 ),
    .sel(\u_PERIPH_TOP/usart_rib_req ),
    .o(\u_PERIPH_TOP/u_USART2RIB/n16 ));  // ../RTL/periph/usart2rib.v(53)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A78C4C0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB840 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCD90 ));  // al_ip/usart_gate.v(1818)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A78F160  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A832EE0 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ));  // al_ip/usart_gate.v(1468)
  AL_DFF_0 \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A78F490  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ));  // al_ip/usart_gate.v(1477)
  AL_DFF_0 \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A826290  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [3]));  // al_ip/usart_gate.v(1594)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8268F0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 [2]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [2]));  // al_ip/usart_gate.v(1558)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A826F50  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 [1]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [1]));  // al_ip/usart_gate.v(1549)
  AL_DFF_0 \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A827060  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [5]));  // al_ip/usart_gate.v(1612)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A827390  (
    .ar(1'b0),
    .as(~reset),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D50E0 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_io_tx));  // al_ip/usart_gate.v(2358)
  AL_DFF_0 \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A827D20  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [4]));  // al_ip/usart_gate.v(1603)
  AL_DFF_0 \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A827F40  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [1]));  // al_ip/usart_gate.v(1576)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A828380  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 [0]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [0]));  // al_ip/usart_gate.v(1540)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8285A0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5BE0 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4480 ));  // al_ip/usart_gate.v(2367)
  AL_DFF_0 \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8298C0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [0]));  // al_ip/usart_gate.v(1567)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A829F20  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2010 ),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD890 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5A80 ));  // al_ip/usart_gate.v(2376)
  AL_DFF_0 \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82A360  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [2]));  // al_ip/usart_gate.v(1585)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82CBC0  (
    .ar(1'b0),
    .as(~reset),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4320 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_rdy ));  // al_ip/usart_gate.v(2385)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82CCD0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D3FB0 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5B30 ));  // al_ip/usart_gate.v(2394)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A876BF0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [3]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [3]));  // al_ip/usart_gate.v(1854)
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'b0000010010001100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A877360  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0A20 ));  // al_ip/usart_gate.v(785)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A877470  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [2]));  // al_ip/usart_gate.v(1881)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A877580  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [5]));  // al_ip/usart_gate.v(1971)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~(~C*~B)))"),
    .INIT(32'b10101010101010101010101000000010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8779C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1100 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA22E0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1940 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [3]));  // al_ip/usart_gate.v(765)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A877AD0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [3]));  // al_ip/usart_gate.v(1953)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A877F10  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 [1]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]));  // al_ip/usart_gate.v(1908)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878130  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [1]));  // al_ip/usart_gate.v(1935)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878240  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [3]));  // al_ip/usart_gate.v(1890)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878350  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [6]));  // al_ip/usart_gate.v(1980)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878460  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [1]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [0]));  // al_ip/usart_gate.v(1998)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878570  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [0]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [0]));  // al_ip/usart_gate.v(1827)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878680  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 [2]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]));  // al_ip/usart_gate.v(1917)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878790  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [2]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [1]));  // al_ip/usart_gate.v(2007)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878AC0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [1]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [1]));  // al_ip/usart_gate.v(1836)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878BD0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 [0]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]));  // al_ip/usart_gate.v(1899)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111000010111111011100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878CE0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1F70 ));  // al_ip/usart_gate.v(775)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878DF0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [7]));  // al_ip/usart_gate.v(1989)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878F00  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [3]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [2]));  // al_ip/usart_gate.v(2016)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879120  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [1]));  // al_ip/usart_gate.v(1872)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'b0000001000000111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879450  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [2]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0760 ));  // al_ip/usart_gate.v(794)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~(~C*~B)))"),
    .INIT(32'b10101010101010101010101000000010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879560  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1F70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0A20 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0760 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [2]));  // al_ip/usart_gate.v(803)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879670  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0]));  // al_ip/usart_gate.v(1926)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879890  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2]));  // al_ip/usart_gate.v(1944)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879BC0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [0]));  // al_ip/usart_gate.v(1863)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879CD0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [4]));  // al_ip/usart_gate.v(1962)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879DE0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [4]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [3]));  // al_ip/usart_gate.v(2025)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879EF0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [5]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [4]));  // al_ip/usart_gate.v(2034)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'b0000001000000111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87A000  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [3]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1940 ));  // al_ip/usart_gate.v(756)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87A110  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [2]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [2]));  // al_ip/usart_gate.v(1845)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87A220  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [6]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [5]));  // al_ip/usart_gate.v(2043)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87A440  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCA20 ),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [7]));  // al_ip/usart_gate.v(2061)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87A550  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [7]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [6]));  // al_ip/usart_gate.v(2052)
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'b01))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87B650  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 [0]));  // al_ip/usart_gate.v(813)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87D850  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [0]),
    .b(1'b1),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830B20 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82ECE0 ,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [0]}));  // al_ip/usart_gate.v(1423)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87D960  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [1]),
    .b(1'b0),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82ECE0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E290 ,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [1]}));  // al_ip/usart_gate.v(1430)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87EC80  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [5]),
    .b(1'b0),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FB50 ),
    .o({open_n86,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [5]}));  // al_ip/usart_gate.v(1458)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87EEA0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [2]),
    .b(1'b0),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E290 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E4A0 ,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [2]}));  // al_ip/usart_gate.v(1437)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F610  (
    .a(1'b1),
    .b(1'b0),
    .c(1'b0),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E3F0 ,open_n87}));  // al_ip/usart_gate.v(1530)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F720  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [4]),
    .b(1'b0),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830020 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FB50 ,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [4]}));  // al_ip/usart_gate.v(1451)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F940  (
    .a(1'b0),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E3F0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E600 ,open_n88}));  // al_ip/usart_gate.v(1488)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87FD80  (
    .a(1'b0),
    .b(1'b0),
    .c(1'b0),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830B20 ,open_n89}));  // al_ip/usart_gate.v(1465)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87FFA0  (
    .a(1'b0),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E600 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E8C0 ,open_n90}));  // al_ip/usart_gate.v(1495)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8800B0  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [2]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E8C0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FCB0 ,open_n91}));  // al_ip/usart_gate.v(1502)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8801C0  (
    .a(1'b0),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [4]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FEC0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830390 ,open_n92}));  // al_ip/usart_gate.v(1516)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A880930  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [3]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FCB0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FEC0 ,open_n93}));  // al_ip/usart_gate.v(1509)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A880B50  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [5]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830390 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A831C50 ,open_n94}));  // al_ip/usart_gate.v(1523)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8814E0  (
    .a(1'b0),
    .b(1'b1),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A831C50 ),
    .o({open_n95,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 }));  // al_ip/usart_gate.v(1535)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A881A30  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4C10 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D3FB0 ));  // al_ip/usart_gate.v(2403)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A881C50  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [3]),
    .b(1'b0),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E4A0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830020 ,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [3]}));  // al_ip/usart_gate.v(1444)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9326A0  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533D80 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533EE0 ,open_n96}));  // al_ip/usart_gate.v(1698)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9327B0  (
    .ar(1'b0),
    .as(~reset),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [3]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A832AC0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCA20 ));  // al_ip/usart_gate.v(2088)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9328C0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [7]));  // al_ip/usart_gate.v(2349)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A932BF0  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533CD0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535380 ,open_n97}));  // al_ip/usart_gate.v(1684)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A932D00  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [0]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [0]));  // al_ip/usart_gate.v(2124)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933140  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [3]));  // al_ip/usart_gate.v(2313)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933250  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]));  // al_ip/usart_gate.v(2295)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933360  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [0]));  // al_ip/usart_gate.v(2286)
  AL_LATCH_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933580  (
    .ar(~reset),
    .as(1'b0),
    .clk(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2F30 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [0]));  // al_ip/usart_gate.v(2223)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9337A0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [1]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [1]));  // al_ip/usart_gate.v(2133)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9338B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0]),
    .b(1'b1),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533280 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5335F0 ,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [0]}));  // al_ip/usart_gate.v(1623)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9339C0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [2]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [2]));  // al_ip/usart_gate.v(2142)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933AD0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [1]),
    .b(1'b0),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5335F0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535BC0 ,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [1]}));  // al_ip/usart_gate.v(1630)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933BE0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [5]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [5]));  // al_ip/usart_gate.v(2169)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933CF0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]));  // al_ip/usart_gate.v(2205)
  AL_LATCH_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933E00  (
    .ar(~reset),
    .as(1'b0),
    .clk(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2F30 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [2]));  // al_ip/usart_gate.v(2241)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933F10  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]));  // al_ip/usart_gate.v(2250)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934130  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [4]),
    .b(1'b0),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533B70 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534880 ,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [4]}));  // al_ip/usart_gate.v(1651)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934240  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [7]),
    .b(1'b0),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534510 ),
    .o({open_n98,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [7]}));  // al_ip/usart_gate.v(1672)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934350  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB2C0 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_vld ));  // al_ip/usart_gate.v(2079)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934460  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [2]));  // al_ip/usart_gate.v(2304)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934570  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB790 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CBF20 ));  // al_ip/usart_gate.v(2097)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934680  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]));  // al_ip/usart_gate.v(2259)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9348A0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(i_io_rx),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB790 ));  // al_ip/usart_gate.v(2106)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934CE0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2]),
    .b(1'b0),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535BC0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533120 ,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [2]}));  // al_ip/usart_gate.v(1637)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934DF0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [4]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [4]));  // al_ip/usart_gate.v(2160)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934F00  (
    .a(1'b0),
    .b(1'b0),
    .c(1'b0),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533280 ,open_n99}));  // al_ip/usart_gate.v(1679)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935010  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]));  // al_ip/usart_gate.v(2214)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935120  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [4]));  // al_ip/usart_gate.v(2322)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935230  (
    .a(1'b1),
    .b(1'b0),
    .c(1'b0),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533CD0 ,open_n100}));  // al_ip/usart_gate.v(1740)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935340  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]));  // al_ip/usart_gate.v(2268)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935560  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [6]));  // al_ip/usart_gate.v(2340)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935670  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]));  // al_ip/usart_gate.v(2196)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935780  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [3]));  // al_ip/usart_gate.v(2277)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935890  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [7]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [7]));  // al_ip/usart_gate.v(2187)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935AB0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB420 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CC810 ));  // al_ip/usart_gate.v(2115)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935CD0  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [3]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [3]));  // al_ip/usart_gate.v(2151)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935DE0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [6]),
    .b(1'b0),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533330 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534510 ,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [6]}));  // al_ip/usart_gate.v(1665)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936000  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [5]));  // al_ip/usart_gate.v(2331)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936110  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [3]),
    .b(1'b0),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533120 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533B70 ,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [3]}));  // al_ip/usart_gate.v(1644)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936220  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [6]),
    .en(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [6]));  // al_ip/usart_gate.v(2178)
  AL_LATCH_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936330  (
    .ar(~reset),
    .as(1'b0),
    .clk(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2F30 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [1]));  // al_ip/usart_gate.v(2232)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936660  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [5]),
    .b(1'b0),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534880 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533330 ,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [5]}));  // al_ip/usart_gate.v(1658)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936770  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535380 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533D80 ,open_n101}));  // al_ip/usart_gate.v(1691)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936BB0  (
    .a(1'b0),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [5]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535430 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534040 ,open_n102}));  // al_ip/usart_gate.v(1719)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A937760  (
    .a(1'b0),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [6]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534040 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535590 ,open_n103}));  // al_ip/usart_gate.v(1726)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A937BA0  (
    .a(1'b0),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [7]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535590 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5340F0 ,open_n104}));  // al_ip/usart_gate.v(1733)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A937CB0  (
    .a(1'b1),
    .b(1'b0),
    .c(1'b0),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534A90 ,open_n105}));  // al_ip/usart_gate.v(1808)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A938640  (
    .a(1'b0),
    .b(1'b1),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5340F0 ),
    .o({open_n106,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 }));  // al_ip/usart_gate.v(1745)
  AL_DFF_X \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A938970  (
    .ar(~reset),
    .as(1'b0),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB6E0 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD470 ));  // al_ip/usart_gate.v(2070)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A938EC0  (
    .a(1'b0),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [4]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534460 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535430 ,open_n107}));  // al_ip/usart_gate.v(1712)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A939EB0  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [3]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533EE0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534460 ,open_n108}));  // al_ip/usart_gate.v(1705)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93AD90  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [6]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5341A0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534250 ,open_n109}));  // al_ip/usart_gate.v(1794)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93B2E0  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [3]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534BF0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534D50 ,open_n110}));  // al_ip/usart_gate.v(1773)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C0B0  (
    .a(1'b0),
    .b(1'b1),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534300 ),
    .o({open_n111,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C93D0 }));  // al_ip/usart_gate.v(1813)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C2D0  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534B40 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5345C0 ,open_n112}));  // al_ip/usart_gate.v(1759)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C600  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [4]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534D50 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535640 ,open_n113}));  // al_ip/usart_gate.v(1780)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C710  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534A90 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534B40 ,open_n114}));  // al_ip/usart_gate.v(1752)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C820  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [5]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535640 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5341A0 ,open_n115}));  // al_ip/usart_gate.v(1787)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93D700  (
    .a(1'b1),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5345C0 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534BF0 ,open_n116}));  // al_ip/usart_gate.v(1766)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93DE70  (
    .a(1'b0),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [7]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534250 ),
    .o({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534300 ,open_n117}));  // al_ip/usart_gate.v(1801)
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(D@C)))"),
    .INIT(16'b1000110011001000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA080  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C9110 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [0]));  // al_ip/usart_gate.v(1186)
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'b00101000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA190  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FFD0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CBF20 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [0]));  // al_ip/usart_gate.v(1236)
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*~B))*~(C)+~A*(D*~B)*~(C)+~(~A)*(D*~B)*C+~A*(D*~B)*C)"),
    .INIT(16'b0011010100000101))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA2A0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0290 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [2]));  // al_ip/usart_gate.v(1270)
  AL_MAP_LUT5 #(
    .EQN("(~B*(~E*~((~D*~A))*~(C)+~E*(~D*~A)*~(C)+~(~E)*(~D*~A)*C+~E*(~D*~A)*C))"),
    .INIT(32'b00000000000100000000001100010011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA3B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FF20 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [0]),
    .e(o_io_tx),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E710 ));  // al_ip/usart_gate.v(1397)
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*B*A))"),
    .INIT(16'b0000000001111111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA4C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F160 ));  // al_ip/usart_gate.v(1109)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*B*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11001000110011111111011111111111),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA5D0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A340 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F580 ));  // al_ip/usart_gate.v(1286)
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*~(B)*~(C)+E*B*~(C)+~(E)*B*C+E*B*C))*~(D)+A*(E*~(B)*~(C)+E*B*~(C)+~(E)*B*C+E*B*C)*~(D)+~(A)*(E*~(B)*~(C)+E*B*~(C)+~(E)*B*C+E*B*C)*D+A*(E*~(B)*~(C)+E*B*~(C)+~(E)*B*C+E*B*C)*D)"),
    .INIT(32'b11001111101010101100000010101010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA6E0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5D780 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A68B0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [0]));  // al_ip/usart_gate.v(266)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA7F0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F370 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F8F0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [6]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [6]));  // al_ip/usart_gate.v(336)
  AL_MAP_LUT5 #(
    .EQN("(A*~((~C*~B))*D*~(E)+A*(~C*~B)*D*~(E)+~(A)*(~C*~B)*~(D)*E+A*(~C*~B)*~(D)*E)"),
    .INIT(32'b00000000000000111010101000000000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA900  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0080 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 [2]));  // al_ip/usart_gate.v(1332)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACAA10  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F4D0 ));  // al_ip/usart_gate.v(355)
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~(C*~B)*~(A)*~(D)+~(C*~B)*A*~(D)+~(~(C*~B))*A*D+~(C*~B)*A*D))"),
    .INIT(32'b00000000000000000101010100110000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACAB20  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0080 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A68B0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F210 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 [1]));  // al_ip/usart_gate.v(246)
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(C*A)))"),
    .INIT(16'b1110110000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACAC30  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DCC0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .d(reset),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 [0]));  // al_ip/usart_gate.v(1369)
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*~B))*~(C)+~A*(D*~B)*~(C)+~(~A)*(D*~B)*C+~A*(D*~B)*C)"),
    .INIT(16'b0011010100000101))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACAD40  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F420 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [1]));  // al_ip/usart_gate.v(1090)
  AL_MAP_LUT5 #(
    .EQN("(E*A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(32'b10001000101000000000000000000000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACAE50  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C93D0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5BBF0 ));  // al_ip/usart_gate.v(1099)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACAF60  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5A80 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9D8A0 ));  // al_ip/usart_gate.v(1407)
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'b0001))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB070  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ),
    .b(o_io_tx),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DE20 ));  // al_ip/usart_gate.v(229)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB180  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CBF20 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C9110 ));  // al_ip/usart_gate.v(1127)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'b1000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB290  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A550 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A340 ));  // al_ip/usart_gate.v(1279)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB3A0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [6]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [6]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F370 ));  // al_ip/usart_gate.v(320)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB4B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [5]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FA50 ));  // al_ip/usart_gate.v(346)
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*A)))"),
    .INIT(16'b1100110010000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB5C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DC10 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [3]));  // al_ip/usart_gate.v(1149)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB6D0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [6]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F8F0 ));  // al_ip/usart_gate.v(329)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB7E0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [7]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DED0 ));  // al_ip/usart_gate.v(286)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'b10101011100010111101111111111111),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB8F0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F420 ));  // al_ip/usart_gate.v(1072)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACBA00  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [4]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [4]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F630 ));  // al_ip/usart_gate.v(372)
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*(D@A))"),
    .INIT(16'b0101000110100010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACBB10  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA01E0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD470 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB6E0 ));  // al_ip/usart_gate.v(1388)
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'b0001000001010000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACBC20  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DA00 ));  // al_ip/usart_gate.v(1342)
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'b00000010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACBD30  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ));  // al_ip/usart_gate.v(1082)
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'b10000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACBE40  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CBF20 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830C80 ));  // al_ip/usart_gate.v(1202)
  AL_MAP_LUT4 #(
    .EQN("(A*(C@(D*B)))"),
    .INIT(16'b0010100010100000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACBF50  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FFD0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CBF20 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [1]));  // al_ip/usart_gate.v(1227)
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*A)))"),
    .INIT(16'b1100100011000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC060  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FF20 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0080 ));  // al_ip/usart_gate.v(1313)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~(E*~C)*~(B)*~(D)+~(E*~C)*B*~(D)+~(~(E*~C))*B*D+~(E*~C)*B*D))"),
    .INIT(32'b00100010000010100010001000000000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC170  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C93D0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ));  // al_ip/usart_gate.v(276)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC280  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9D950 ));  // al_ip/usart_gate.v(303)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC390  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FA50 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F4D0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [5]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [5]));  // al_ip/usart_gate.v(362)
  AL_MAP_LUT4 #(
    .EQN("(A*(D@(C*B)))"),
    .INIT(16'b0010101010000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC4A0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FFD0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830C80 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [3]));  // al_ip/usart_gate.v(1210)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'b10111010000000001011101010111011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC5B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E710 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9D8A0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .e(o_io_tx),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EDF0 ));  // al_ip/usart_gate.v(1414)
  AL_MAP_LUT5 #(
    .EQN("(A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'b10111011101100001000110010000000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC6C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A68B0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5D780 ));  // al_ip/usart_gate.v(256)
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'b10000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC7D0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C9110 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DC10 ));  // al_ip/usart_gate.v(1134)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC8E0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F630 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0340 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [4]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [4]));  // al_ip/usart_gate.v(388)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC9F0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F9A0 ));  // al_ip/usart_gate.v(407)
  AL_MAP_LUT4 #(
    .EQN("(B*(A*~(C)*~(D)+~(A)*C*~(D)+A*~(C)*D+~(A)*C*D+A*C*D))"),
    .INIT(16'b1100100001001000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACCB00  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DC10 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [2]));  // al_ip/usart_gate.v(1158)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACCC10  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [4]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0340 ));  // al_ip/usart_gate.v(381)
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*~B))*~(C)+~A*(D*~B)*~(C)+~(~A)*(D*~B)*C+~A*(D*~B)*C)"),
    .INIT(16'b0011010100000101))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACCD20  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F580 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [3]));  // al_ip/usart_gate.v(1296)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACCE30  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [3]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E240 ));  // al_ip/usart_gate.v(398)
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'b00101000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACCF40  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FFD0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830C80 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [2]));  // al_ip/usart_gate.v(1219)
  AL_MAP_LUT5 #(
    .EQN("(B*~(~A*~(E@(D*C))))"),
    .INIT(32'b10001100110011001100100010001000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD050  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C9110 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [1]));  // al_ip/usart_gate.v(1176)
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'b0000000010000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD160  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C95E0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DAB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ));  // al_ip/usart_gate.v(1244)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD270  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E240 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F9A0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [3]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [3]));  // al_ip/usart_gate.v(414)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD380  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F000 ));  // al_ip/usart_gate.v(424)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'b1000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD490  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A550 ));  // al_ip/usart_gate.v(1253)
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*A)"),
    .INIT(32'b00000000100000000000000000000000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD5A0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C95E0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DAB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCA20 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA01E0 ));  // al_ip/usart_gate.v(1378)
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'b0001))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD6B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C95E0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FFD0 ));  // al_ip/usart_gate.v(1195)
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'b00000100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD7C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ));  // al_ip/usart_gate.v(295)
  AL_MAP_LUT5 #(
    .EQN("(~B*~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*~(C)+~B*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)+~(~B)*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C+~B*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C)"),
    .INIT(32'b11110011010100111010001100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD8D0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [0]),
    .e(o_io_tx),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5F070 ));  // al_ip/usart_gate.v(219)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD9E0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DED0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9D950 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [7]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [7]));  // al_ip/usart_gate.v(310)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'b1000000000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACDAF0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ));  // al_ip/usart_gate.v(1167)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~C*~B))"),
    .INIT(32'b10101010101010101010101010101000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACDC00  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ));  // al_ip/usart_gate.v(1322)
  AL_MAP_LUT5 #(
    .EQN("~((~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*~(C)*~(E)+(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*C*~(E)+~((~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))*C*E+(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*C*E)"),
    .INIT(32'b00001111000011110101010111001100),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACDD10  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EDF0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5F070 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DE20 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D50E0 ));  // al_ip/usart_gate.v(236)
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'b0000000000010000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACDE20  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5BBF0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F160 ),
    .c(reset),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 [1]));  // al_ip/usart_gate.v(1118)
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'b0001))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACDF30  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ));  // al_ip/usart_gate.v(1142)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*B*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11001000110011111111011111111111),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE040  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A550 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0290 ));  // al_ip/usart_gate.v(1260)
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'b10000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE150  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FF20 ));  // al_ip/usart_gate.v(1305)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~A*~(D*B)))"),
    .INIT(16'b0000111000001010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE260  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DA00 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4480 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 [0]));  // al_ip/usart_gate.v(1351)
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*A))"),
    .INIT(16'b0000000001110000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE370  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DCC0 ));  // al_ip/usart_gate.v(1360)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE480  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DF80 ));  // al_ip/usart_gate.v(459)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE590  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E920 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F6E0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [0]));  // al_ip/usart_gate.v(492)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE7B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FB00 ));  // al_ip/usart_gate.v(433)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'b0000010000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACED00  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FF20 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ));  // al_ip/usart_gate.v(520)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACF580  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F000 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FB00 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [2]));  // al_ip/usart_gate.v(440)
  AL_MAP_LUT5 #(
    .EQN("(D*(B*~((C*~A))*~(E)+B*(C*~A)*~(E)+~(B)*(C*~A)*E+B*(C*~A)*E))"),
    .INIT(32'b01010000000000001100110000000000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACF690  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FC60 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5BBF0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ),
    .d(reset),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 [2]));  // al_ip/usart_gate.v(510)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACF7A0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [1]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A7020 [1]));  // al_ip/usart_gate.v(537)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD0020  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F6E0 ));  // al_ip/usart_gate.v(485)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD0680  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E7C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DF80 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [1]));  // al_ip/usart_gate.v(466)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD0DF0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E920 ));  // al_ip/usart_gate.v(476)
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'b11001000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD1340  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FC60 ));  // al_ip/usart_gate.v(502)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD1670  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA63600 ));  // al_ip/usart_gate.v(529)
  AL_MAP_LUT5 #(
    .EQN("(A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'b11111010110010100011101000001010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD1780  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A7020 [1]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA60730 ));  // al_ip/usart_gate.v(545)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD2220  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E7C0 ));  // al_ip/usart_gate.v(450)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'b10101010000011001111111100111111),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD2BB0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [7]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FDC0 ));  // al_ip/usart_gate.v(603)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111000010111111011100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD2DD0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E0E0 ));  // al_ip/usart_gate.v(565)
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'b0000010010001100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD3100  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [6]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EA80 ));  // al_ip/usart_gate.v(633)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'b0000001000000111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD3320  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [5]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EC90 ));  // al_ip/usart_gate.v(680)
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'b0000010010001100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD3A90  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [5]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [6]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EBE0 ));  // al_ip/usart_gate.v(671)
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'b0000010010001100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD3CB0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [3]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [4]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA22E0 ));  // al_ip/usart_gate.v(747)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'b0000001000000111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD4530  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [6]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [6]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E9D0 ));  // al_ip/usart_gate.v(642)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~(~C*~B)))"),
    .INIT(32'b10101010101010101010101000000010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD4640  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E190 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EA80 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E9D0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [6]));  // al_ip/usart_gate.v(651)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111001101010000000000000101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD4860  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FDC0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [7]));  // al_ip/usart_gate.v(613)
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'b0000010010001100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD5740  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F790 ));  // al_ip/usart_gate.v(575)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111000010111111011100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD5960  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [6]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E190 ));  // al_ip/usart_gate.v(623)
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'b0000010010001100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD5A70  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [4]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EF50 ));  // al_ip/usart_gate.v(709)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'b0000001000000111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD5C90  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FD10 ));  // al_ip/usart_gate.v(584)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111000010111111011100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD5DA0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [4]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EEA0 ));  // al_ip/usart_gate.v(699)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~(~C*~B)))"),
    .INIT(32'b10101010101010101010101000000010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD5EB0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EB30 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EBE0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EC90 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [5]));  // al_ip/usart_gate.v(689)
  AL_MAP_LUT5 #(
    .EQN("((B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)*~(E)*~(D)+(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)*E*~(D)+~((B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))*E*D+(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)*E*D)"),
    .INIT(32'b11111111101011000000000010101100),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD62F0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA63600 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA60730 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [1]));  // al_ip/usart_gate.v(555)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111000010111111011100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6510  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [5]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [6]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EB30 ));  // al_ip/usart_gate.v(661)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'b0000001000000111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6620  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [4]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [4]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1AA0 ));  // al_ip/usart_gate.v(718)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~(~C*~B)))"),
    .INIT(32'b10101010101010101010101000000010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6730  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EEA0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EF50 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1AA0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [4]));  // al_ip/usart_gate.v(727)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111000010111111011100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6840  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [3]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [4]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1100 ));  // al_ip/usart_gate.v(737)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~(~C*~B)))"),
    .INIT(32'b10101010101010101010101000000010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6B70  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E0E0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F790 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FD10 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [0]));  // al_ip/usart_gate.v(593)
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'b0110))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6C80  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 [1]));  // al_ip/usart_gate.v(861)
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'b00000010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6FB0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ));  // al_ip/usart_gate.v(954)
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(B*~(D*~C)))"),
    .INIT(16'b1110101011101110))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD72E0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4480 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5B30 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D3FB0 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5BE0 ));  // al_ip/usart_gate.v(918)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'b1000000000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD73F0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A832EE0 ));  // al_ip/usart_gate.v(936)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'b1000000000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7500  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C95E0 ));  // al_ip/usart_gate.v(978)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'b1000000000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7610  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DAB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DB60 ));  // al_ip/usart_gate.v(1003)
  AL_MAP_LUT4 #(
    .EQN("(D*~((~C*B))*~(A)+D*(~C*B)*~(A)+~(D)*(~C*B)*A+D*(~C*B)*A)"),
    .INIT(16'b0101110100001000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7720  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCA20 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CC810 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB420 ));  // al_ip/usart_gate.v(994)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7940  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [0]));  // al_ip/usart_gate.v(854)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'b1000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7A50  (
    .a(\u_PERIPH_TOP/u_USART2RIB/tx_en ),
    .b(\u_PERIPH_TOP/u_USART2RIB/tx_rdy ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ));  // al_ip/usart_gate.v(875)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7B60  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [5]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [5]));  // al_ip/usart_gate.v(819)
  AL_MAP_LUT4 #(
    .EQN("~(D@C@B@A)"),
    .INIT(16'b1001011001101001))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7C70  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [6]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E500 ));  // al_ip/usart_gate.v(890)
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~C)*~(A)*~(B)+~(D*~C)*A*~(B)+~(~(D*~C))*A*B+~(D*~C)*A*B)"),
    .INIT(16'b0100011101000100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7D80  (
    .a(\u_PERIPH_TOP/u_USART2RIB/tx_en ),
    .b(\u_PERIPH_TOP/u_USART2RIB/tx_rdy ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5B30 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D3FB0 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4320 ));  // al_ip/usart_gate.v(927)
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'b10100010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7E90  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA03F0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB840 ));  // al_ip/usart_gate.v(1021)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD81C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [4]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [4]));  // al_ip/usart_gate.v(826)
  AL_MAP_LUT4 #(
    .EQN("(B*~((D@C))*~(A)+B*(D@C)*~(A)+~(B)*(D@C)*A+B*(D@C)*A)"),
    .INIT(16'b0100111011100100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8600  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DB60 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCD90 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD470 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCA20 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA03F0 ));  // al_ip/usart_gate.v(1012)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'b0000001000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8710  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4480 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ));  // al_ip/usart_gate.v(1029)
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'b0000000000000001))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8820  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A68B0 [0]));  // al_ip/usart_gate.v(1047)
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'b1111101100000010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8930  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D3FB0 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4C10 ));  // al_ip/usart_gate.v(909)
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'b0101111100001000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8A40  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C93D0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_vld ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A550340 ));  // al_ip/usart_gate.v(945)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'b1000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8D70  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F210 ));  // al_ip/usart_gate.v(1056)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8E80  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DAB0 ));  // al_ip/usart_gate.v(962)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'b1000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8F90  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C95E0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A832AC0 ));  // al_ip/usart_gate.v(987)
  AL_MAP_LUT5 #(
    .EQN("~(E@D@C@B@A)"),
    .INIT(32'b01101001100101101001011001101001),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD90A0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E500 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [2]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [3]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [4]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2010 ));  // al_ip/usart_gate.v(899)
  AL_MAP_LUT4 #(
    .EQN("~(~D*C*B*A)"),
    .INIT(16'b1111111101111111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD91B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A68B0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F210 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2F30 ));  // al_ip/usart_gate.v(1063)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD92C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [3]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [3]));  // al_ip/usart_gate.v(833)
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'b0000000000000010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD93D0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD890 ));  // al_ip/usart_gate.v(1038)
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'b01111000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD95F0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 [2]));  // al_ip/usart_gate.v(882)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD9920  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [1]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [1]));  // al_ip/usart_gate.v(847)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD9C50  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [2]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [2]));  // al_ip/usart_gate.v(840)
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'b1110))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD9D60  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCD90 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CC810 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/rx_err ));  // al_ip/usart_gate.v(868)
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(A)*~(C)+(D*~B)*A*~(C)+~((D*~B))*A*C+(D*~B)*A*C)"),
    .INIT(16'b1010001110100000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD9E70  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A550340 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DAB0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_vld ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB2C0 ));  // al_ip/usart_gate.v(969)
  AL_DFF_X \u_internal_reset/reg0_b0  (
    .ar(~n1),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_internal_reset/synch_regs_q [0]));  // ../RTL/core/reset.v(16)
  AL_DFF_X \u_internal_reset/reg0_b1  (
    .ar(~n1),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_internal_reset/synch_regs_q [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_internal_reset/synch_regs_q [1]));  // ../RTL/core/reset.v(16)
  AL_DFF_X \u_internal_reset/reg0_b2  (
    .ar(~n1),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_internal_reset/synch_regs_q [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_internal_reset/synch_regs_q [2]));  // ../RTL/core/reset.v(16)
  AL_DFF_X \u_internal_reset/reg0_b3  (
    .ar(~n1),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_internal_reset/synch_regs_q [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_internal_reset/synch_regs_q [3]));  // ../RTL/core/reset.v(16)
  AL_DFF_X \u_internal_reset/reg0_b4  (
    .ar(~n1),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_internal_reset/synch_regs_q [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(reset));  // ../RTL/core/reset.v(16)
  EG_LOGIC_BUFG \u_pll/bufg_feedback  (
    .i(\u_pll/clk0_buf ),
    .o(clk_84mhz));  // al_ip/pll.v(34)
  EG_PHY_PLL #(
    .CLKC0_CPHASE(11),
    .CLKC0_DIV(12),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(1),
    .CLKC1_DIV(1),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("DISABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(1),
    .CLKC2_DIV(1),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("DISABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(7),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(0),
    .GMC_TEST(14),
    .ICP_CURRENT(9),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(2),
    .LPF_CAPACITOR(2),
    .LPF_RESISTOR(8),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(2),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \u_pll/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(clk_84mhz),
    .load_reg(1'b0),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(i_clk),
    .reset(n0),
    .stdby(1'b0),
    .clkc({open_n118,open_n119,open_n120,open_n121,\u_pll/clk0_buf }),
    .extlock(extlock));  // al_ip/pll.v(57)

endmodule 

module CORE_TOP  // ../RTL/soc_top/core_top.v(8)
  (
  i_clk,
  i_ribp_gnt,
  i_ribp_rdata,
  i_ribp_rsp,
  i_ribx_gnt,
  i_ribx_rdata,
  i_ribx_rsp,
  i_rstn,
  o_ribp_addr,
  o_ribp_mask,
  o_ribp_rdy,
  o_ribp_req,
  o_ribp_wdata,
  o_ribp_wrcs,
  o_ribx_addr,
  o_ribx_mask,
  o_ribx_rdy,
  o_ribx_req,
  o_ribx_wdata,
  o_ribx_wrcs
  );

  input i_clk;  // ../RTL/soc_top/core_top.v(9)
  input i_ribp_gnt;  // ../RTL/soc_top/core_top.v(31)
  input [31:0] i_ribp_rdata;  // ../RTL/soc_top/core_top.v(29)
  input i_ribp_rsp;  // ../RTL/soc_top/core_top.v(32)
  input i_ribx_gnt;  // ../RTL/soc_top/core_top.v(19)
  input [31:0] i_ribx_rdata;  // ../RTL/soc_top/core_top.v(17)
  input i_ribx_rsp;  // ../RTL/soc_top/core_top.v(20)
  input i_rstn;  // ../RTL/soc_top/core_top.v(10)
  output [31:0] o_ribp_addr;  // ../RTL/soc_top/core_top.v(25)
  output [3:0] o_ribp_mask;  // ../RTL/soc_top/core_top.v(27)
  output o_ribp_rdy;  // ../RTL/soc_top/core_top.v(33)
  output o_ribp_req;  // ../RTL/soc_top/core_top.v(30)
  output [31:0] o_ribp_wdata;  // ../RTL/soc_top/core_top.v(28)
  output o_ribp_wrcs;  // ../RTL/soc_top/core_top.v(26)
  output [31:0] o_ribx_addr;  // ../RTL/soc_top/core_top.v(13)
  output [3:0] o_ribx_mask;  // ../RTL/soc_top/core_top.v(15)
  output o_ribx_rdy;  // ../RTL/soc_top/core_top.v(21)
  output o_ribx_req;  // ../RTL/soc_top/core_top.v(18)
  output [31:0] o_ribx_wdata;  // ../RTL/soc_top/core_top.v(16)
  output o_ribx_wrcs;  // ../RTL/soc_top/core_top.v(14)

  wire [1:0] \RIB_ARB0/sel_tag ;  // ../RTL/core/rib.v(78)
  wire [7:0] \RIB_ARB0/sel_tag_id ;  // ../RTL/core/rib.v(113)
  wire [31:0] \RIB_ARB1/n20 ;
  wire [1:0] \RIB_ARB1/n7 ;
  wire [2:0] \RIB_ARB1/sel_tag ;  // ../RTL/core/rib.v(78)
  wire [7:0] \RIB_ARB1/sel_tag_id ;  // ../RTL/core/rib.v(113)
  wire [1:0] \RIB_ARB2/sel_tag ;  // ../RTL/core/rib.v(216)
  wire [1:0] \RIB_ARB2/sel_tag_id ;  // ../RTL/core/rib.v(252)
  wire [31:0] arb1_rdata1;  // ../RTL/soc_top/core_top.v(173)
  wire [31:0] arb2_addr0;  // ../RTL/soc_top/core_top.v(241)
  wire [3:0] arb2_mask0;  // ../RTL/soc_top/core_top.v(243)
  wire [31:0] arb2_rdata0;  // ../RTL/soc_top/core_top.v(245)
  wire [31:0] arb2_wdata0;  // ../RTL/soc_top/core_top.v(244)
  wire [31:0] rib_addr0;  // ../RTL/soc_top/core_top.v(37)
  wire [31:0] rib_addr1;  // ../RTL/soc_top/core_top.v(48)
  wire [3:0] rib_mask1;  // ../RTL/soc_top/core_top.v(50)
  wire [31:0] rib_rdata0;  // ../RTL/soc_top/core_top.v(41)
  wire [31:0] rib_rdata1;  // ../RTL/soc_top/core_top.v(52)
  wire [31:0] rib_wdata1;  // ../RTL/soc_top/core_top.v(51)
  wire [3:0] \u_DTCM_CTRL/bram_wea ;  // ../RTL/periph/bram2rib.v(27)
  wire [3:0] \u_ITCM_CTRL/bram_wea ;  // ../RTL/periph/bram2rib.v(98)
  wire \RIB_ARB0/default_cs ;  // ../RTL/core/rib.v(112)
  wire \RIB_ARB0/default_cs_neg ;
  wire \RIB_ARB0/handshake_rdy ;  // ../RTL/core/rib.v(114)
  wire \RIB_ARB0/handshake_rdy_last ;  // ../RTL/core/rib.v(117)
  wire \RIB_ARB0/mux3_b0_sel_is_0_o ;
  wire \RIB_ARB0/n2 ;
  wire \RIB_ARB0/n3 ;
  wire \RIB_ARB0/n5 ;
  wire \RIB_ARB0/n6 ;
  wire \RIB_ARB0/sel_tag_id[0]_neg ;
  wire \RIB_ARB1/default_cs ;  // ../RTL/core/rib.v(112)
  wire \RIB_ARB1/handshake_rdy ;  // ../RTL/core/rib.v(114)
  wire \RIB_ARB1/handshake_rdy_last ;  // ../RTL/core/rib.v(117)
  wire \RIB_ARB1/n0 ;
  wire \RIB_ARB1/n1 ;
  wire \RIB_ARB1/n13 ;
  wire \RIB_ARB1/n2 ;
  wire \RIB_ARB1/n3 ;
  wire \RIB_ARB1/n5 ;
  wire \RIB_ARB1/n6 ;
  wire \RIB_ARB2/handshake_rdy ;  // ../RTL/core/rib.v(253)
  wire \RIB_ARB2/handshake_rdy_last ;  // ../RTL/core/rib.v(256)
  wire \RIB_ARB2/mux4_b0_sel_is_2_o ;
  wire \RIB_ARB2/n1 ;
  wire \RIB_ARB2/n2 ;
  wire \RIB_ARB2/n6 ;
  wire \RIB_ARB2/n7 ;
  wire arb0_gnt0;  // ../RTL/soc_top/core_top.v(95)
  wire arb0_req0;  // ../RTL/soc_top/core_top.v(94)
  wire arb0_rsp0;  // ../RTL/soc_top/core_top.v(96)
  wire arb1_gnt0;  // ../RTL/soc_top/core_top.v(165)
  wire arb1_req0;  // ../RTL/soc_top/core_top.v(164)
  wire arb1_req1;  // ../RTL/soc_top/core_top.v(174)
  wire arb1_rsp0;  // ../RTL/soc_top/core_top.v(166)
  wire arb1_rsp1;  // ../RTL/soc_top/core_top.v(176)
  wire arb2_req0;  // ../RTL/soc_top/core_top.v(246)
  wire arb2_rsp0;  // ../RTL/soc_top/core_top.v(248)
  wire arb2_wrcs0;  // ../RTL/soc_top/core_top.v(242)
  wire rib_gnt1;  // ../RTL/soc_top/core_top.v(54)
  wire rib_req0;  // ../RTL/soc_top/core_top.v(42)
  wire rib_req1;  // ../RTL/soc_top/core_top.v(53)
  wire rib_rsp1;  // ../RTL/soc_top/core_top.v(55)
  wire rib_wrcs1;  // ../RTL/soc_top/core_top.v(49)
  wire \u_DTCM_CTRL/n0 ;
  wire \u_ITCM_CTRL/n0 ;

  assign o_ribp_addr[31] = rib_addr1[31];
  assign o_ribp_addr[30] = rib_addr1[30];
  assign o_ribp_addr[29] = rib_addr1[29];
  assign o_ribp_addr[28] = rib_addr1[28];
  assign o_ribp_addr[27] = rib_addr1[27];
  assign o_ribp_addr[26] = rib_addr1[26];
  assign o_ribp_addr[25] = rib_addr1[25];
  assign o_ribp_addr[24] = rib_addr1[24];
  assign o_ribp_addr[15] = rib_addr1[15];
  assign o_ribp_addr[14] = rib_addr1[14];
  assign o_ribp_addr[13] = rib_addr1[13];
  assign o_ribp_addr[12] = rib_addr1[12];
  assign o_ribp_addr[11] = rib_addr1[11];
  assign o_ribp_addr[10] = rib_addr1[10];
  assign o_ribp_addr[9] = rib_addr1[9];
  assign o_ribp_addr[8] = rib_addr1[8];
  assign o_ribp_addr[7] = rib_addr1[7];
  assign o_ribp_addr[6] = rib_addr1[6];
  assign o_ribp_addr[5] = rib_addr1[5];
  assign o_ribp_addr[4] = rib_addr1[4];
  assign o_ribp_addr[3] = rib_addr1[3];
  assign o_ribp_addr[2] = rib_addr1[2];
  assign o_ribp_addr[1] = 1'b0;
  assign o_ribp_addr[0] = 1'b0;
  assign o_ribp_mask[3] = rib_mask1[3];
  assign o_ribp_mask[2] = rib_mask1[2];
  assign o_ribp_mask[1] = rib_mask1[1];
  assign o_ribp_mask[0] = rib_mask1[0];
  assign o_ribp_wdata[31] = rib_wdata1[31];
  assign o_ribp_wdata[30] = rib_wdata1[30];
  assign o_ribp_wdata[29] = rib_wdata1[29];
  assign o_ribp_wdata[28] = rib_wdata1[28];
  assign o_ribp_wdata[27] = rib_wdata1[27];
  assign o_ribp_wdata[26] = rib_wdata1[26];
  assign o_ribp_wdata[25] = rib_wdata1[25];
  assign o_ribp_wdata[24] = rib_wdata1[24];
  assign o_ribp_wdata[23] = rib_wdata1[23];
  assign o_ribp_wdata[22] = rib_wdata1[22];
  assign o_ribp_wdata[21] = rib_wdata1[21];
  assign o_ribp_wdata[20] = rib_wdata1[20];
  assign o_ribp_wdata[19] = rib_wdata1[19];
  assign o_ribp_wdata[18] = rib_wdata1[18];
  assign o_ribp_wdata[17] = rib_wdata1[17];
  assign o_ribp_wdata[16] = rib_wdata1[16];
  assign o_ribp_wdata[15] = rib_wdata1[15];
  assign o_ribp_wdata[14] = rib_wdata1[14];
  assign o_ribp_wdata[13] = rib_wdata1[13];
  assign o_ribp_wdata[12] = rib_wdata1[12];
  assign o_ribp_wdata[11] = rib_wdata1[11];
  assign o_ribp_wdata[10] = rib_wdata1[10];
  assign o_ribp_wdata[9] = rib_wdata1[9];
  assign o_ribp_wdata[8] = rib_wdata1[8];
  assign o_ribp_wdata[7] = rib_wdata1[7];
  assign o_ribp_wdata[6] = rib_wdata1[6];
  assign o_ribp_wdata[5] = rib_wdata1[5];
  assign o_ribp_wdata[4] = rib_wdata1[4];
  assign o_ribp_wdata[3] = rib_wdata1[3];
  assign o_ribp_wdata[2] = rib_wdata1[2];
  assign o_ribp_wdata[1] = rib_wdata1[1];
  assign o_ribp_wdata[0] = rib_wdata1[0];
  assign o_ribp_wrcs = rib_wrcs1;
  not \RIB_ARB0/default_cs_inv  (\RIB_ARB0/default_cs_neg , \RIB_ARB0/default_cs );
  AL_DFF_X \RIB_ARB0/default_cs_reg  (
    .ar(1'b0),
    .as(~i_rstn),
    .clk(i_clk),
    .d(\RIB_ARB0/n3 ),
    .en(\RIB_ARB0/n6 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\RIB_ARB0/default_cs ));  // ../RTL/core/rib.v(121)
  eq_w8 \RIB_ARB0/eq0  (
    .i0(rib_addr0[31:24]),
    .i1(8'b00000000),
    .o(\RIB_ARB0/sel_tag [0]));  // ../RTL/core/rib.v(83)
  eq_w8 \RIB_ARB0/eq1  (
    .i0(rib_addr0[31:24]),
    .i1(8'b00000010),
    .o(\RIB_ARB0/sel_tag [1]));  // ../RTL/core/rib.v(83)
  AL_DFF_X \RIB_ARB0/handshake_rdy_last_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\RIB_ARB0/handshake_rdy ),
    .en(\RIB_ARB0/n6 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\RIB_ARB0/handshake_rdy_last ));  // ../RTL/core/rib.v(121)
  AL_MUX \RIB_ARB0/mux3_b0  (
    .i0(1'b0),
    .i1(arb2_rdata0[0]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[0]));
  and \RIB_ARB0/mux3_b0_sel_is_0  (\RIB_ARB0/mux3_b0_sel_is_0_o , \RIB_ARB0/default_cs_neg , \RIB_ARB0/sel_tag_id[0]_neg );
  AL_MUX \RIB_ARB0/mux3_b1  (
    .i0(1'b0),
    .i1(arb2_rdata0[1]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[1]));
  AL_MUX \RIB_ARB0/mux3_b10  (
    .i0(1'b0),
    .i1(arb2_rdata0[10]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[10]));
  AL_MUX \RIB_ARB0/mux3_b11  (
    .i0(1'b0),
    .i1(arb2_rdata0[11]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[11]));
  AL_MUX \RIB_ARB0/mux3_b12  (
    .i0(1'b0),
    .i1(arb2_rdata0[12]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[12]));
  AL_MUX \RIB_ARB0/mux3_b13  (
    .i0(1'b0),
    .i1(arb2_rdata0[13]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[13]));
  AL_MUX \RIB_ARB0/mux3_b14  (
    .i0(1'b0),
    .i1(arb2_rdata0[14]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[14]));
  AL_MUX \RIB_ARB0/mux3_b15  (
    .i0(1'b0),
    .i1(arb2_rdata0[15]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[15]));
  AL_MUX \RIB_ARB0/mux3_b16  (
    .i0(1'b0),
    .i1(arb2_rdata0[16]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[16]));
  AL_MUX \RIB_ARB0/mux3_b17  (
    .i0(1'b0),
    .i1(arb2_rdata0[17]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[17]));
  AL_MUX \RIB_ARB0/mux3_b18  (
    .i0(1'b0),
    .i1(arb2_rdata0[18]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[18]));
  AL_MUX \RIB_ARB0/mux3_b19  (
    .i0(1'b0),
    .i1(arb2_rdata0[19]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[19]));
  AL_MUX \RIB_ARB0/mux3_b2  (
    .i0(1'b0),
    .i1(arb2_rdata0[2]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[2]));
  AL_MUX \RIB_ARB0/mux3_b20  (
    .i0(1'b0),
    .i1(arb2_rdata0[20]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[20]));
  AL_MUX \RIB_ARB0/mux3_b21  (
    .i0(1'b0),
    .i1(arb2_rdata0[21]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[21]));
  AL_MUX \RIB_ARB0/mux3_b22  (
    .i0(1'b0),
    .i1(arb2_rdata0[22]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[22]));
  AL_MUX \RIB_ARB0/mux3_b23  (
    .i0(1'b0),
    .i1(arb2_rdata0[23]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[23]));
  AL_MUX \RIB_ARB0/mux3_b24  (
    .i0(1'b0),
    .i1(arb2_rdata0[24]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[24]));
  AL_MUX \RIB_ARB0/mux3_b25  (
    .i0(1'b0),
    .i1(arb2_rdata0[25]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[25]));
  AL_MUX \RIB_ARB0/mux3_b26  (
    .i0(1'b0),
    .i1(arb2_rdata0[26]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[26]));
  AL_MUX \RIB_ARB0/mux3_b27  (
    .i0(1'b0),
    .i1(arb2_rdata0[27]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[27]));
  AL_MUX \RIB_ARB0/mux3_b28  (
    .i0(1'b0),
    .i1(arb2_rdata0[28]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[28]));
  AL_MUX \RIB_ARB0/mux3_b29  (
    .i0(1'b0),
    .i1(arb2_rdata0[29]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[29]));
  AL_MUX \RIB_ARB0/mux3_b3  (
    .i0(1'b0),
    .i1(arb2_rdata0[3]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[3]));
  AL_MUX \RIB_ARB0/mux3_b30  (
    .i0(1'b0),
    .i1(arb2_rdata0[30]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[30]));
  AL_MUX \RIB_ARB0/mux3_b31  (
    .i0(1'b0),
    .i1(arb2_rdata0[31]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[31]));
  AL_MUX \RIB_ARB0/mux3_b4  (
    .i0(1'b0),
    .i1(arb2_rdata0[4]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[4]));
  AL_MUX \RIB_ARB0/mux3_b5  (
    .i0(1'b0),
    .i1(arb2_rdata0[5]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[5]));
  AL_MUX \RIB_ARB0/mux3_b6  (
    .i0(1'b0),
    .i1(arb2_rdata0[6]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[6]));
  AL_MUX \RIB_ARB0/mux3_b7  (
    .i0(1'b0),
    .i1(arb2_rdata0[7]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[7]));
  AL_MUX \RIB_ARB0/mux3_b8  (
    .i0(1'b0),
    .i1(arb2_rdata0[8]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[8]));
  AL_MUX \RIB_ARB0/mux3_b9  (
    .i0(1'b0),
    .i1(arb2_rdata0[9]),
    .sel(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .o(rib_rdata0[9]));
  AL_DFF_X \RIB_ARB0/reg0_b0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\RIB_ARB0/sel_tag [1]),
    .en(\RIB_ARB0/n6 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\RIB_ARB0/sel_tag_id [0]));  // ../RTL/core/rib.v(121)
  not \RIB_ARB0/sel_tag_id[0]_inv  (\RIB_ARB0/sel_tag_id[0]_neg , \RIB_ARB0/sel_tag_id [0]);
  and \RIB_ARB0/u14  (arb0_req0, rib_req0, \RIB_ARB0/sel_tag [0]);  // ../RTL/core/rib.v(90)
  not \RIB_ARB0/u23  (\RIB_ARB0/n3 , \RIB_ARB0/n2 );  // ../RTL/core/rib.v(105)
  and \RIB_ARB0/u25  (\RIB_ARB0/handshake_rdy , rib_req0, arb0_gnt0);  // ../RTL/core/rib.v(114)
  not \RIB_ARB0/u31  (\RIB_ARB0/n5 , \RIB_ARB0/handshake_rdy_last );  // ../RTL/core/rib.v(128)
  or \RIB_ARB0/u32  (\RIB_ARB0/n6 , arb0_rsp0, \RIB_ARB0/n5 );  // ../RTL/core/rib.v(128)
  or \RIB_ARB0/u33  (\RIB_ARB0/n2 , \RIB_ARB0/sel_tag [0], \RIB_ARB0/sel_tag [1]);  // ../RTL/core/rib.v(105)
  AL_DFF_X \RIB_ARB1/default_cs_reg  (
    .ar(1'b0),
    .as(~i_rstn),
    .clk(i_clk),
    .d(\RIB_ARB1/n3 ),
    .en(\RIB_ARB1/n6 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\RIB_ARB1/default_cs ));  // ../RTL/core/rib.v(121)
  eq_w8 \RIB_ARB1/eq0  (
    .i0(rib_addr1[31:24]),
    .i1(8'b00000000),
    .o(\RIB_ARB1/sel_tag [0]));  // ../RTL/core/rib.v(83)
  eq_w8 \RIB_ARB1/eq1  (
    .i0(rib_addr1[31:24]),
    .i1(8'b00000001),
    .o(\RIB_ARB1/sel_tag [1]));  // ../RTL/core/rib.v(83)
  eq_w8 \RIB_ARB1/eq2  (
    .i0(rib_addr1[31:24]),
    .i1(8'b00000010),
    .o(\RIB_ARB1/sel_tag [2]));  // ../RTL/core/rib.v(83)
  AL_DFF_X \RIB_ARB1/handshake_rdy_last_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\RIB_ARB1/handshake_rdy ),
    .en(\RIB_ARB1/n6 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\RIB_ARB1/handshake_rdy_last ));  // ../RTL/core/rib.v(121)
  binary_mux_s1_w1 \RIB_ARB1/mux1_b0  (
    .i0(\RIB_ARB1/sel_tag [1]),
    .i1(1'b0),
    .sel(\RIB_ARB1/sel_tag [2]),
    .o(\RIB_ARB1/n7 [0]));  // ../RTL/core/rib.v(69)
  binary_mux_s1_w1 \RIB_ARB1/mux1_b1  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\RIB_ARB1/sel_tag [2]),
    .o(\RIB_ARB1/n7 [1]));  // ../RTL/core/rib.v(69)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b0  (
    .i0(arb2_rdata0[0]),
    .i1(arb1_rdata1[0]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [0]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b1  (
    .i0(arb2_rdata0[1]),
    .i1(arb1_rdata1[1]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [1]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b10  (
    .i0(arb2_rdata0[10]),
    .i1(arb1_rdata1[10]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [10]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b11  (
    .i0(arb2_rdata0[11]),
    .i1(arb1_rdata1[11]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [11]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b12  (
    .i0(arb2_rdata0[12]),
    .i1(arb1_rdata1[12]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [12]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b13  (
    .i0(arb2_rdata0[13]),
    .i1(arb1_rdata1[13]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [13]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b14  (
    .i0(arb2_rdata0[14]),
    .i1(arb1_rdata1[14]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [14]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b15  (
    .i0(arb2_rdata0[15]),
    .i1(arb1_rdata1[15]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [15]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b16  (
    .i0(arb2_rdata0[16]),
    .i1(arb1_rdata1[16]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [16]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b17  (
    .i0(arb2_rdata0[17]),
    .i1(arb1_rdata1[17]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [17]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b18  (
    .i0(arb2_rdata0[18]),
    .i1(arb1_rdata1[18]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [18]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b19  (
    .i0(arb2_rdata0[19]),
    .i1(arb1_rdata1[19]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [19]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b2  (
    .i0(arb2_rdata0[2]),
    .i1(arb1_rdata1[2]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [2]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b20  (
    .i0(arb2_rdata0[20]),
    .i1(arb1_rdata1[20]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [20]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b21  (
    .i0(arb2_rdata0[21]),
    .i1(arb1_rdata1[21]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [21]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b22  (
    .i0(arb2_rdata0[22]),
    .i1(arb1_rdata1[22]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [22]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b23  (
    .i0(arb2_rdata0[23]),
    .i1(arb1_rdata1[23]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [23]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b24  (
    .i0(arb2_rdata0[24]),
    .i1(arb1_rdata1[24]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [24]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b25  (
    .i0(arb2_rdata0[25]),
    .i1(arb1_rdata1[25]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [25]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b26  (
    .i0(arb2_rdata0[26]),
    .i1(arb1_rdata1[26]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [26]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b27  (
    .i0(arb2_rdata0[27]),
    .i1(arb1_rdata1[27]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [27]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b28  (
    .i0(arb2_rdata0[28]),
    .i1(arb1_rdata1[28]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [28]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b29  (
    .i0(arb2_rdata0[29]),
    .i1(arb1_rdata1[29]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [29]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b3  (
    .i0(arb2_rdata0[3]),
    .i1(arb1_rdata1[3]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [3]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b30  (
    .i0(arb2_rdata0[30]),
    .i1(arb1_rdata1[30]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [30]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b31  (
    .i0(arb2_rdata0[31]),
    .i1(arb1_rdata1[31]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [31]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b4  (
    .i0(arb2_rdata0[4]),
    .i1(arb1_rdata1[4]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [4]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b5  (
    .i0(arb2_rdata0[5]),
    .i1(arb1_rdata1[5]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [5]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b6  (
    .i0(arb2_rdata0[6]),
    .i1(arb1_rdata1[6]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [6]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b7  (
    .i0(arb2_rdata0[7]),
    .i1(arb1_rdata1[7]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [7]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b8  (
    .i0(arb2_rdata0[8]),
    .i1(arb1_rdata1[8]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [8]));  // ../RTL/core/rib.v(146)
  binary_mux_s2_w1 \RIB_ARB1/mux3_b9  (
    .i0(arb2_rdata0[9]),
    .i1(arb1_rdata1[9]),
    .i2(1'b0),
    .i3(1'bx),
    .sel(\RIB_ARB1/sel_tag_id [1:0]),
    .o(\RIB_ARB1/n20 [9]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b0  (
    .i0(\RIB_ARB1/n20 [0]),
    .i1(i_ribp_rdata[0]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[0]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b1  (
    .i0(\RIB_ARB1/n20 [1]),
    .i1(i_ribp_rdata[1]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[1]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b10  (
    .i0(\RIB_ARB1/n20 [10]),
    .i1(i_ribp_rdata[10]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[10]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b11  (
    .i0(\RIB_ARB1/n20 [11]),
    .i1(i_ribp_rdata[11]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[11]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b12  (
    .i0(\RIB_ARB1/n20 [12]),
    .i1(i_ribp_rdata[12]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[12]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b13  (
    .i0(\RIB_ARB1/n20 [13]),
    .i1(i_ribp_rdata[13]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[13]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b14  (
    .i0(\RIB_ARB1/n20 [14]),
    .i1(i_ribp_rdata[14]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[14]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b15  (
    .i0(\RIB_ARB1/n20 [15]),
    .i1(i_ribp_rdata[15]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[15]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b16  (
    .i0(\RIB_ARB1/n20 [16]),
    .i1(i_ribp_rdata[16]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[16]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b17  (
    .i0(\RIB_ARB1/n20 [17]),
    .i1(i_ribp_rdata[17]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[17]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b18  (
    .i0(\RIB_ARB1/n20 [18]),
    .i1(i_ribp_rdata[18]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[18]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b19  (
    .i0(\RIB_ARB1/n20 [19]),
    .i1(i_ribp_rdata[19]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[19]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b2  (
    .i0(\RIB_ARB1/n20 [2]),
    .i1(i_ribp_rdata[2]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[2]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b20  (
    .i0(\RIB_ARB1/n20 [20]),
    .i1(i_ribp_rdata[20]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[20]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b21  (
    .i0(\RIB_ARB1/n20 [21]),
    .i1(i_ribp_rdata[21]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[21]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b22  (
    .i0(\RIB_ARB1/n20 [22]),
    .i1(i_ribp_rdata[22]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[22]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b23  (
    .i0(\RIB_ARB1/n20 [23]),
    .i1(i_ribp_rdata[23]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[23]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b24  (
    .i0(\RIB_ARB1/n20 [24]),
    .i1(i_ribp_rdata[24]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[24]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b25  (
    .i0(\RIB_ARB1/n20 [25]),
    .i1(i_ribp_rdata[25]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[25]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b26  (
    .i0(\RIB_ARB1/n20 [26]),
    .i1(i_ribp_rdata[26]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[26]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b27  (
    .i0(\RIB_ARB1/n20 [27]),
    .i1(i_ribp_rdata[27]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[27]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b28  (
    .i0(\RIB_ARB1/n20 [28]),
    .i1(i_ribp_rdata[28]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[28]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b29  (
    .i0(\RIB_ARB1/n20 [29]),
    .i1(i_ribp_rdata[29]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[29]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b3  (
    .i0(\RIB_ARB1/n20 [3]),
    .i1(i_ribp_rdata[3]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[3]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b30  (
    .i0(\RIB_ARB1/n20 [30]),
    .i1(i_ribp_rdata[30]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[30]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b31  (
    .i0(\RIB_ARB1/n20 [31]),
    .i1(i_ribp_rdata[31]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[31]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b4  (
    .i0(\RIB_ARB1/n20 [4]),
    .i1(i_ribp_rdata[4]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[4]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b5  (
    .i0(\RIB_ARB1/n20 [5]),
    .i1(i_ribp_rdata[5]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[5]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b6  (
    .i0(\RIB_ARB1/n20 [6]),
    .i1(i_ribp_rdata[6]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[6]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b7  (
    .i0(\RIB_ARB1/n20 [7]),
    .i1(i_ribp_rdata[7]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[7]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b8  (
    .i0(\RIB_ARB1/n20 [8]),
    .i1(i_ribp_rdata[8]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[8]));  // ../RTL/core/rib.v(146)
  binary_mux_s1_w1 \RIB_ARB1/mux4_b9  (
    .i0(\RIB_ARB1/n20 [9]),
    .i1(i_ribp_rdata[9]),
    .sel(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[9]));  // ../RTL/core/rib.v(146)
  AL_DFF_X \RIB_ARB1/reg0_b0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\RIB_ARB1/n7 [0]),
    .en(\RIB_ARB1/n6 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\RIB_ARB1/sel_tag_id [0]));  // ../RTL/core/rib.v(121)
  AL_DFF_X \RIB_ARB1/reg0_b1  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\RIB_ARB1/n7 [1]),
    .en(\RIB_ARB1/n6 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\RIB_ARB1/sel_tag_id [1]));  // ../RTL/core/rib.v(121)
  or \RIB_ARB1/u129  (\RIB_ARB1/n2 , \RIB_ARB1/sel_tag [0], \RIB_ARB1/n13 );  // ../RTL/core/rib.v(105)
  or \RIB_ARB1/u195  (\RIB_ARB1/n1 , arb1_rsp0, arb1_rsp1);  // ../RTL/core/rib.v(97)
  or \RIB_ARB1/u196  (\RIB_ARB1/n0 , arb1_gnt0, arb1_req1);  // ../RTL/core/rib.v(95)
  and \RIB_ARB1/u197  (arb1_req1, rib_req1, \RIB_ARB1/sel_tag [1]);  // ../RTL/core/rib.v(90)
  and \RIB_ARB1/u20  (arb1_req0, rib_req1, \RIB_ARB1/sel_tag [0]);  // ../RTL/core/rib.v(90)
  or \RIB_ARB1/u21  (rib_gnt1, \RIB_ARB1/n0 , i_ribp_gnt);  // ../RTL/core/rib.v(95)
  or \RIB_ARB1/u23  (rib_rsp1, \RIB_ARB1/n1 , i_ribp_rsp);  // ../RTL/core/rib.v(97)
  not \RIB_ARB1/u29  (\RIB_ARB1/n3 , \RIB_ARB1/n2 );  // ../RTL/core/rib.v(105)
  and \RIB_ARB1/u30  (o_ribp_req, rib_req1, \RIB_ARB1/n3 );  // ../RTL/core/rib.v(105)
  and \RIB_ARB1/u31  (\RIB_ARB1/handshake_rdy , rib_req1, rib_gnt1);  // ../RTL/core/rib.v(114)
  not \RIB_ARB1/u37  (\RIB_ARB1/n5 , \RIB_ARB1/handshake_rdy_last );  // ../RTL/core/rib.v(128)
  or \RIB_ARB1/u38  (\RIB_ARB1/n6 , rib_rsp1, \RIB_ARB1/n5 );  // ../RTL/core/rib.v(128)
  or \RIB_ARB1/u39  (\RIB_ARB1/n13 , \RIB_ARB1/sel_tag [1], \RIB_ARB1/sel_tag [2]);  // ../RTL/core/rib.v(105)
  eq_w1 \RIB_ARB2/eq0  (
    .i0(1'b0),
    .i1(\RIB_ARB2/sel_tag_id [0]),
    .o(\RIB_ARB2/n6 ));  // ../RTL/core/rib.v(276)
  eq_w1 \RIB_ARB2/eq1  (
    .i0(1'b1),
    .i1(\RIB_ARB2/sel_tag_id [0]),
    .o(\RIB_ARB2/n7 ));  // ../RTL/core/rib.v(276)
  AL_DFF_X \RIB_ARB2/handshake_rdy_last_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\RIB_ARB2/handshake_rdy ),
    .en(\RIB_ARB2/n2 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\RIB_ARB2/handshake_rdy_last ));  // ../RTL/core/rib.v(260)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b10  (
    .i0(rib_addr0[10]),
    .i1(rib_addr1[10]),
    .sel(arb1_req0),
    .o(arb2_addr0[10]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b11  (
    .i0(rib_addr0[11]),
    .i1(rib_addr1[11]),
    .sel(arb1_req0),
    .o(arb2_addr0[11]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b12  (
    .i0(rib_addr0[12]),
    .i1(rib_addr1[12]),
    .sel(arb1_req0),
    .o(arb2_addr0[12]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b13  (
    .i0(rib_addr0[13]),
    .i1(rib_addr1[13]),
    .sel(arb1_req0),
    .o(arb2_addr0[13]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b14  (
    .i0(rib_addr0[14]),
    .i1(rib_addr1[14]),
    .sel(arb1_req0),
    .o(arb2_addr0[14]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b15  (
    .i0(rib_addr0[15]),
    .i1(rib_addr1[15]),
    .sel(arb1_req0),
    .o(arb2_addr0[15]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b2  (
    .i0(rib_addr0[2]),
    .i1(rib_addr1[2]),
    .sel(arb1_req0),
    .o(arb2_addr0[2]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b3  (
    .i0(rib_addr0[3]),
    .i1(rib_addr1[3]),
    .sel(arb1_req0),
    .o(arb2_addr0[3]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b4  (
    .i0(rib_addr0[4]),
    .i1(rib_addr1[4]),
    .sel(arb1_req0),
    .o(arb2_addr0[4]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b5  (
    .i0(rib_addr0[5]),
    .i1(rib_addr1[5]),
    .sel(arb1_req0),
    .o(arb2_addr0[5]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b6  (
    .i0(rib_addr0[6]),
    .i1(rib_addr1[6]),
    .sel(arb1_req0),
    .o(arb2_addr0[6]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b7  (
    .i0(rib_addr0[7]),
    .i1(rib_addr1[7]),
    .sel(arb1_req0),
    .o(arb2_addr0[7]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b8  (
    .i0(rib_addr0[8]),
    .i1(rib_addr1[8]),
    .sel(arb1_req0),
    .o(arb2_addr0[8]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux0_b9  (
    .i0(rib_addr0[9]),
    .i1(rib_addr1[9]),
    .sel(arb1_req0),
    .o(arb2_addr0[9]));  // ../RTL/core/rib.v(238)
  binary_mux_s1_w1 \RIB_ARB2/mux1_b0  (
    .i0(1'b1),
    .i1(rib_mask1[0]),
    .sel(arb1_req0),
    .o(arb2_mask0[0]));  // ../RTL/core/rib.v(242)
  binary_mux_s1_w1 \RIB_ARB2/mux1_b1  (
    .i0(1'b1),
    .i1(rib_mask1[1]),
    .sel(arb1_req0),
    .o(arb2_mask0[1]));  // ../RTL/core/rib.v(242)
  binary_mux_s1_w1 \RIB_ARB2/mux1_b2  (
    .i0(1'b1),
    .i1(rib_mask1[2]),
    .sel(arb1_req0),
    .o(arb2_mask0[2]));  // ../RTL/core/rib.v(242)
  binary_mux_s1_w1 \RIB_ARB2/mux1_b3  (
    .i0(1'b1),
    .i1(rib_mask1[3]),
    .sel(arb1_req0),
    .o(arb2_mask0[3]));  // ../RTL/core/rib.v(242)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b0  (
    .i0(1'b0),
    .i1(rib_wdata1[0]),
    .sel(arb1_req0),
    .o(arb2_wdata0[0]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b1  (
    .i0(1'b0),
    .i1(rib_wdata1[1]),
    .sel(arb1_req0),
    .o(arb2_wdata0[1]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b10  (
    .i0(1'b0),
    .i1(rib_wdata1[10]),
    .sel(arb1_req0),
    .o(arb2_wdata0[10]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b11  (
    .i0(1'b0),
    .i1(rib_wdata1[11]),
    .sel(arb1_req0),
    .o(arb2_wdata0[11]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b12  (
    .i0(1'b0),
    .i1(rib_wdata1[12]),
    .sel(arb1_req0),
    .o(arb2_wdata0[12]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b13  (
    .i0(1'b0),
    .i1(rib_wdata1[13]),
    .sel(arb1_req0),
    .o(arb2_wdata0[13]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b14  (
    .i0(1'b0),
    .i1(rib_wdata1[14]),
    .sel(arb1_req0),
    .o(arb2_wdata0[14]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b15  (
    .i0(1'b0),
    .i1(rib_wdata1[15]),
    .sel(arb1_req0),
    .o(arb2_wdata0[15]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b16  (
    .i0(1'b0),
    .i1(rib_wdata1[16]),
    .sel(arb1_req0),
    .o(arb2_wdata0[16]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b17  (
    .i0(1'b0),
    .i1(rib_wdata1[17]),
    .sel(arb1_req0),
    .o(arb2_wdata0[17]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b18  (
    .i0(1'b0),
    .i1(rib_wdata1[18]),
    .sel(arb1_req0),
    .o(arb2_wdata0[18]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b19  (
    .i0(1'b0),
    .i1(rib_wdata1[19]),
    .sel(arb1_req0),
    .o(arb2_wdata0[19]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b2  (
    .i0(1'b0),
    .i1(rib_wdata1[2]),
    .sel(arb1_req0),
    .o(arb2_wdata0[2]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b20  (
    .i0(1'b0),
    .i1(rib_wdata1[20]),
    .sel(arb1_req0),
    .o(arb2_wdata0[20]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b21  (
    .i0(1'b0),
    .i1(rib_wdata1[21]),
    .sel(arb1_req0),
    .o(arb2_wdata0[21]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b22  (
    .i0(1'b0),
    .i1(rib_wdata1[22]),
    .sel(arb1_req0),
    .o(arb2_wdata0[22]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b23  (
    .i0(1'b0),
    .i1(rib_wdata1[23]),
    .sel(arb1_req0),
    .o(arb2_wdata0[23]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b24  (
    .i0(1'b0),
    .i1(rib_wdata1[24]),
    .sel(arb1_req0),
    .o(arb2_wdata0[24]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b25  (
    .i0(1'b0),
    .i1(rib_wdata1[25]),
    .sel(arb1_req0),
    .o(arb2_wdata0[25]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b26  (
    .i0(1'b0),
    .i1(rib_wdata1[26]),
    .sel(arb1_req0),
    .o(arb2_wdata0[26]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b27  (
    .i0(1'b0),
    .i1(rib_wdata1[27]),
    .sel(arb1_req0),
    .o(arb2_wdata0[27]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b28  (
    .i0(1'b0),
    .i1(rib_wdata1[28]),
    .sel(arb1_req0),
    .o(arb2_wdata0[28]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b29  (
    .i0(1'b0),
    .i1(rib_wdata1[29]),
    .sel(arb1_req0),
    .o(arb2_wdata0[29]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b3  (
    .i0(1'b0),
    .i1(rib_wdata1[3]),
    .sel(arb1_req0),
    .o(arb2_wdata0[3]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b30  (
    .i0(1'b0),
    .i1(rib_wdata1[30]),
    .sel(arb1_req0),
    .o(arb2_wdata0[30]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b31  (
    .i0(1'b0),
    .i1(rib_wdata1[31]),
    .sel(arb1_req0),
    .o(arb2_wdata0[31]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b4  (
    .i0(1'b0),
    .i1(rib_wdata1[4]),
    .sel(arb1_req0),
    .o(arb2_wdata0[4]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b5  (
    .i0(1'b0),
    .i1(rib_wdata1[5]),
    .sel(arb1_req0),
    .o(arb2_wdata0[5]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b6  (
    .i0(1'b0),
    .i1(rib_wdata1[6]),
    .sel(arb1_req0),
    .o(arb2_wdata0[6]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b7  (
    .i0(1'b0),
    .i1(rib_wdata1[7]),
    .sel(arb1_req0),
    .o(arb2_wdata0[7]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b8  (
    .i0(1'b0),
    .i1(rib_wdata1[8]),
    .sel(arb1_req0),
    .o(arb2_wdata0[8]));  // ../RTL/core/rib.v(244)
  binary_mux_s1_w1 \RIB_ARB2/mux2_b9  (
    .i0(1'b0),
    .i1(rib_wdata1[9]),
    .sel(arb1_req0),
    .o(arb2_wdata0[9]));  // ../RTL/core/rib.v(244)
  and \RIB_ARB2/mux4_b0_sel_is_2  (\RIB_ARB2/mux4_b0_sel_is_2_o , i_rstn, \RIB_ARB2/n2 );
  AL_DFF_X \RIB_ARB2/reg0_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(arb1_req0),
    .en(\RIB_ARB2/mux4_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\RIB_ARB2/sel_tag_id [0]));  // ../RTL/core/rib.v(260)
  and \RIB_ARB2/u14  (arb0_rsp0, \RIB_ARB2/n6 , arb2_rsp0);  // ../RTL/core/rib.v(276)
  AL_MUX \RIB_ARB2/u17  (
    .i0(1'b0),
    .i1(rib_wrcs1),
    .sel(arb1_req0),
    .o(arb2_wrcs0));  // ../RTL/core/rib.v(240)
  and \RIB_ARB2/u20  (arb0_gnt0, \RIB_ARB2/sel_tag [0], arb2_req0);  // ../RTL/core/rib.v(231)
  and \RIB_ARB2/u21  (\RIB_ARB2/handshake_rdy , arb2_req0, arb2_req0);  // ../RTL/core/rib.v(253)
  not \RIB_ARB2/u27  (\RIB_ARB2/n1 , \RIB_ARB2/handshake_rdy_last );  // ../RTL/core/rib.v(265)
  or \RIB_ARB2/u28  (\RIB_ARB2/n2 , arb2_rsp0, \RIB_ARB2/n1 );  // ../RTL/core/rib.v(265)
  or \RIB_ARB2/u31  (arb2_req0, arb0_req0, arb1_req0);  // ../RTL/core/rib.v(246)
  and \RIB_ARB2/u86  (arb1_gnt0, arb1_req0, arb2_req0);  // ../RTL/core/rib.v(231)
  and \RIB_ARB2/u87  (arb1_rsp0, \RIB_ARB2/n7 , arb2_rsp0);  // ../RTL/core/rib.v(276)
  not \RIB_ARB2/u9  (\RIB_ARB2/sel_tag [0], arb1_req0);  // ../RTL/core/rib.v(221)
  AL_DFF_X \u_DTCM_CTRL/handshake_rdy_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(arb1_req1),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(arb1_rsp1));  // ../RTL/periph/bram2rib.v(37)
  binary_mux_s1_w1 \u_DTCM_CTRL/mux0_b0  (
    .i0(1'b0),
    .i1(rib_mask1[0]),
    .sel(\u_DTCM_CTRL/n0 ),
    .o(\u_DTCM_CTRL/bram_wea [0]));  // ../RTL/periph/bram2rib.v(27)
  binary_mux_s1_w1 \u_DTCM_CTRL/mux0_b1  (
    .i0(1'b0),
    .i1(rib_mask1[1]),
    .sel(\u_DTCM_CTRL/n0 ),
    .o(\u_DTCM_CTRL/bram_wea [1]));  // ../RTL/periph/bram2rib.v(27)
  binary_mux_s1_w1 \u_DTCM_CTRL/mux0_b2  (
    .i0(1'b0),
    .i1(rib_mask1[2]),
    .sel(\u_DTCM_CTRL/n0 ),
    .o(\u_DTCM_CTRL/bram_wea [2]));  // ../RTL/periph/bram2rib.v(27)
  binary_mux_s1_w1 \u_DTCM_CTRL/mux0_b3  (
    .i0(1'b0),
    .i1(rib_mask1[3]),
    .sel(\u_DTCM_CTRL/n0 ),
    .o(\u_DTCM_CTRL/bram_wea [3]));  // ../RTL/periph/bram2rib.v(27)
  and \u_DTCM_CTRL/u2  (\u_DTCM_CTRL/n0 , rib_wrcs1, arb1_req1);  // ../RTL/periph/bram2rib.v(27)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("NONE"),
    .ADDR_WIDTH_A(14),
    .ADDR_WIDTH_B(14),
    .BYTE_A(4),
    .BYTE_B(4),
    .BYTE_ENABLE(8),
    .DATA_DEPTH_A(16384),
    .DATA_DEPTH_B(16384),
    .DATA_WIDTH_A(32),
    .DATA_WIDTH_B(32),
    .DEBUGGABLE("NO"),
    .FILL_ALL("00000000000000000000000000000000"),
    .IMPLEMENT("32K"),
    .MODE("SP"),
    .PACKABLE("NO"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst  (
    .addra(rib_addr1[15:2]),
    .addrb(14'b00000000000000),
    .bea(\u_DTCM_CTRL/bram_wea ),
    .beb(4'b0000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(i_clk),
    .clkb(1'b0),
    .dia(rib_wdata1),
    .dib(32'b00000000000000000000000000000000),
    .ocea(1'b0),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(1'b0),
    .web(1'b0),
    .doa(arb1_rdata1));  // al_ip/bram_dtcm.v(53)
  AL_DFF_X \u_ITCM_CTRL/handshake_rdy_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(arb2_req0),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(arb2_rsp0));  // ../RTL/periph/bram2rib.v(110)
  binary_mux_s1_w1 \u_ITCM_CTRL/mux0_b0  (
    .i0(1'b0),
    .i1(arb2_mask0[0]),
    .sel(\u_ITCM_CTRL/n0 ),
    .o(\u_ITCM_CTRL/bram_wea [0]));  // ../RTL/periph/bram2rib.v(98)
  binary_mux_s1_w1 \u_ITCM_CTRL/mux0_b1  (
    .i0(1'b0),
    .i1(arb2_mask0[1]),
    .sel(\u_ITCM_CTRL/n0 ),
    .o(\u_ITCM_CTRL/bram_wea [1]));  // ../RTL/periph/bram2rib.v(98)
  binary_mux_s1_w1 \u_ITCM_CTRL/mux0_b2  (
    .i0(1'b0),
    .i1(arb2_mask0[2]),
    .sel(\u_ITCM_CTRL/n0 ),
    .o(\u_ITCM_CTRL/bram_wea [2]));  // ../RTL/periph/bram2rib.v(98)
  binary_mux_s1_w1 \u_ITCM_CTRL/mux0_b3  (
    .i0(1'b0),
    .i1(arb2_mask0[3]),
    .sel(\u_ITCM_CTRL/n0 ),
    .o(\u_ITCM_CTRL/bram_wea [3]));  // ../RTL/periph/bram2rib.v(98)
  and \u_ITCM_CTRL/u2  (\u_ITCM_CTRL/n0 , arb2_wrcs0, arb2_req0);  // ../RTL/periph/bram2rib.v(98)
  EG_LOGIC_BRAM #(
    //.FORCE_KEEP("OFF"),
    //.INIT_FILE("../../../../EIDE/ritter mcu/mem.dat"),
    .ADDR_WIDTH_A(14),
    .ADDR_WIDTH_B(14),
    .BYTE_A(4),
    .BYTE_B(4),
    .BYTE_ENABLE(8),
    .DATA_DEPTH_A(16384),
    .DATA_DEPTH_B(16384),
    .DATA_WIDTH_A(32),
    .DATA_WIDTH_B(32),
    .DEBUGGABLE("NO"),
    .FILL_ALL("NONE"),
    .IMPLEMENT("9K(FAST)"),
    .MODE("SP"),
    .PACKABLE("NO"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst  (
    .addra(arb2_addr0[15:2]),
    .addrb(14'b00000000000000),
    .bea(\u_ITCM_CTRL/bram_wea ),
    .beb(4'b0000),
    .cea(1'b1),
    .ceb(1'b0),
    .clka(i_clk),
    .clkb(1'b0),
    .dia(arb2_wdata0),
    .dib(32'b00000000000000000000000000000000),
    .ocea(1'b0),
    .oceb(1'b0),
    .rsta(1'b0),
    .rstb(1'b0),
    .wea(1'b0),
    .web(1'b0),
    .doa(arb2_rdata0));  // al_ip/bram_itcm.v(53)
  RITTER_TOP u_RITTER_TOP (
    .i_clk(i_clk),
    .i_ribm_gnt0(arb0_gnt0),
    .i_ribm_gnt1(rib_gnt1),
    .i_ribm_rdata0(rib_rdata0),
    .i_ribm_rdata1(rib_rdata1),
    .i_ribm_rsp0(arb0_rsp0),
    .i_ribm_rsp1(rib_rsp1),
    .i_rstn(i_rstn),
    .o_ribm_addr0({rib_addr0[31:24],open_n64,open_n65,open_n66,open_n67,open_n68,open_n69,open_n70,open_n71,rib_addr0[15:2],open_n72,open_n73}),
    .o_ribm_addr1({rib_addr1[31:24],open_n74,open_n75,open_n76,open_n77,open_n78,open_n79,open_n80,open_n81,rib_addr1[15:2],open_n82,open_n83}),
    .o_ribm_mask1(rib_mask1),
    .o_ribm_req0(rib_req0),
    .o_ribm_req1(rib_req1),
    .o_ribm_wdata1(rib_wdata1),
    .o_ribm_wrcs1(rib_wrcs1));  // ../RTL/soc_top/core_top.v(59)

endmodule 

module AL_DFF_X
  (
  ar,
  as,
  clk,
  d,
  en,
  sr,
  ss,
  q
  );

  input ar;
  input as;
  input clk;
  input d;
  input en;
  input sr;
  input ss;
  output q;

  wire enout;
  wire srout;
  wire ssout;

  AL_MUX u_en (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset (
    .i0(ssout),
    .i1(1'b0),
    .sel(sr),
    .o(srout));
  AL_DFF u_seq (
    .clk(clk),
    .d(srout),
    .reset(ar),
    .set(as),
    .q(q));
  AL_MUX u_set (
    .i0(enout),
    .i1(1'b1),
    .sel(ss),
    .o(ssout));

endmodule 

module eq_w8
  (
  i0,
  i1,
  o
  );

  input [7:0] i0;
  input [7:0] i1;
  output o;

  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[4]_i1[4_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;

  not none_diff (o, \or_or_or_xor_i0[0]_i_o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[4]_i1[4_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_or_xor_i0[4]_i1[4  (\or_or_xor_i0[4]_i1[4_o , \or_xor_i0[4]_i1[4]_o_o , \or_xor_i0[6]_i1[6]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \xor_i0[3]_i1[3]_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \xor_i0[7]_i1[7]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);

endmodule 

module binary_mux_s1_w1
  (
  i0,
  i1,
  sel,
  o
  );

  input i0;
  input i1;
  input sel;
  output o;


  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel),
    .o(o));

endmodule 

module add_pu64_pu64_o64
  (
  i0,
  i1,
  o
  );

  input [63:0] i0;
  input [63:0] i1;
  output [63:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a32;
  wire net_a33;
  wire net_a34;
  wire net_a35;
  wire net_a36;
  wire net_a37;
  wire net_a38;
  wire net_a39;
  wire net_a4;
  wire net_a40;
  wire net_a41;
  wire net_a42;
  wire net_a43;
  wire net_a44;
  wire net_a45;
  wire net_a46;
  wire net_a47;
  wire net_a48;
  wire net_a49;
  wire net_a5;
  wire net_a50;
  wire net_a51;
  wire net_a52;
  wire net_a53;
  wire net_a54;
  wire net_a55;
  wire net_a56;
  wire net_a57;
  wire net_a58;
  wire net_a59;
  wire net_a6;
  wire net_a60;
  wire net_a61;
  wire net_a62;
  wire net_a63;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b32;
  wire net_b33;
  wire net_b34;
  wire net_b35;
  wire net_b36;
  wire net_b37;
  wire net_b38;
  wire net_b39;
  wire net_b4;
  wire net_b40;
  wire net_b41;
  wire net_b42;
  wire net_b43;
  wire net_b44;
  wire net_b45;
  wire net_b46;
  wire net_b47;
  wire net_b48;
  wire net_b49;
  wire net_b5;
  wire net_b50;
  wire net_b51;
  wire net_b52;
  wire net_b53;
  wire net_b54;
  wire net_b55;
  wire net_b56;
  wire net_b57;
  wire net_b58;
  wire net_b59;
  wire net_b6;
  wire net_b60;
  wire net_b61;
  wire net_b62;
  wire net_b63;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout32;
  wire net_cout33;
  wire net_cout34;
  wire net_cout35;
  wire net_cout36;
  wire net_cout37;
  wire net_cout38;
  wire net_cout39;
  wire net_cout4;
  wire net_cout40;
  wire net_cout41;
  wire net_cout42;
  wire net_cout43;
  wire net_cout44;
  wire net_cout45;
  wire net_cout46;
  wire net_cout47;
  wire net_cout48;
  wire net_cout49;
  wire net_cout5;
  wire net_cout50;
  wire net_cout51;
  wire net_cout52;
  wire net_cout53;
  wire net_cout54;
  wire net_cout55;
  wire net_cout56;
  wire net_cout57;
  wire net_cout58;
  wire net_cout59;
  wire net_cout6;
  wire net_cout60;
  wire net_cout61;
  wire net_cout62;
  wire net_cout63;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum32;
  wire net_sum33;
  wire net_sum34;
  wire net_sum35;
  wire net_sum36;
  wire net_sum37;
  wire net_sum38;
  wire net_sum39;
  wire net_sum4;
  wire net_sum40;
  wire net_sum41;
  wire net_sum42;
  wire net_sum43;
  wire net_sum44;
  wire net_sum45;
  wire net_sum46;
  wire net_sum47;
  wire net_sum48;
  wire net_sum49;
  wire net_sum5;
  wire net_sum50;
  wire net_sum51;
  wire net_sum52;
  wire net_sum53;
  wire net_sum54;
  wire net_sum55;
  wire net_sum56;
  wire net_sum57;
  wire net_sum58;
  wire net_sum59;
  wire net_sum6;
  wire net_sum60;
  wire net_sum61;
  wire net_sum62;
  wire net_sum63;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a63 = i0[63];
  assign net_a62 = i0[62];
  assign net_a61 = i0[61];
  assign net_a60 = i0[60];
  assign net_a59 = i0[59];
  assign net_a58 = i0[58];
  assign net_a57 = i0[57];
  assign net_a56 = i0[56];
  assign net_a55 = i0[55];
  assign net_a54 = i0[54];
  assign net_a53 = i0[53];
  assign net_a52 = i0[52];
  assign net_a51 = i0[51];
  assign net_a50 = i0[50];
  assign net_a49 = i0[49];
  assign net_a48 = i0[48];
  assign net_a47 = i0[47];
  assign net_a46 = i0[46];
  assign net_a45 = i0[45];
  assign net_a44 = i0[44];
  assign net_a43 = i0[43];
  assign net_a42 = i0[42];
  assign net_a41 = i0[41];
  assign net_a40 = i0[40];
  assign net_a39 = i0[39];
  assign net_a38 = i0[38];
  assign net_a37 = i0[37];
  assign net_a36 = i0[36];
  assign net_a35 = i0[35];
  assign net_a34 = i0[34];
  assign net_a33 = i0[33];
  assign net_a32 = i0[32];
  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b63 = i1[63];
  assign net_b62 = i1[62];
  assign net_b61 = i1[61];
  assign net_b60 = i1[60];
  assign net_b59 = i1[59];
  assign net_b58 = i1[58];
  assign net_b57 = i1[57];
  assign net_b56 = i1[56];
  assign net_b55 = i1[55];
  assign net_b54 = i1[54];
  assign net_b53 = i1[53];
  assign net_b52 = i1[52];
  assign net_b51 = i1[51];
  assign net_b50 = i1[50];
  assign net_b49 = i1[49];
  assign net_b48 = i1[48];
  assign net_b47 = i1[47];
  assign net_b46 = i1[46];
  assign net_b45 = i1[45];
  assign net_b44 = i1[44];
  assign net_b43 = i1[43];
  assign net_b42 = i1[42];
  assign net_b41 = i1[41];
  assign net_b40 = i1[40];
  assign net_b39 = i1[39];
  assign net_b38 = i1[38];
  assign net_b37 = i1[37];
  assign net_b36 = i1[36];
  assign net_b35 = i1[35];
  assign net_b34 = i1[34];
  assign net_b33 = i1[33];
  assign net_b32 = i1[32];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[63] = net_sum63;
  assign o[62] = net_sum62;
  assign o[61] = net_sum61;
  assign o[60] = net_sum60;
  assign o[59] = net_sum59;
  assign o[58] = net_sum58;
  assign o[57] = net_sum57;
  assign o[56] = net_sum56;
  assign o[55] = net_sum55;
  assign o[54] = net_sum54;
  assign o[53] = net_sum53;
  assign o[52] = net_sum52;
  assign o[51] = net_sum51;
  assign o[50] = net_sum50;
  assign o[49] = net_sum49;
  assign o[48] = net_sum48;
  assign o[47] = net_sum47;
  assign o[46] = net_sum46;
  assign o[45] = net_sum45;
  assign o[44] = net_sum44;
  assign o[43] = net_sum43;
  assign o[42] = net_sum42;
  assign o[41] = net_sum41;
  assign o[40] = net_sum40;
  assign o[39] = net_sum39;
  assign o[38] = net_sum38;
  assign o[37] = net_sum37;
  assign o[36] = net_sum36;
  assign o[35] = net_sum35;
  assign o[34] = net_sum34;
  assign o[33] = net_sum33;
  assign o[32] = net_sum32;
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_32 (
    .a(net_a32),
    .b(net_b32),
    .c(net_cout31),
    .cout(net_cout32),
    .sum(net_sum32));
  AL_FADD comp_33 (
    .a(net_a33),
    .b(net_b33),
    .c(net_cout32),
    .cout(net_cout33),
    .sum(net_sum33));
  AL_FADD comp_34 (
    .a(net_a34),
    .b(net_b34),
    .c(net_cout33),
    .cout(net_cout34),
    .sum(net_sum34));
  AL_FADD comp_35 (
    .a(net_a35),
    .b(net_b35),
    .c(net_cout34),
    .cout(net_cout35),
    .sum(net_sum35));
  AL_FADD comp_36 (
    .a(net_a36),
    .b(net_b36),
    .c(net_cout35),
    .cout(net_cout36),
    .sum(net_sum36));
  AL_FADD comp_37 (
    .a(net_a37),
    .b(net_b37),
    .c(net_cout36),
    .cout(net_cout37),
    .sum(net_sum37));
  AL_FADD comp_38 (
    .a(net_a38),
    .b(net_b38),
    .c(net_cout37),
    .cout(net_cout38),
    .sum(net_sum38));
  AL_FADD comp_39 (
    .a(net_a39),
    .b(net_b39),
    .c(net_cout38),
    .cout(net_cout39),
    .sum(net_sum39));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_40 (
    .a(net_a40),
    .b(net_b40),
    .c(net_cout39),
    .cout(net_cout40),
    .sum(net_sum40));
  AL_FADD comp_41 (
    .a(net_a41),
    .b(net_b41),
    .c(net_cout40),
    .cout(net_cout41),
    .sum(net_sum41));
  AL_FADD comp_42 (
    .a(net_a42),
    .b(net_b42),
    .c(net_cout41),
    .cout(net_cout42),
    .sum(net_sum42));
  AL_FADD comp_43 (
    .a(net_a43),
    .b(net_b43),
    .c(net_cout42),
    .cout(net_cout43),
    .sum(net_sum43));
  AL_FADD comp_44 (
    .a(net_a44),
    .b(net_b44),
    .c(net_cout43),
    .cout(net_cout44),
    .sum(net_sum44));
  AL_FADD comp_45 (
    .a(net_a45),
    .b(net_b45),
    .c(net_cout44),
    .cout(net_cout45),
    .sum(net_sum45));
  AL_FADD comp_46 (
    .a(net_a46),
    .b(net_b46),
    .c(net_cout45),
    .cout(net_cout46),
    .sum(net_sum46));
  AL_FADD comp_47 (
    .a(net_a47),
    .b(net_b47),
    .c(net_cout46),
    .cout(net_cout47),
    .sum(net_sum47));
  AL_FADD comp_48 (
    .a(net_a48),
    .b(net_b48),
    .c(net_cout47),
    .cout(net_cout48),
    .sum(net_sum48));
  AL_FADD comp_49 (
    .a(net_a49),
    .b(net_b49),
    .c(net_cout48),
    .cout(net_cout49),
    .sum(net_sum49));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_50 (
    .a(net_a50),
    .b(net_b50),
    .c(net_cout49),
    .cout(net_cout50),
    .sum(net_sum50));
  AL_FADD comp_51 (
    .a(net_a51),
    .b(net_b51),
    .c(net_cout50),
    .cout(net_cout51),
    .sum(net_sum51));
  AL_FADD comp_52 (
    .a(net_a52),
    .b(net_b52),
    .c(net_cout51),
    .cout(net_cout52),
    .sum(net_sum52));
  AL_FADD comp_53 (
    .a(net_a53),
    .b(net_b53),
    .c(net_cout52),
    .cout(net_cout53),
    .sum(net_sum53));
  AL_FADD comp_54 (
    .a(net_a54),
    .b(net_b54),
    .c(net_cout53),
    .cout(net_cout54),
    .sum(net_sum54));
  AL_FADD comp_55 (
    .a(net_a55),
    .b(net_b55),
    .c(net_cout54),
    .cout(net_cout55),
    .sum(net_sum55));
  AL_FADD comp_56 (
    .a(net_a56),
    .b(net_b56),
    .c(net_cout55),
    .cout(net_cout56),
    .sum(net_sum56));
  AL_FADD comp_57 (
    .a(net_a57),
    .b(net_b57),
    .c(net_cout56),
    .cout(net_cout57),
    .sum(net_sum57));
  AL_FADD comp_58 (
    .a(net_a58),
    .b(net_b58),
    .c(net_cout57),
    .cout(net_cout58),
    .sum(net_sum58));
  AL_FADD comp_59 (
    .a(net_a59),
    .b(net_b59),
    .c(net_cout58),
    .cout(net_cout59),
    .sum(net_sum59));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_60 (
    .a(net_a60),
    .b(net_b60),
    .c(net_cout59),
    .cout(net_cout60),
    .sum(net_sum60));
  AL_FADD comp_61 (
    .a(net_a61),
    .b(net_b61),
    .c(net_cout60),
    .cout(net_cout61),
    .sum(net_sum61));
  AL_FADD comp_62 (
    .a(net_a62),
    .b(net_b62),
    .c(net_cout61),
    .cout(net_cout62),
    .sum(net_sum62));
  AL_FADD comp_63 (
    .a(net_a63),
    .b(net_b63),
    .c(net_cout62),
    .cout(net_cout63),
    .sum(net_sum63));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module eq_w16
  (
  i0,
  i1,
  o
  );

  input [15:0] i0;
  input [15:0] i1;
  output o;

  wire \or_or_or_or_xor_i0[0_o ;
  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_or_xor_i0[8]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[12]_i1[_o ;
  wire \or_or_xor_i0[4]_i1[4_o ;
  wire \or_or_xor_i0[8]_i1[8_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[10]_i1[10]_o ;
  wire \or_xor_i0[12]_i1[12]_o ;
  wire \or_xor_i0[14]_i1[14]_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[8]_i1[8]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[12]_i1[12]_o ;
  wire \xor_i0[13]_i1[13]_o ;
  wire \xor_i0[14]_i1[14]_o ;
  wire \xor_i0[15]_i1[15]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, \or_or_or_or_xor_i0[0_o );
  or \or_or_or_or_xor_i0[0  (\or_or_or_or_xor_i0[0_o , \or_or_or_xor_i0[0]_i_o , \or_or_or_xor_i0[8]_i_o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[4]_i1[4_o );
  or \or_or_or_xor_i0[8]_i  (\or_or_or_xor_i0[8]_i_o , \or_or_xor_i0[8]_i1[8_o , \or_or_xor_i0[12]_i1[_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_or_xor_i0[12]_i1[  (\or_or_xor_i0[12]_i1[_o , \or_xor_i0[12]_i1[12]_o , \or_xor_i0[14]_i1[14]_o );
  or \or_or_xor_i0[4]_i1[4  (\or_or_xor_i0[4]_i1[4_o , \or_xor_i0[4]_i1[4]_o_o , \or_xor_i0[6]_i1[6]_o_o );
  or \or_or_xor_i0[8]_i1[8  (\or_or_xor_i0[8]_i1[8_o , \or_xor_i0[8]_i1[8]_o_o , \or_xor_i0[10]_i1[10]_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[10]_i1[10]  (\or_xor_i0[10]_i1[10]_o , \xor_i0[10]_i1[10]_o , \xor_i0[11]_i1[11]_o );
  or \or_xor_i0[12]_i1[12]  (\or_xor_i0[12]_i1[12]_o , \xor_i0[12]_i1[12]_o , \xor_i0[13]_i1[13]_o );
  or \or_xor_i0[14]_i1[14]  (\or_xor_i0[14]_i1[14]_o , \xor_i0[14]_i1[14]_o , \xor_i0[15]_i1[15]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \xor_i0[3]_i1[3]_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \xor_i0[7]_i1[7]_o );
  or \or_xor_i0[8]_i1[8]_o  (\or_xor_i0[8]_i1[8]_o_o , \xor_i0[8]_i1[8]_o , \xor_i0[9]_i1[9]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (\xor_i0[12]_i1[12]_o , i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (\xor_i0[13]_i1[13]_o , i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (\xor_i0[14]_i1[14]_o , i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (\xor_i0[15]_i1[15]_o , i0[15], i1[15]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module binary_mux_s4_w1
  (
  i0,
  i1,
  i10,
  i11,
  i12,
  i13,
  i14,
  i15,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  sel,
  o
  );

  input i0;
  input i1;
  input i10;
  input i11;
  input i12;
  input i13;
  input i14;
  input i15;
  input i2;
  input i3;
  input i4;
  input i5;
  input i6;
  input i7;
  input i8;
  input i9;
  input [3:0] sel;
  output o;

  wire  B0_0;
  wire  B0_1;
  wire  B0_2;
  wire  B0_3;
  wire  B0_4;
  wire  B0_5;
  wire  B0_6;
  wire  B0_7;
  wire  B1_0;
  wire  B1_1;
  wire  B1_2;
  wire  B1_3;
  wire  B2_0;
  wire  B2_1;

  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel[0]),
    .o(B0_0));
  AL_MUX al_mux_b0_0_1 (
    .i0(i2),
    .i1(i3),
    .sel(sel[0]),
    .o(B0_1));
  AL_MUX al_mux_b0_0_2 (
    .i0(i4),
    .i1(i5),
    .sel(sel[0]),
    .o(B0_2));
  AL_MUX al_mux_b0_0_3 (
    .i0(i6),
    .i1(i7),
    .sel(sel[0]),
    .o(B0_3));
  AL_MUX al_mux_b0_0_4 (
    .i0(i8),
    .i1(i9),
    .sel(sel[0]),
    .o(B0_4));
  AL_MUX al_mux_b0_0_5 (
    .i0(i10),
    .i1(i11),
    .sel(sel[0]),
    .o(B0_5));
  AL_MUX al_mux_b0_0_6 (
    .i0(i12),
    .i1(i13),
    .sel(sel[0]),
    .o(B0_6));
  AL_MUX al_mux_b0_0_7 (
    .i0(i14),
    .i1(i15),
    .sel(sel[0]),
    .o(B0_7));
  AL_MUX al_mux_b0_1_0 (
    .i0(B0_0),
    .i1(B0_1),
    .sel(sel[1]),
    .o(B1_0));
  AL_MUX al_mux_b0_1_1 (
    .i0(B0_2),
    .i1(B0_3),
    .sel(sel[1]),
    .o(B1_1));
  AL_MUX al_mux_b0_1_2 (
    .i0(B0_4),
    .i1(B0_5),
    .sel(sel[1]),
    .o(B1_2));
  AL_MUX al_mux_b0_1_3 (
    .i0(B0_6),
    .i1(B0_7),
    .sel(sel[1]),
    .o(B1_3));
  AL_MUX al_mux_b0_2_0 (
    .i0(B1_0),
    .i1(B1_1),
    .sel(sel[2]),
    .o(B2_0));
  AL_MUX al_mux_b0_2_1 (
    .i0(B1_2),
    .i1(B1_3),
    .sel(sel[2]),
    .o(B2_1));
  AL_MUX al_mux_b0_3_0 (
    .i0(B2_0),
    .i1(B2_1),
    .sel(sel[3]),
    .o(o));

endmodule 

module AL_DFF_0
  (
  ar,
  as,
  clk,
  d,
  en,
  sr,
  ss,
  q
  );

  input ar;
  input as;
  input clk;
  input d;
  input en;
  input sr;
  input ss;
  output q;

  wire enout;
  wire srout;
  wire ssout;

  AL_MUX u_en (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset (
    .i0(ssout),
    .i1(1'b0),
    .sel(sr),
    .o(srout));
  AL_DFF #(
    .INI(1'b0))
    u_seq (
    .clk(clk),
    .d(srout),
    .reset(ar),
    .set(as),
    .q(q));
  AL_MUX u_set (
    .i0(enout),
    .i1(1'b1),
    .sel(ss),
    .o(ssout));

endmodule 

module AL_LATCH_X
  (
  ar,
  as,
  clk,
  d,
  en,
  sr,
  ss,
  q
  );

  input ar;
  input as;
  input clk;
  input d;
  input en;
  input sr;
  input ss;
  output q;

  wire enout;
  wire srout;
  wire ssout;

  AL_MUX u_en (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset (
    .i0(ssout),
    .i1(1'b0),
    .sel(sr),
    .o(srout));
  AL_LATCH u_seq (
    .clk(clk),
    .d(srout),
    .reset(ar),
    .set(as),
    .q(q));
  AL_MUX u_set (
    .i0(enout),
    .i1(1'b1),
    .sel(ss),
    .o(ssout));

endmodule 

module binary_mux_s2_w1
  (
  i0,
  i1,
  i2,
  i3,
  sel,
  o
  );

  input i0;
  input i1;
  input i2;
  input i3;
  input [1:0] sel;
  output o;

  wire  B0_0;
  wire  B0_1;

  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel[0]),
    .o(B0_0));
  AL_MUX al_mux_b0_0_1 (
    .i0(i2),
    .i1(i3),
    .sel(sel[0]),
    .o(B0_1));
  AL_MUX al_mux_b0_1_0 (
    .i0(B0_0),
    .i1(B0_1),
    .sel(sel[1]),
    .o(o));

endmodule 

module eq_w1
  (
  i0,
  i1,
  o
  );

  input i0;
  input i1;
  output o;

  wire xor_i0_i1_o;

  not none_diff (o, xor_i0_i1_o);
  xor xor_i0_i1 (xor_i0_i1_o, i0, i1);

endmodule 

module RITTER_TOP  // ../RTL/core/ritter_top.v(6)
  (
  i_clk,
  i_ribm_gnt0,
  i_ribm_gnt1,
  i_ribm_rdata0,
  i_ribm_rdata1,
  i_ribm_rsp0,
  i_ribm_rsp1,
  i_rstn,
  o_ribm_addr0,
  o_ribm_addr1,
  o_ribm_mask0,
  o_ribm_mask1,
  o_ribm_rdy0,
  o_ribm_rdy1,
  o_ribm_req0,
  o_ribm_req1,
  o_ribm_wdata0,
  o_ribm_wdata1,
  o_ribm_wrcs0,
  o_ribm_wrcs1
  );

  input i_clk;  // ../RTL/core/ritter_top.v(7)
  input i_ribm_gnt0;  // ../RTL/core/ritter_top.v(17)
  input i_ribm_gnt1;  // ../RTL/core/ritter_top.v(27)
  input [31:0] i_ribm_rdata0;  // ../RTL/core/ritter_top.v(15)
  input [31:0] i_ribm_rdata1;  // ../RTL/core/ritter_top.v(25)
  input i_ribm_rsp0;  // ../RTL/core/ritter_top.v(18)
  input i_ribm_rsp1;  // ../RTL/core/ritter_top.v(28)
  input i_rstn;  // ../RTL/core/ritter_top.v(8)
  output [31:0] o_ribm_addr0;  // ../RTL/core/ritter_top.v(11)
  output [31:0] o_ribm_addr1;  // ../RTL/core/ritter_top.v(21)
  output [3:0] o_ribm_mask0;  // ../RTL/core/ritter_top.v(13)
  output [3:0] o_ribm_mask1;  // ../RTL/core/ritter_top.v(23)
  output o_ribm_rdy0;  // ../RTL/core/ritter_top.v(19)
  output o_ribm_rdy1;  // ../RTL/core/ritter_top.v(29)
  output o_ribm_req0;  // ../RTL/core/ritter_top.v(16)
  output o_ribm_req1;  // ../RTL/core/ritter_top.v(26)
  output [31:0] o_ribm_wdata0;  // ../RTL/core/ritter_top.v(14)
  output [31:0] o_ribm_wdata1;  // ../RTL/core/ritter_top.v(24)
  output o_ribm_wrcs0;  // ../RTL/core/ritter_top.v(12)
  output o_ribm_wrcs1;  // ../RTL/core/ritter_top.v(22)

  wire [31:0] bpu_csr_zimm;  // ../RTL/core/ritter_top.v(153)
  wire [11:0] bpu_csridx;  // ../RTL/core/ritter_top.v(151)
  wire [9:0] bpu_decinfo;  // ../RTL/core/ritter_top.v(155)
  wire [5:0] bpu_decinfo_grp;  // ../RTL/core/ritter_top.v(154)
  wire [31:0] bpu_exu_op1;  // ../RTL/core/ritter_top.v(143)
  wire [31:0] bpu_exu_op2;  // ../RTL/core/ritter_top.v(144)
  wire [31:0] bpu_iaddr;  // ../RTL/core/ritter_top.v(156)
  wire [31:0] bpu_imm;  // ../RTL/core/ritter_top.v(146)
  wire [31:0] bpu_jaddr;  // ../RTL/core/ritter_top.v(141)
  wire [31:0] bpu_jaddr_gen;  // ../RTL/core/ritter_top.v(79)
  wire [4:0] bpu_rdidx;  // ../RTL/core/ritter_top.v(148)
  wire [31:0] bpu_rs2rdata;  // ../RTL/core/ritter_top.v(145)
  wire [31:0] csr_rdata;  // ../RTL/core/ritter_top.v(200)
  wire [4:0] ctrl2bpu_rs1idx;  // ../RTL/core/ritter_top.v(34)
  wire [4:0] ctrl2bpu_rs2idx;  // ../RTL/core/ritter_top.v(36)
  wire [4:0] ctrl2exu_rdidx0;  // ../RTL/core/ritter_top.v(39)
  wire [4:0] ctrl2exu_rdidx1;  // ../RTL/core/ritter_top.v(42)
  wire [4:0] ctrl2exu_rdidx2;  // ../RTL/core/ritter_top.v(44)
  wire [31:0] dis_csr_rdata;  // ../RTL/core/ritter_top.v(230)
  wire [31:0] dis_csr_zimm;  // ../RTL/core/ritter_top.v(231)
  wire [11:0] dis_csridx;  // ../RTL/core/ritter_top.v(229)
  wire [9:0] dis_decinfo;  // ../RTL/core/ritter_top.v(234)
  wire [5:0] dis_decinfo_grp;  // ../RTL/core/ritter_top.v(233)
  wire [31:0] dis_exu_op1;  // ../RTL/core/ritter_top.v(222)
  wire [31:0] dis_exu_op2;  // ../RTL/core/ritter_top.v(223)
  wire [31:0] dis_iaddr;  // ../RTL/core/ritter_top.v(235)
  wire [31:0] dis_imm;  // ../RTL/core/ritter_top.v(225)
  wire [4:0] dis_rdidx;  // ../RTL/core/ritter_top.v(227)
  wire [31:0] dis_rs2rdata;  // ../RTL/core/ritter_top.v(224)
  wire [31:0] exu_jaddr;  // ../RTL/core/ritter_top.v(296)
  wire [31:0] exu_jaddr_gen;  // ../RTL/core/ritter_top.v(81)
  wire [4:0] exu_rdidx0;  // ../RTL/core/ritter_top.v(284)
  wire [4:0] exu_rdidx1;  // ../RTL/core/ritter_top.v(288)
  wire [4:0] exu_rdidx2;  // ../RTL/core/ritter_top.v(292)
  wire [31:0] exu_rdwdata0;  // ../RTL/core/ritter_top.v(285)
  wire [31:0] exu_rdwdata1;  // ../RTL/core/ritter_top.v(289)
  wire [31:0] exu_rdwdata2;  // ../RTL/core/ritter_top.v(293)
  wire [31:0] ifu2bpu_data;  // ../RTL/core/ritter_top.v(117)
  wire [31:0] ifu2bpu_iaddr;  // ../RTL/core/ritter_top.v(116)
  wire [31:0] ifu_iaddr;  // ../RTL/core/ritter_top.v(83)
  wire [5:0] \u_DISPATCH/n5 ;
  wire [31:0] \u_IFU/fetch_addr ;  // ../RTL/core/ifu.v(80)
  wire [0:0] \u_IFU/fifo_cnt ;  // ../RTL/core/ifu.v(130)
  wire [31:0] \u_IFU/jump_addr ;  // ../RTL/core/ifu.v(62)
  wire [0:0] \u_IFU/u_IFU_FIFO/hptr ;  // ../RTL/core/fifos.v(120)
  wire [0:0] \u_IFU/u_IFU_FIFO/hptr_1 ;  // ../RTL/core/fifos.v(124)
  wire [0:0] \u_IFU/u_IFU_FIFO/n10 ;
  wire [1:0] \u_IFU/u_IFU_FIFO/n11 ;
  wire [0:0] \u_IFU/u_IFU_FIFO/n2 ;
  wire [31:0] \u_IFU/u_IFU_PC/n10 ;
  wire [29:0] \u_IFU/u_IFU_PC/n2 ;
  wire [29:0] \u_IFU/u_IFU_PC/n3 ;
  wire [29:0] \u_IFU/u_IFU_PC/n4 ;
  wire [31:0] \u_IFU/u_IFU_PC/n5 ;
  wire [31:0] \u_IFU/u_IFU_PC/n9 ;
  wire [31:0] \u_IFU/u_IFU_PC/pc ;  // ../RTL/core/ifu_pc.v(23)
  wire [8:0] \u_IFU2BPU/fifo_cnt ;  // ../RTL/core/ifu2bpu.v(37)
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/eptr ;  // ../RTL/core/fifos.v(36)
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/eptr_1 ;  // ../RTL/core/fifos.v(42)
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/hptr ;  // ../RTL/core/fifos.v(36)
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/hptr_1 ;  // ../RTL/core/fifos.v(40)
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n10 ;
  wire [4:0] \u_IFU2BPU/u_SYNC_FIFO/n13 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n14 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n15 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n16 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n2 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n20 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n21 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n22 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n23 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n24 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n5 ;
  wire [31:0] \u_PIPE_CTRL/n1 ;
  wire [31:0] \u_PIPE_CTRL/n11 ;
  wire [31:0] \u_PIPE_CTRL/n12 ;
  wire [31:0] \u_PIPE_CTRL/n14 ;
  wire [31:0] \u_PIPE_CTRL/n15 ;
  wire [31:0] \u_PIPE_CTRL/n3 ;
  wire [31:0] \u_PIPE_CTRL/n4 ;
  wire [31:0] \u_PIPE_CTRL/n6 ;
  wire [31:0] \u_PIPE_CTRL/n7 ;
  wire [31:0] \u_PIPE_CTRL/n9 ;
  wire [4:0] \u_WB/n34 ;
  wire [31:0] \u_WB/n35 ;
  wire [4:0] \u_WB/rdidx0 ;  // ../RTL/core/wb.v(48)
  wire [4:0] \u_WB/rdidx1 ;  // ../RTL/core/wb.v(49)
  wire [4:0] \u_WB/rdidx2 ;  // ../RTL/core/wb.v(50)
  wire [31:0] \u_WB/rdwdata0 ;  // ../RTL/core/wb.v(51)
  wire [31:0] \u_WB/rdwdata1 ;  // ../RTL/core/wb.v(52)
  wire [31:0] \u_WB/rdwdata2 ;  // ../RTL/core/wb.v(53)
  wire [31:0] wb_csr_wdata;  // ../RTL/core/ritter_top.v(204)
  wire [11:0] wb_csridx;  // ../RTL/core/ritter_top.v(203)
  wire [4:0] wb_rdidx;  // ../RTL/core/ritter_top.v(137)
  wire [31:0] wb_rdwdata;  // ../RTL/core/ritter_top.v(138)
  wire bpu2ifu_vld;  // ../RTL/core/ritter_top.v(86)
  wire bpu_csrwren;  // ../RTL/core/ritter_top.v(150)
  wire bpu_inst_vld;  // ../RTL/core/ritter_top.v(142)
  wire bpu_rdwen;  // ../RTL/core/ritter_top.v(147)
  wire bpu_taken;  // ../RTL/core/ritter_top.v(140)
  wire bpu_taken_gen;  // ../RTL/core/ritter_top.v(78)
  wire ctrl2bpu_rs1ren;  // ../RTL/core/ritter_top.v(33)
  wire ctrl2bpu_rs2ren;  // ../RTL/core/ritter_top.v(35)
  wire ctrl2bpu_wait;  // ../RTL/core/ritter_top.v(50)
  wire ctrl2dis_flush;  // ../RTL/core/ritter_top.v(52)
  wire ctrl2dis_wait;  // ../RTL/core/ritter_top.v(51)
  wire ctrl2exu_rdwen0;  // ../RTL/core/ritter_top.v(38)
  wire ctrl2exu_rdwen1;  // ../RTL/core/ritter_top.v(41)
  wire ctrl2exu_rdwen2;  // ../RTL/core/ritter_top.v(43)
  wire ctrl2exu_resource_match;  // ../RTL/core/ritter_top.v(46)
  wire ctrl2wb_match;  // ../RTL/core/ritter_top.v(47)
  wire dis_rdwen;  // ../RTL/core/ritter_top.v(226)
  wire exu_rdwen0;  // ../RTL/core/ritter_top.v(283)
  wire exu_rdwen1;  // ../RTL/core/ritter_top.v(287)
  wire exu_rdwen2;  // ../RTL/core/ritter_top.v(291)
  wire exu_taken;  // ../RTL/core/ritter_top.v(295)
  wire exu_taken_gen;  // ../RTL/core/ritter_top.v(80)
  wire ifu2bpu_data_vld;  // ../RTL/core/ritter_top.v(115)
  wire ifu_data_vld;  // ../RTL/core/ritter_top.v(82)
  wire ifu_fetch_vld;  // ../RTL/core/ritter_top.v(88)
  wire n0;
  wire n0_neg;
  wire n1;
  wire n2;
  wire n3;
  wire n4;
  wire n5;
  wire \u_DISPATCH/mux12_b0_sel_is_2_o ;
  wire \u_DISPATCH/n1 ;
  wire \u_DISPATCH/n2 ;
  wire \u_DISPATCH/n28 ;
  wire \u_DISPATCH/n3 ;
  wire \u_DISPATCH/n4 ;
  wire \u_IFU/data_vld ;  // ../RTL/core/ifu.v(79)
  wire \u_IFU/jump_flag ;  // ../RTL/core/ifu.v(61)
  wire \u_IFU/n0 ;
  wire \u_IFU/pc_vld ;  // ../RTL/core/ifu.v(77)
  wire \u_IFU/u_IFU_FETCH/handshake_rdy_last ;  // ../RTL/core/ifu_fetch.v(70)
  wire \u_IFU/u_IFU_FETCH/n1 ;
  wire \u_IFU/u_IFU_FETCH/n2 ;
  wire \u_IFU/u_IFU_FETCH/n2_neg ;
  wire \u_IFU/u_IFU_FETCH/n3 ;
  wire \u_IFU/u_IFU_FETCH/n4 ;
  wire \u_IFU/u_IFU_FETCH/n5 ;
  wire \u_IFU/u_IFU_FETCH/n7 ;
  wire \u_IFU/u_IFU_FETCH/u20_sel_is_2_o ;
  wire \u_IFU/u_IFU_FIFO/hptr[0]_neg ;
  wire \u_IFU/u_IFU_FIFO/mux4_b32_sel_is_1_o ;
  wire \u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ;
  wire \u_IFU/u_IFU_FIFO/n12 ;
  wire \u_IFU/u_IFU_FIFO/n13 ;
  wire \u_IFU/u_IFU_FIFO/n9 ;
  wire \u_IFU/u_IFU_PC/n1 ;
  wire \u_IFU/u_IFU_PC/n7 ;
  wire \u_IFU/u_IFU_PC/n8 ;
  wire \u_IFU2BPU/fifo_empty ;  // ../RTL/core/ifu2bpu.v(35)
  wire \u_IFU2BPU/fifo_full ;  // ../RTL/core/ifu2bpu.v(34)
  wire \u_IFU2BPU/n0 ;
  wire \u_IFU2BPU/n2 ;
  wire \u_IFU2BPU/u_SYNC_FIFO/n0 ;
  wire \u_IFU2BPU/u_SYNC_FIFO/n12 ;
  wire \u_IFU2BPU/u_SYNC_FIFO/n17 ;
  wire \u_IFU2BPU/u_SYNC_FIFO/n18 ;
  wire \u_IFU2BPU/u_SYNC_FIFO/n19 ;
  wire \u_IFU2BPU/u_SYNC_FIFO/n3 ;
  wire \u_IFU2BPU/u_SYNC_FIFO/n7 ;
  wire \u_IFU2BPU/u_SYNC_FIFO/n8 ;
  wire \u_IFU2BPU/u_SYNC_FIFO/n9 ;
  wire \u_IFU2BPU/u_SYNC_FIFO/u11_sel_is_0_o ;
  wire \u_PIPE_CTRL/n0 ;
  wire \u_PIPE_CTRL/n10 ;
  wire \u_PIPE_CTRL/n13 ;
  wire \u_PIPE_CTRL/n16 ;
  wire \u_PIPE_CTRL/n2 ;
  wire \u_PIPE_CTRL/n5 ;
  wire \u_PIPE_CTRL/n8 ;
  wire \u_PIPE_CTRL/read_after_write ;  // ../RTL/core/pipe_ctrl.v(51)
  wire \u_PIPE_CTRL/rs1_match ;  // ../RTL/core/pipe_ctrl.v(41)
  wire \u_PIPE_CTRL/rs2_match ;  // ../RTL/core/pipe_ctrl.v(45)
  wire \u_WB/mux10_b0_sel_is_2_o ;
  wire \u_WB/n0 ;
  wire \u_WB/n1 ;
  wire \u_WB/n12 ;
  wire \u_WB/n13 ;
  wire \u_WB/n15 ;
  wire \u_WB/n16 ;
  wire \u_WB/n2 ;
  wire \u_WB/n29 ;
  wire \u_WB/n3 ;
  wire \u_WB/n30 ;
  wire \u_WB/n31 ;
  wire \u_WB/n32 ;
  wire \u_WB/n33 ;
  wire \u_WB/n37 ;
  wire \u_WB/n4 ;
  wire \u_WB/n5 ;
  wire \u_WB/n6 ;
  wire \u_WB/n7 ;
  wire \u_WB/n8 ;
  wire \u_WB/rdwen0 ;  // ../RTL/core/wb.v(45)
  wire \u_WB/rdwen1 ;  // ../RTL/core/wb.v(46)
  wire \u_WB/rdwen2 ;  // ../RTL/core/wb.v(47)
  wire \u_WB/rdwen2_neg ;
  wire \u_WB/u13_sel_is_2_o ;
  wire \u_WB/u14_sel_is_3_o ;
  wire \u_WB/u15_sel_is_3_o ;
  wire wb_csr_wen;  // ../RTL/core/ritter_top.v(202)
  wire wb_rdwen;  // ../RTL/core/ritter_top.v(136)

  assign o_ribm_addr0[1] = 1'b0;
  assign o_ribm_addr0[0] = 1'b0;
  assign o_ribm_addr1[1] = 1'b0;
  assign o_ribm_addr1[0] = 1'b0;
  assign o_ribm_mask0[3] = 1'b1;
  assign o_ribm_mask0[2] = 1'b1;
  assign o_ribm_mask0[1] = 1'b1;
  assign o_ribm_mask0[0] = 1'b1;
  assign o_ribm_rdy0 = i_ribm_rsp0;
  assign o_ribm_wdata0[31] = 1'b0;
  assign o_ribm_wdata0[30] = 1'b0;
  assign o_ribm_wdata0[29] = 1'b0;
  assign o_ribm_wdata0[28] = 1'b0;
  assign o_ribm_wdata0[27] = 1'b0;
  assign o_ribm_wdata0[26] = 1'b0;
  assign o_ribm_wdata0[25] = 1'b0;
  assign o_ribm_wdata0[24] = 1'b0;
  assign o_ribm_wdata0[23] = 1'b0;
  assign o_ribm_wdata0[22] = 1'b0;
  assign o_ribm_wdata0[21] = 1'b0;
  assign o_ribm_wdata0[20] = 1'b0;
  assign o_ribm_wdata0[19] = 1'b0;
  assign o_ribm_wdata0[18] = 1'b0;
  assign o_ribm_wdata0[17] = 1'b0;
  assign o_ribm_wdata0[16] = 1'b0;
  assign o_ribm_wdata0[15] = 1'b0;
  assign o_ribm_wdata0[14] = 1'b0;
  assign o_ribm_wdata0[13] = 1'b0;
  assign o_ribm_wdata0[12] = 1'b0;
  assign o_ribm_wdata0[11] = 1'b0;
  assign o_ribm_wdata0[10] = 1'b0;
  assign o_ribm_wdata0[9] = 1'b0;
  assign o_ribm_wdata0[8] = 1'b0;
  assign o_ribm_wdata0[7] = 1'b0;
  assign o_ribm_wdata0[6] = 1'b0;
  assign o_ribm_wdata0[5] = 1'b0;
  assign o_ribm_wdata0[4] = 1'b0;
  assign o_ribm_wdata0[3] = 1'b0;
  assign o_ribm_wdata0[2] = 1'b0;
  assign o_ribm_wdata0[1] = 1'b0;
  assign o_ribm_wdata0[0] = 1'b0;
  assign o_ribm_wrcs0 = 1'b0;
  not n0_inv (n0_neg, n0);
  or u1 (n0, bpu_taken_gen, exu_taken_gen);  // ../RTL/core/ritter_top.v(88)
  AL_MUX u2 (
    .i0(bpu2ifu_vld),
    .i1(1'b1),
    .sel(n0),
    .o(ifu_fetch_vld));  // ../RTL/core/ritter_top.v(88)
  not u3 (n1, ctrl2bpu_wait);  // ../RTL/core/ritter_top.v(122)
  not u4 (n2, ctrl2dis_wait);  // ../RTL/core/ritter_top.v(241)
  or u5 (n3, n0, ctrl2dis_flush);  // ../RTL/core/ritter_top.v(242)
  or u6 (n4, exu_taken_gen, ctrl2dis_wait);  // ../RTL/core/ritter_top.v(301)
  not u7 (n5, n4);  // ../RTL/core/ritter_top.v(301)
  BPU u_BPU (
    .i_clk(i_clk),
    .i_data(ifu2bpu_data),
    .i_data_vld(ifu2bpu_data_vld),
    .i_flush(n0),
    .i_iaddr(ifu2bpu_iaddr),
    .i_rd_wdata(wb_rdwdata),
    .i_rdidx(wb_rdidx),
    .i_rdwen(wb_rdwen),
    .i_rstn(i_rstn),
    .i_stop(ctrl2bpu_wait),
    .o_bpu_jaddr(bpu_jaddr),
    .o_bpu_rs1idx(ctrl2bpu_rs1idx),
    .o_bpu_rs1ren(ctrl2bpu_rs1ren),
    .o_bpu_rs2idx(ctrl2bpu_rs2idx),
    .o_bpu_rs2ren(ctrl2bpu_rs2ren),
    .o_bpu_taken(bpu_taken),
    .o_csr_ren(bpu_csrwren),
    .o_csr_zimm({open_n0,open_n1,open_n2,open_n3,open_n4,open_n5,open_n6,open_n7,open_n8,open_n9,open_n10,open_n11,open_n12,open_n13,open_n14,open_n15,open_n16,open_n17,open_n18,open_n19,open_n20,open_n21,open_n22,open_n23,open_n24,open_n25,open_n26,bpu_csr_zimm[4:0]}),
    .o_csridx(bpu_csridx),
    .o_decinfo({bpu_decinfo[9:1],open_n27}),
    .o_decinfo_grp(bpu_decinfo_grp),
    .o_exu_op1(bpu_exu_op1),
    .o_exu_op2(bpu_exu_op2),
    .o_iaddr(bpu_iaddr),
    .o_imm(bpu_imm),
    .o_inst_vld(bpu_inst_vld),
    .o_rdidx(bpu_rdidx),
    .o_rdwen(bpu_rdwen),
    .o_rs2rdata(bpu_rs2rdata));  // ../RTL/core/ritter_top.v(157)
  CSR_REGFILE u_CSR_REGFILE (
    .i_clk(i_clk),
    .i_csr_ren(bpu_csrwren),
    .i_csr_ridx(bpu_csridx),
    .i_csr_wdata(wb_csr_wdata),
    .i_csr_wen(wb_csr_wen),
    .i_csr_widx(wb_csridx),
    .i_rstn(i_rstn),
    .o_csr_rdata(csr_rdata));  // ../RTL/core/ritter_top.v(206)
  binary_mux_s1_w1 \u_DISPATCH/mux0_b0  (
    .i0(bpu_decinfo_grp[0]),
    .i1(1'b0),
    .sel(\u_DISPATCH/n3 ),
    .o(\u_DISPATCH/n5 [0]));  // ../RTL/core/dispatch.v(106)
  binary_mux_s1_w1 \u_DISPATCH/mux0_b1  (
    .i0(bpu_decinfo_grp[1]),
    .i1(1'b0),
    .sel(\u_DISPATCH/n3 ),
    .o(\u_DISPATCH/n5 [1]));  // ../RTL/core/dispatch.v(106)
  binary_mux_s1_w1 \u_DISPATCH/mux0_b2  (
    .i0(bpu_decinfo_grp[2]),
    .i1(1'b0),
    .sel(\u_DISPATCH/n3 ),
    .o(\u_DISPATCH/n5 [2]));  // ../RTL/core/dispatch.v(106)
  binary_mux_s1_w1 \u_DISPATCH/mux0_b3  (
    .i0(bpu_decinfo_grp[3]),
    .i1(1'b0),
    .sel(\u_DISPATCH/n3 ),
    .o(\u_DISPATCH/n5 [3]));  // ../RTL/core/dispatch.v(106)
  binary_mux_s1_w1 \u_DISPATCH/mux0_b4  (
    .i0(bpu_decinfo_grp[4]),
    .i1(1'b0),
    .sel(\u_DISPATCH/n3 ),
    .o(\u_DISPATCH/n5 [4]));  // ../RTL/core/dispatch.v(106)
  binary_mux_s1_w1 \u_DISPATCH/mux0_b5  (
    .i0(bpu_decinfo_grp[5]),
    .i1(1'b0),
    .sel(\u_DISPATCH/n3 ),
    .o(\u_DISPATCH/n5 [5]));  // ../RTL/core/dispatch.v(106)
  and \u_DISPATCH/mux12_b0_sel_is_2  (\u_DISPATCH/mux12_b0_sel_is_2_o , i_rstn, \u_DISPATCH/n1 );
  AL_DFF_X \u_DISPATCH/o_bpu_taken_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DISPATCH/n28 ),
    .en(\u_DISPATCH/n1 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_taken_gen));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/o_rdwen_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DISPATCH/n4 ),
    .en(\u_DISPATCH/n1 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rdwen));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg0_b0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DISPATCH/n5 [0]),
    .en(\u_DISPATCH/n1 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo_grp[0]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg0_b1  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DISPATCH/n5 [1]),
    .en(\u_DISPATCH/n1 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo_grp[1]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg0_b2  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DISPATCH/n5 [2]),
    .en(\u_DISPATCH/n1 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo_grp[2]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg0_b3  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DISPATCH/n5 [3]),
    .en(\u_DISPATCH/n1 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo_grp[3]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg0_b4  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DISPATCH/n5 [4]),
    .en(\u_DISPATCH/n1 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo_grp[4]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg0_b5  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DISPATCH/n5 [5]),
    .en(\u_DISPATCH/n1 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo_grp[5]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[0]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[0]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[1]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[1]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[10]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[10]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[11]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[11]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[12]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[12]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[13]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[13]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[14]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[14]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[15]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[15]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[16]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[16]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[17]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[17]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[18]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[18]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[19]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[19]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[2]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[2]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[20]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[20]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[21]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[21]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[22]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[22]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[23]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[23]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[24]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[24]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[25]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[25]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[26]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[26]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[27]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[27]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[28]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[28]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[29]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[29]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[3]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[3]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[30]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[30]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[31]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[31]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[4]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[4]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[5]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[5]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[6]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[6]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[7]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[7]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[8]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[8]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg10_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_iaddr[9]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_iaddr[9]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg11_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[0]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[0]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[1]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[1]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[10]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[10]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[11]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[11]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[12]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[12]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[13]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[13]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[14]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[14]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[15]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[15]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[16]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[16]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[17]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[17]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[18]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[18]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[19]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[19]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[2]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[2]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[20]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[20]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[21]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[21]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[22]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[22]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[23]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[23]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[24]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[24]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[25]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[25]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[26]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[26]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[27]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[27]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[28]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[28]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[29]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[29]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[3]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[3]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[30]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[30]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[31]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[31]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[4]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[4]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[5]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[5]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[6]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[6]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[7]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[7]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[8]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[8]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg11_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_jaddr[9]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(bpu_jaddr_gen[9]));  // ../RTL/core/dispatch.v(113)
  AL_DFF_X \u_DISPATCH/reg1_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[0]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[0]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[1]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[1]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[10]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[10]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[11]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[11]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[12]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[12]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[13]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[13]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[14]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[14]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[15]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[15]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[16]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[16]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[17]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[17]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[18]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[18]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[19]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[19]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[2]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[2]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[20]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[20]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[21]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[21]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[22]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[22]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[23]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[23]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[24]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[24]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[25]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[25]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[26]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[26]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[27]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[27]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[28]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[28]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[29]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[29]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[3]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[3]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[30]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[30]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[31]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[31]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[4]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[4]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[5]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[5]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[6]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[6]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[7]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[7]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[8]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[8]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg1_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op1[9]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op1[9]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[0]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[0]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[1]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[1]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[10]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[10]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[11]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[11]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[12]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[12]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[13]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[13]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[14]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[14]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[15]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[15]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[16]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[16]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[17]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[17]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[18]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[18]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[19]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[19]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[2]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[2]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[20]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[20]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[21]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[21]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[22]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[22]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[23]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[23]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[24]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[24]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[25]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[25]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[26]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[26]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[27]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[27]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[28]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[28]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[29]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[29]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[3]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[3]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[30]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[30]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[31]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[31]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[4]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[4]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[5]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[5]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[6]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[6]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[7]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[7]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[8]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[8]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg2_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_exu_op2[9]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_exu_op2[9]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[0]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[0]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[1]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[1]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[10]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[10]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[11]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[11]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[12]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[12]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[13]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[13]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[14]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[14]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[15]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[15]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[16]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[16]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[17]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[17]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[18]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[18]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[19]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[19]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[2]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[2]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[20]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[20]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[21]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[21]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[22]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[22]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[23]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[23]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[24]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[24]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[25]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[25]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[26]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[26]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[27]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[27]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[28]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[28]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[29]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[29]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[3]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[3]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[30]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[30]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[31]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[31]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[4]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[4]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[5]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[5]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[6]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[6]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[7]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[7]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[8]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[8]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg3_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rs2rdata[9]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rs2rdata[9]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[0]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[0]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[1]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[1]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[10]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[10]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[11]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[11]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[12]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[12]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[13]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[13]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[14]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[14]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[15]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[15]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[16]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[16]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[17]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[17]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[18]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[18]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[19]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[19]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[2]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[2]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[20]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[20]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[21]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[21]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[22]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[22]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[23]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[23]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[24]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[24]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[25]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[25]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[26]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[26]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[27]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[27]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[28]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[28]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[29]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[29]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[3]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[3]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[30]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[30]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[31]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[31]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[4]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[4]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[5]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[5]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[6]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[6]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[7]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[7]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[8]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[8]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg4_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_imm[9]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_imm[9]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg5_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rdidx[0]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rdidx[0]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg5_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rdidx[1]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rdidx[1]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg5_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rdidx[2]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rdidx[2]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg5_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rdidx[3]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rdidx[3]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg5_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_rdidx[4]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_rdidx[4]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg6_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csridx[0]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csridx[0]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg6_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csridx[1]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csridx[1]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg6_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csridx[10]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csridx[10]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg6_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csridx[11]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csridx[11]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg6_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csridx[2]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csridx[2]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg6_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csridx[3]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csridx[3]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg6_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csridx[4]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csridx[4]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg6_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csridx[5]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csridx[5]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg6_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csridx[6]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csridx[6]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg6_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csridx[7]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csridx[7]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg6_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csridx[8]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csridx[8]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg6_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csridx[9]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csridx[9]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[0]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[0]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[1]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[1]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[10]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[10]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[11]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[11]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[12]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[12]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[13]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[13]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[14]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[14]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[15]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[15]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[16]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[16]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[17]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[17]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[18]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[18]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[19]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[19]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[2]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[2]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[20]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[20]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[21]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[21]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[22]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[22]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[23]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[23]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[24]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[24]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[25]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[25]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[26]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[26]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[27]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[27]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[28]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[28]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[29]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[29]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[3]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[3]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[30]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[30]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[31]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[31]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[4]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[4]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[5]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[5]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[6]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[6]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[7]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[7]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[8]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[8]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg7_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(csr_rdata[9]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_rdata[9]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csr_zimm[0]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[0]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csr_zimm[1]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[1]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[10]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[11]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[12]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[13]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[14]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[15]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[16]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[17]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[18]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[19]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csr_zimm[2]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[2]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[20]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[21]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[22]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[23]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[24]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[25]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[26]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[27]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[28]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[29]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csr_zimm[3]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[3]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[30]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[31]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_csr_zimm[4]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[4]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[5]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[6]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[7]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[8]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg8_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(1'b0),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_csr_zimm[9]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg9_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_decinfo[1]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo[1]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg9_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_decinfo[2]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo[2]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg9_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_decinfo[3]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo[3]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg9_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_decinfo[4]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo[4]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg9_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_decinfo[5]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo[5]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg9_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_decinfo[6]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo[6]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg9_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_decinfo[7]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo[7]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg9_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_decinfo[8]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo[8]));  // ../RTL/core/dispatch.v(90)
  AL_DFF_X \u_DISPATCH/reg9_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(bpu_decinfo[9]),
    .en(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(dis_decinfo[9]));  // ../RTL/core/dispatch.v(90)
  or \u_DISPATCH/u2  (\u_DISPATCH/n1 , n2, n3);  // ../RTL/core/dispatch.v(94)
  not \u_DISPATCH/u3  (\u_DISPATCH/n2 , bpu_inst_vld);  // ../RTL/core/dispatch.v(99)
  or \u_DISPATCH/u4  (\u_DISPATCH/n3 , n3, \u_DISPATCH/n2 );  // ../RTL/core/dispatch.v(99)
  AL_MUX \u_DISPATCH/u5  (
    .i0(bpu_rdwen),
    .i1(1'b0),
    .sel(\u_DISPATCH/n3 ),
    .o(\u_DISPATCH/n4 ));  // ../RTL/core/dispatch.v(99)
  AL_MUX \u_DISPATCH/u7  (
    .i0(bpu_taken),
    .i1(1'b0),
    .sel(\u_DISPATCH/n3 ),
    .o(\u_DISPATCH/n28 ));  // ../RTL/core/dispatch.v(117)
  EXU u_EXU (
    .i_clk(i_clk),
    .i_csr_rdata(dis_csr_rdata),
    .i_csr_zimm(dis_csr_zimm),
    .i_csridx(dis_csridx),
    .i_decinfo({dis_decinfo[9:1],1'b0}),
    .i_decinfo_grp(dis_decinfo_grp),
    .i_exu_op1(dis_exu_op1),
    .i_exu_op2(dis_exu_op2),
    .i_iaddr(dis_iaddr),
    .i_imm(dis_imm),
    .i_rdidx(dis_rdidx),
    .i_rdwen(dis_rdwen),
    .i_ribm_gnt(i_ribm_gnt1),
    .i_ribm_rdata(i_ribm_rdata1),
    .i_ribm_rsp(i_ribm_rsp1),
    .i_rs2rdata(dis_rs2rdata),
    .i_rstn(i_rstn),
    .i_vld(n5),
    .o_csr_wdata(wb_csr_wdata),
    .o_csr_wen(wb_csr_wen),
    .o_csridx(wb_csridx),
    .o_exu_jaddr(exu_jaddr),
    .o_exu_rdidx0(ctrl2exu_rdidx0),
    .o_exu_rdidx1(ctrl2exu_rdidx1),
    .o_exu_rdidx2(ctrl2exu_rdidx2),
    .o_exu_rdwen0(ctrl2exu_rdwen0),
    .o_exu_rdwen1(ctrl2exu_rdwen1),
    .o_exu_rdwen2(ctrl2exu_rdwen2),
    .o_exu_resource_match(ctrl2exu_resource_match),
    .o_exu_taken(exu_taken),
    .o_rdidx0(exu_rdidx0),
    .o_rdidx1(exu_rdidx1),
    .o_rdidx2(exu_rdidx2),
    .o_rdwdata0(exu_rdwdata0),
    .o_rdwdata1(exu_rdwdata1),
    .o_rdwdata2(exu_rdwdata2),
    .o_rdwen0(exu_rdwen0),
    .o_rdwen1(exu_rdwen1),
    .o_rdwen2(exu_rdwen2),
    .o_ribm_addr({o_ribm_addr1[31:24],open_n30,open_n31,open_n32,open_n33,open_n34,open_n35,open_n36,open_n37,o_ribm_addr1[15:2],open_n38,open_n39}),
    .o_ribm_mask(o_ribm_mask1),
    .o_ribm_req(o_ribm_req1),
    .o_ribm_wdata(o_ribm_wdata1),
    .o_ribm_wrcs(o_ribm_wrcs1));  // ../RTL/core/ritter_top.v(297)
  and \u_IFU/u1  (\u_IFU/n0 , ifu_fetch_vld, \u_IFU/data_vld );  // ../RTL/core/ifu.v(161)
  and \u_IFU/u3  (ifu_data_vld, \u_IFU/n0 , \u_IFU/fifo_cnt [0]);  // ../RTL/core/ifu.v(161)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b0  (
    .i0(bpu_jaddr_gen[0]),
    .i1(exu_jaddr_gen[0]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [0]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b1  (
    .i0(bpu_jaddr_gen[1]),
    .i1(exu_jaddr_gen[1]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [1]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b10  (
    .i0(bpu_jaddr_gen[10]),
    .i1(exu_jaddr_gen[10]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [10]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b11  (
    .i0(bpu_jaddr_gen[11]),
    .i1(exu_jaddr_gen[11]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [11]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b12  (
    .i0(bpu_jaddr_gen[12]),
    .i1(exu_jaddr_gen[12]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [12]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b13  (
    .i0(bpu_jaddr_gen[13]),
    .i1(exu_jaddr_gen[13]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [13]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b14  (
    .i0(bpu_jaddr_gen[14]),
    .i1(exu_jaddr_gen[14]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [14]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b15  (
    .i0(bpu_jaddr_gen[15]),
    .i1(exu_jaddr_gen[15]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [15]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b16  (
    .i0(bpu_jaddr_gen[16]),
    .i1(exu_jaddr_gen[16]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [16]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b17  (
    .i0(bpu_jaddr_gen[17]),
    .i1(exu_jaddr_gen[17]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [17]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b18  (
    .i0(bpu_jaddr_gen[18]),
    .i1(exu_jaddr_gen[18]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [18]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b19  (
    .i0(bpu_jaddr_gen[19]),
    .i1(exu_jaddr_gen[19]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [19]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b2  (
    .i0(bpu_jaddr_gen[2]),
    .i1(exu_jaddr_gen[2]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [2]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b20  (
    .i0(bpu_jaddr_gen[20]),
    .i1(exu_jaddr_gen[20]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [20]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b21  (
    .i0(bpu_jaddr_gen[21]),
    .i1(exu_jaddr_gen[21]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [21]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b22  (
    .i0(bpu_jaddr_gen[22]),
    .i1(exu_jaddr_gen[22]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [22]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b23  (
    .i0(bpu_jaddr_gen[23]),
    .i1(exu_jaddr_gen[23]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [23]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b24  (
    .i0(bpu_jaddr_gen[24]),
    .i1(exu_jaddr_gen[24]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [24]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b25  (
    .i0(bpu_jaddr_gen[25]),
    .i1(exu_jaddr_gen[25]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [25]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b26  (
    .i0(bpu_jaddr_gen[26]),
    .i1(exu_jaddr_gen[26]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [26]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b27  (
    .i0(bpu_jaddr_gen[27]),
    .i1(exu_jaddr_gen[27]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [27]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b28  (
    .i0(bpu_jaddr_gen[28]),
    .i1(exu_jaddr_gen[28]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [28]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b29  (
    .i0(bpu_jaddr_gen[29]),
    .i1(exu_jaddr_gen[29]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [29]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b3  (
    .i0(bpu_jaddr_gen[3]),
    .i1(exu_jaddr_gen[3]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [3]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b30  (
    .i0(bpu_jaddr_gen[30]),
    .i1(exu_jaddr_gen[30]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [30]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b31  (
    .i0(bpu_jaddr_gen[31]),
    .i1(exu_jaddr_gen[31]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [31]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b4  (
    .i0(bpu_jaddr_gen[4]),
    .i1(exu_jaddr_gen[4]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [4]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b5  (
    .i0(bpu_jaddr_gen[5]),
    .i1(exu_jaddr_gen[5]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [5]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b6  (
    .i0(bpu_jaddr_gen[6]),
    .i1(exu_jaddr_gen[6]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [6]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b7  (
    .i0(bpu_jaddr_gen[7]),
    .i1(exu_jaddr_gen[7]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [7]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b8  (
    .i0(bpu_jaddr_gen[8]),
    .i1(exu_jaddr_gen[8]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [8]));  // ../RTL/core/ifu_bju.v(35)
  binary_mux_s1_w1 \u_IFU/u_IFU_BJU/mux0_b9  (
    .i0(bpu_jaddr_gen[9]),
    .i1(exu_jaddr_gen[9]),
    .sel(exu_taken_gen),
    .o(\u_IFU/jump_addr [9]));  // ../RTL/core/ifu_bju.v(35)
  or \u_IFU/u_IFU_BJU/u0  (\u_IFU/jump_flag , exu_taken_gen, bpu_taken_gen);  // ../RTL/core/ifu_bju.v(33)
  AL_DFF_X \u_IFU/u_IFU_FETCH/handshake_rdy_last_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_FETCH/n7 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_FETCH/handshake_rdy_last ));  // ../RTL/core/ifu_fetch.v(75)
  not \u_IFU/u_IFU_FETCH/n2_inv  (\u_IFU/u_IFU_FETCH/n2_neg , \u_IFU/u_IFU_FETCH/n2 );
  and \u_IFU/u_IFU_FETCH/u10  (\u_IFU/data_vld , \u_IFU/u_IFU_FETCH/handshake_rdy_last , i_ribm_rsp0);  // ../RTL/core/ifu_fetch.v(72)
  not \u_IFU/u_IFU_FETCH/u14  (\u_IFU/u_IFU_FETCH/n1 , \u_IFU/pc_vld );  // ../RTL/core/ifu_fetch.v(80)
  and \u_IFU/u_IFU_FETCH/u15  (\u_IFU/u_IFU_FETCH/n2 , \u_IFU/jump_flag , \u_IFU/u_IFU_FETCH/n1 );  // ../RTL/core/ifu_fetch.v(80)
  not \u_IFU/u_IFU_FETCH/u16  (\u_IFU/u_IFU_FETCH/n3 , \u_IFU/u_IFU_FETCH/handshake_rdy_last );  // ../RTL/core/ifu_fetch.v(85)
  or \u_IFU/u_IFU_FETCH/u17  (\u_IFU/u_IFU_FETCH/n4 , i_ribm_rsp0, \u_IFU/u_IFU_FETCH/n3 );  // ../RTL/core/ifu_fetch.v(85)
  AL_MUX \u_IFU/u_IFU_FETCH/u18  (
    .i0(\u_IFU/u_IFU_FETCH/handshake_rdy_last ),
    .i1(\u_IFU/pc_vld ),
    .sel(\u_IFU/u_IFU_FETCH/n4 ),
    .o(\u_IFU/u_IFU_FETCH/n5 ));  // ../RTL/core/ifu_fetch.v(85)
  AL_MUX \u_IFU/u_IFU_FETCH/u20  (
    .i0(1'b0),
    .i1(\u_IFU/u_IFU_FETCH/n5 ),
    .sel(\u_IFU/u_IFU_FETCH/u20_sel_is_2_o ),
    .o(\u_IFU/u_IFU_FETCH/n7 ));
  and \u_IFU/u_IFU_FETCH/u20_sel_is_2  (\u_IFU/u_IFU_FETCH/u20_sel_is_2_o , \u_IFU/u_IFU_FETCH/n2_neg , ifu_fetch_vld);
  and \u_IFU/u_IFU_FETCH/u6  (o_ribm_req0, i_rstn, ifu_fetch_vld);  // ../RTL/core/ifu_fetch.v(63)
  and \u_IFU/u_IFU_FETCH/u8  (\u_IFU/pc_vld , o_ribm_req0, i_ribm_gnt0);  // ../RTL/core/ifu_fetch.v(67)
  add_pu1_pu1_o1 \u_IFU/u_IFU_FIFO/add0  (
    .i0(\u_IFU/u_IFU_FIFO/hptr ),
    .i1(1'b1),
    .o(\u_IFU/u_IFU_FIFO/n2 ));  // ../RTL/core/fifos.v(124)
  add_pu1_pu1_o1 \u_IFU/u_IFU_FIFO/add2  (
    .i0(\u_IFU/fifo_cnt ),
    .i1(1'b1),
    .o(\u_IFU/u_IFU_FIFO/n10 ));  // ../RTL/core/fifos.v(154)
  not \u_IFU/u_IFU_FIFO/hptr[0]_inv  (\u_IFU/u_IFU_FIFO/hptr[0]_neg , \u_IFU/u_IFU_FIFO/hptr [0]);
  AL_DFF_X \u_IFU/u_IFU_FIFO/hptr_reg[0]  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_FIFO/hptr_1 ),
    .en(\u_IFU/pc_vld ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_FIFO/hptr ));  // ../RTL/core/fifos.v(131)
  binary_mux_s1_w1 \u_IFU/u_IFU_FIFO/mux0_b0  (
    .i0(\u_IFU/u_IFU_FIFO/n2 ),
    .i1(1'b0),
    .sel(\u_IFU/u_IFU_FIFO/hptr[0]_neg ),
    .o(\u_IFU/u_IFU_FIFO/hptr_1 ));  // ../RTL/core/fifos.v(124)
  and \u_IFU/u_IFU_FIFO/mux4_b32_sel_is_1  (\u_IFU/u_IFU_FIFO/mux4_b32_sel_is_1_o , \u_IFU/pc_vld , \u_IFU/u_IFU_FIFO/hptr[0]_neg );
  and \u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2  (\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o , i_rstn, \u_IFU/u_IFU_FIFO/mux4_b32_sel_is_1_o );
  AL_DFF_X \u_IFU/u_IFU_FIFO/o_fifo_cnt_reg[0]  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_FIFO/n13 ),
    .en(~\u_IFU/u_IFU_FIFO/n9 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/fifo_cnt ));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/fetch_addr [0]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[0]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/fetch_addr [1]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[1]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[10]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[10]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[11]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[11]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[12]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[12]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[13]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[13]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[14]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[14]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[15]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[15]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[16]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[16]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[17]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[17]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[18]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[18]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[19]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[19]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[2]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[2]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[20]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[20]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[21]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[21]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[22]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[22]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[23]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[23]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[24]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[24]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[25]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[25]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[26]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[26]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[27]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[27]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[28]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[28]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[29]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[29]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[3]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[3]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[30]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[30]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[31]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[31]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[4]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[4]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[5]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[5]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[6]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[6]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[7]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[7]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[8]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[8]));  // ../RTL/core/fifos.v(131)
  AL_DFF_X \u_IFU/u_IFU_FIFO/reg0_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_ribm_addr0[9]),
    .en(\u_IFU/u_IFU_FIFO/mux5_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(ifu_iaddr[9]));  // ../RTL/core/fifos.v(131)
  add_pu1_mu1_o1 \u_IFU/u_IFU_FIFO/sub0  (
    .i0(\u_IFU/fifo_cnt ),
    .i1(1'b1),
    .o(\u_IFU/u_IFU_FIFO/n11 [0]));  // ../RTL/core/fifos.v(157)
  and \u_IFU/u_IFU_FIFO/u12  (\u_IFU/u_IFU_FIFO/n9 , \u_IFU/pc_vld , i_ribm_rsp0);  // ../RTL/core/fifos.v(150)
  AL_MUX \u_IFU/u_IFU_FIFO/u13  (
    .i0(\u_IFU/fifo_cnt ),
    .i1(\u_IFU/u_IFU_FIFO/n11 [0]),
    .sel(i_ribm_rsp0),
    .o(\u_IFU/u_IFU_FIFO/n12 ));  // ../RTL/core/fifos.v(156)
  AL_MUX \u_IFU/u_IFU_FIFO/u14  (
    .i0(\u_IFU/u_IFU_FIFO/n12 ),
    .i1(\u_IFU/u_IFU_FIFO/n10 ),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_FIFO/n13 ));  // ../RTL/core/fifos.v(153)
  add_pu30_pu30_o30 \u_IFU/u_IFU_PC/add0  (
    .i0(\u_IFU/jump_addr [31:2]),
    .i1(30'b000000000000000000000000000001),
    .o(\u_IFU/u_IFU_PC/n2 ));  // ../RTL/core/ifu_pc.v(32)
  add_pu30_pu30_o30 \u_IFU/u_IFU_PC/add1  (
    .i0(\u_IFU/u_IFU_PC/pc [31:2]),
    .i1(30'b000000000000000000000000000001),
    .o(\u_IFU/u_IFU_PC/n4 ));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b0  (
    .i0(\u_IFU/u_IFU_PC/pc [0]),
    .i1(\u_IFU/jump_addr [0]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/fetch_addr [0]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b1  (
    .i0(\u_IFU/u_IFU_PC/pc [1]),
    .i1(\u_IFU/jump_addr [1]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/fetch_addr [1]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b10  (
    .i0(\u_IFU/u_IFU_PC/n4 [8]),
    .i1(\u_IFU/u_IFU_PC/n3 [8]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [10]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b11  (
    .i0(\u_IFU/u_IFU_PC/n4 [9]),
    .i1(\u_IFU/u_IFU_PC/n3 [9]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [11]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b12  (
    .i0(\u_IFU/u_IFU_PC/n4 [10]),
    .i1(\u_IFU/u_IFU_PC/n3 [10]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [12]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b13  (
    .i0(\u_IFU/u_IFU_PC/n4 [11]),
    .i1(\u_IFU/u_IFU_PC/n3 [11]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [13]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b14  (
    .i0(\u_IFU/u_IFU_PC/n4 [12]),
    .i1(\u_IFU/u_IFU_PC/n3 [12]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [14]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b15  (
    .i0(\u_IFU/u_IFU_PC/n4 [13]),
    .i1(\u_IFU/u_IFU_PC/n3 [13]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [15]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b16  (
    .i0(\u_IFU/u_IFU_PC/n4 [14]),
    .i1(\u_IFU/u_IFU_PC/n3 [14]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [16]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b17  (
    .i0(\u_IFU/u_IFU_PC/n4 [15]),
    .i1(\u_IFU/u_IFU_PC/n3 [15]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [17]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b18  (
    .i0(\u_IFU/u_IFU_PC/n4 [16]),
    .i1(\u_IFU/u_IFU_PC/n3 [16]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [18]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b19  (
    .i0(\u_IFU/u_IFU_PC/n4 [17]),
    .i1(\u_IFU/u_IFU_PC/n3 [17]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [19]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b2  (
    .i0(\u_IFU/u_IFU_PC/n4 [0]),
    .i1(\u_IFU/u_IFU_PC/n3 [0]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [2]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b20  (
    .i0(\u_IFU/u_IFU_PC/n4 [18]),
    .i1(\u_IFU/u_IFU_PC/n3 [18]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [20]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b21  (
    .i0(\u_IFU/u_IFU_PC/n4 [19]),
    .i1(\u_IFU/u_IFU_PC/n3 [19]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [21]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b22  (
    .i0(\u_IFU/u_IFU_PC/n4 [20]),
    .i1(\u_IFU/u_IFU_PC/n3 [20]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [22]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b23  (
    .i0(\u_IFU/u_IFU_PC/n4 [21]),
    .i1(\u_IFU/u_IFU_PC/n3 [21]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [23]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b24  (
    .i0(\u_IFU/u_IFU_PC/n4 [22]),
    .i1(\u_IFU/u_IFU_PC/n3 [22]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [24]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b25  (
    .i0(\u_IFU/u_IFU_PC/n4 [23]),
    .i1(\u_IFU/u_IFU_PC/n3 [23]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [25]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b26  (
    .i0(\u_IFU/u_IFU_PC/n4 [24]),
    .i1(\u_IFU/u_IFU_PC/n3 [24]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [26]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b27  (
    .i0(\u_IFU/u_IFU_PC/n4 [25]),
    .i1(\u_IFU/u_IFU_PC/n3 [25]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [27]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b28  (
    .i0(\u_IFU/u_IFU_PC/n4 [26]),
    .i1(\u_IFU/u_IFU_PC/n3 [26]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [28]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b29  (
    .i0(\u_IFU/u_IFU_PC/n4 [27]),
    .i1(\u_IFU/u_IFU_PC/n3 [27]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [29]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b3  (
    .i0(\u_IFU/u_IFU_PC/n4 [1]),
    .i1(\u_IFU/u_IFU_PC/n3 [1]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [3]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b30  (
    .i0(\u_IFU/u_IFU_PC/n4 [28]),
    .i1(\u_IFU/u_IFU_PC/n3 [28]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [30]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b31  (
    .i0(\u_IFU/u_IFU_PC/n4 [29]),
    .i1(\u_IFU/u_IFU_PC/n3 [29]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [31]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b4  (
    .i0(\u_IFU/u_IFU_PC/n4 [2]),
    .i1(\u_IFU/u_IFU_PC/n3 [2]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [4]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b5  (
    .i0(\u_IFU/u_IFU_PC/n4 [3]),
    .i1(\u_IFU/u_IFU_PC/n3 [3]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [5]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b6  (
    .i0(\u_IFU/u_IFU_PC/n4 [4]),
    .i1(\u_IFU/u_IFU_PC/n3 [4]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [6]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b7  (
    .i0(\u_IFU/u_IFU_PC/n4 [5]),
    .i1(\u_IFU/u_IFU_PC/n3 [5]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [7]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b8  (
    .i0(\u_IFU/u_IFU_PC/n4 [6]),
    .i1(\u_IFU/u_IFU_PC/n3 [6]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [8]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux0_b9  (
    .i0(\u_IFU/u_IFU_PC/n4 [7]),
    .i1(\u_IFU/u_IFU_PC/n3 [7]),
    .sel(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n5 [9]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b0  (
    .i0(\u_IFU/u_IFU_PC/pc [0]),
    .i1(ifu_iaddr[0]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [0]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b1  (
    .i0(\u_IFU/u_IFU_PC/pc [1]),
    .i1(ifu_iaddr[1]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [1]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b10  (
    .i0(\u_IFU/u_IFU_PC/pc [10]),
    .i1(ifu_iaddr[10]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [10]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b11  (
    .i0(\u_IFU/u_IFU_PC/pc [11]),
    .i1(ifu_iaddr[11]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [11]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b12  (
    .i0(\u_IFU/u_IFU_PC/pc [12]),
    .i1(ifu_iaddr[12]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [12]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b13  (
    .i0(\u_IFU/u_IFU_PC/pc [13]),
    .i1(ifu_iaddr[13]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [13]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b14  (
    .i0(\u_IFU/u_IFU_PC/pc [14]),
    .i1(ifu_iaddr[14]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [14]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b15  (
    .i0(\u_IFU/u_IFU_PC/pc [15]),
    .i1(ifu_iaddr[15]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [15]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b16  (
    .i0(\u_IFU/u_IFU_PC/pc [16]),
    .i1(ifu_iaddr[16]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [16]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b17  (
    .i0(\u_IFU/u_IFU_PC/pc [17]),
    .i1(ifu_iaddr[17]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [17]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b18  (
    .i0(\u_IFU/u_IFU_PC/pc [18]),
    .i1(ifu_iaddr[18]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [18]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b19  (
    .i0(\u_IFU/u_IFU_PC/pc [19]),
    .i1(ifu_iaddr[19]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [19]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b2  (
    .i0(\u_IFU/u_IFU_PC/pc [2]),
    .i1(ifu_iaddr[2]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [2]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b20  (
    .i0(\u_IFU/u_IFU_PC/pc [20]),
    .i1(ifu_iaddr[20]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [20]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b21  (
    .i0(\u_IFU/u_IFU_PC/pc [21]),
    .i1(ifu_iaddr[21]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [21]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b22  (
    .i0(\u_IFU/u_IFU_PC/pc [22]),
    .i1(ifu_iaddr[22]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [22]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b23  (
    .i0(\u_IFU/u_IFU_PC/pc [23]),
    .i1(ifu_iaddr[23]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [23]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b24  (
    .i0(\u_IFU/u_IFU_PC/pc [24]),
    .i1(ifu_iaddr[24]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [24]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b25  (
    .i0(\u_IFU/u_IFU_PC/pc [25]),
    .i1(ifu_iaddr[25]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [25]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b26  (
    .i0(\u_IFU/u_IFU_PC/pc [26]),
    .i1(ifu_iaddr[26]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [26]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b27  (
    .i0(\u_IFU/u_IFU_PC/pc [27]),
    .i1(ifu_iaddr[27]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [27]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b28  (
    .i0(\u_IFU/u_IFU_PC/pc [28]),
    .i1(ifu_iaddr[28]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [28]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b29  (
    .i0(\u_IFU/u_IFU_PC/pc [29]),
    .i1(ifu_iaddr[29]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [29]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b3  (
    .i0(\u_IFU/u_IFU_PC/pc [3]),
    .i1(ifu_iaddr[3]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [3]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b30  (
    .i0(\u_IFU/u_IFU_PC/pc [30]),
    .i1(ifu_iaddr[30]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [30]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b31  (
    .i0(\u_IFU/u_IFU_PC/pc [31]),
    .i1(ifu_iaddr[31]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [31]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b4  (
    .i0(\u_IFU/u_IFU_PC/pc [4]),
    .i1(ifu_iaddr[4]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [4]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b5  (
    .i0(\u_IFU/u_IFU_PC/pc [5]),
    .i1(ifu_iaddr[5]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [5]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b6  (
    .i0(\u_IFU/u_IFU_PC/pc [6]),
    .i1(ifu_iaddr[6]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [6]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b7  (
    .i0(\u_IFU/u_IFU_PC/pc [7]),
    .i1(ifu_iaddr[7]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [7]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b8  (
    .i0(\u_IFU/u_IFU_PC/pc [8]),
    .i1(ifu_iaddr[8]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [8]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux1_b9  (
    .i0(\u_IFU/u_IFU_PC/pc [9]),
    .i1(ifu_iaddr[9]),
    .sel(\u_IFU/u_IFU_PC/n8 ),
    .o(\u_IFU/u_IFU_PC/n9 [9]));  // ../RTL/core/ifu_pc.v(34)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b0  (
    .i0(\u_IFU/u_IFU_PC/n9 [0]),
    .i1(\u_IFU/fetch_addr [0]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [0]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b1  (
    .i0(\u_IFU/u_IFU_PC/n9 [1]),
    .i1(\u_IFU/fetch_addr [1]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [1]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b10  (
    .i0(\u_IFU/u_IFU_PC/n9 [10]),
    .i1(\u_IFU/u_IFU_PC/n5 [10]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [10]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b11  (
    .i0(\u_IFU/u_IFU_PC/n9 [11]),
    .i1(\u_IFU/u_IFU_PC/n5 [11]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [11]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b12  (
    .i0(\u_IFU/u_IFU_PC/n9 [12]),
    .i1(\u_IFU/u_IFU_PC/n5 [12]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [12]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b13  (
    .i0(\u_IFU/u_IFU_PC/n9 [13]),
    .i1(\u_IFU/u_IFU_PC/n5 [13]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [13]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b14  (
    .i0(\u_IFU/u_IFU_PC/n9 [14]),
    .i1(\u_IFU/u_IFU_PC/n5 [14]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [14]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b15  (
    .i0(\u_IFU/u_IFU_PC/n9 [15]),
    .i1(\u_IFU/u_IFU_PC/n5 [15]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [15]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b16  (
    .i0(\u_IFU/u_IFU_PC/n9 [16]),
    .i1(\u_IFU/u_IFU_PC/n5 [16]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [16]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b17  (
    .i0(\u_IFU/u_IFU_PC/n9 [17]),
    .i1(\u_IFU/u_IFU_PC/n5 [17]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [17]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b18  (
    .i0(\u_IFU/u_IFU_PC/n9 [18]),
    .i1(\u_IFU/u_IFU_PC/n5 [18]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [18]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b19  (
    .i0(\u_IFU/u_IFU_PC/n9 [19]),
    .i1(\u_IFU/u_IFU_PC/n5 [19]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [19]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b2  (
    .i0(\u_IFU/u_IFU_PC/n9 [2]),
    .i1(\u_IFU/u_IFU_PC/n5 [2]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [2]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b20  (
    .i0(\u_IFU/u_IFU_PC/n9 [20]),
    .i1(\u_IFU/u_IFU_PC/n5 [20]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [20]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b21  (
    .i0(\u_IFU/u_IFU_PC/n9 [21]),
    .i1(\u_IFU/u_IFU_PC/n5 [21]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [21]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b22  (
    .i0(\u_IFU/u_IFU_PC/n9 [22]),
    .i1(\u_IFU/u_IFU_PC/n5 [22]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [22]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b23  (
    .i0(\u_IFU/u_IFU_PC/n9 [23]),
    .i1(\u_IFU/u_IFU_PC/n5 [23]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [23]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b24  (
    .i0(\u_IFU/u_IFU_PC/n9 [24]),
    .i1(\u_IFU/u_IFU_PC/n5 [24]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [24]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b25  (
    .i0(\u_IFU/u_IFU_PC/n9 [25]),
    .i1(\u_IFU/u_IFU_PC/n5 [25]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [25]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b26  (
    .i0(\u_IFU/u_IFU_PC/n9 [26]),
    .i1(\u_IFU/u_IFU_PC/n5 [26]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [26]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b27  (
    .i0(\u_IFU/u_IFU_PC/n9 [27]),
    .i1(\u_IFU/u_IFU_PC/n5 [27]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [27]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b28  (
    .i0(\u_IFU/u_IFU_PC/n9 [28]),
    .i1(\u_IFU/u_IFU_PC/n5 [28]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [28]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b29  (
    .i0(\u_IFU/u_IFU_PC/n9 [29]),
    .i1(\u_IFU/u_IFU_PC/n5 [29]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [29]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b3  (
    .i0(\u_IFU/u_IFU_PC/n9 [3]),
    .i1(\u_IFU/u_IFU_PC/n5 [3]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [3]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b30  (
    .i0(\u_IFU/u_IFU_PC/n9 [30]),
    .i1(\u_IFU/u_IFU_PC/n5 [30]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [30]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b31  (
    .i0(\u_IFU/u_IFU_PC/n9 [31]),
    .i1(\u_IFU/u_IFU_PC/n5 [31]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [31]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b4  (
    .i0(\u_IFU/u_IFU_PC/n9 [4]),
    .i1(\u_IFU/u_IFU_PC/n5 [4]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [4]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b5  (
    .i0(\u_IFU/u_IFU_PC/n9 [5]),
    .i1(\u_IFU/u_IFU_PC/n5 [5]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [5]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b6  (
    .i0(\u_IFU/u_IFU_PC/n9 [6]),
    .i1(\u_IFU/u_IFU_PC/n5 [6]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [6]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b7  (
    .i0(\u_IFU/u_IFU_PC/n9 [7]),
    .i1(\u_IFU/u_IFU_PC/n5 [7]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [7]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b8  (
    .i0(\u_IFU/u_IFU_PC/n9 [8]),
    .i1(\u_IFU/u_IFU_PC/n5 [8]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [8]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux2_b9  (
    .i0(\u_IFU/u_IFU_PC/n9 [9]),
    .i1(\u_IFU/u_IFU_PC/n5 [9]),
    .sel(\u_IFU/u_IFU_PC/n1 ),
    .o(\u_IFU/u_IFU_PC/n10 [9]));  // ../RTL/core/ifu_pc.v(31)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b0  (
    .i0(\u_IFU/jump_addr [2]),
    .i1(\u_IFU/u_IFU_PC/n2 [0]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [0]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b1  (
    .i0(\u_IFU/jump_addr [3]),
    .i1(\u_IFU/u_IFU_PC/n2 [1]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [1]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b10  (
    .i0(\u_IFU/jump_addr [12]),
    .i1(\u_IFU/u_IFU_PC/n2 [10]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [10]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b11  (
    .i0(\u_IFU/jump_addr [13]),
    .i1(\u_IFU/u_IFU_PC/n2 [11]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [11]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b12  (
    .i0(\u_IFU/jump_addr [14]),
    .i1(\u_IFU/u_IFU_PC/n2 [12]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [12]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b13  (
    .i0(\u_IFU/jump_addr [15]),
    .i1(\u_IFU/u_IFU_PC/n2 [13]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [13]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b14  (
    .i0(\u_IFU/jump_addr [16]),
    .i1(\u_IFU/u_IFU_PC/n2 [14]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [14]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b15  (
    .i0(\u_IFU/jump_addr [17]),
    .i1(\u_IFU/u_IFU_PC/n2 [15]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [15]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b16  (
    .i0(\u_IFU/jump_addr [18]),
    .i1(\u_IFU/u_IFU_PC/n2 [16]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [16]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b17  (
    .i0(\u_IFU/jump_addr [19]),
    .i1(\u_IFU/u_IFU_PC/n2 [17]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [17]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b18  (
    .i0(\u_IFU/jump_addr [20]),
    .i1(\u_IFU/u_IFU_PC/n2 [18]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [18]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b19  (
    .i0(\u_IFU/jump_addr [21]),
    .i1(\u_IFU/u_IFU_PC/n2 [19]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [19]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b2  (
    .i0(\u_IFU/jump_addr [4]),
    .i1(\u_IFU/u_IFU_PC/n2 [2]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [2]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b20  (
    .i0(\u_IFU/jump_addr [22]),
    .i1(\u_IFU/u_IFU_PC/n2 [20]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [20]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b21  (
    .i0(\u_IFU/jump_addr [23]),
    .i1(\u_IFU/u_IFU_PC/n2 [21]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [21]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b22  (
    .i0(\u_IFU/jump_addr [24]),
    .i1(\u_IFU/u_IFU_PC/n2 [22]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [22]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b23  (
    .i0(\u_IFU/jump_addr [25]),
    .i1(\u_IFU/u_IFU_PC/n2 [23]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [23]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b24  (
    .i0(\u_IFU/jump_addr [26]),
    .i1(\u_IFU/u_IFU_PC/n2 [24]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [24]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b25  (
    .i0(\u_IFU/jump_addr [27]),
    .i1(\u_IFU/u_IFU_PC/n2 [25]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [25]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b26  (
    .i0(\u_IFU/jump_addr [28]),
    .i1(\u_IFU/u_IFU_PC/n2 [26]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [26]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b27  (
    .i0(\u_IFU/jump_addr [29]),
    .i1(\u_IFU/u_IFU_PC/n2 [27]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [27]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b28  (
    .i0(\u_IFU/jump_addr [30]),
    .i1(\u_IFU/u_IFU_PC/n2 [28]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [28]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b29  (
    .i0(\u_IFU/jump_addr [31]),
    .i1(\u_IFU/u_IFU_PC/n2 [29]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [29]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b3  (
    .i0(\u_IFU/jump_addr [5]),
    .i1(\u_IFU/u_IFU_PC/n2 [3]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [3]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b4  (
    .i0(\u_IFU/jump_addr [6]),
    .i1(\u_IFU/u_IFU_PC/n2 [4]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [4]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b5  (
    .i0(\u_IFU/jump_addr [7]),
    .i1(\u_IFU/u_IFU_PC/n2 [5]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [5]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b6  (
    .i0(\u_IFU/jump_addr [8]),
    .i1(\u_IFU/u_IFU_PC/n2 [6]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [6]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b7  (
    .i0(\u_IFU/jump_addr [9]),
    .i1(\u_IFU/u_IFU_PC/n2 [7]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [7]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b8  (
    .i0(\u_IFU/jump_addr [10]),
    .i1(\u_IFU/u_IFU_PC/n2 [8]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [8]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux3_b9  (
    .i0(\u_IFU/jump_addr [11]),
    .i1(\u_IFU/u_IFU_PC/n2 [9]),
    .sel(\u_IFU/pc_vld ),
    .o(\u_IFU/u_IFU_PC/n3 [9]));  // ../RTL/core/ifu_pc.v(32)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b10  (
    .i0(\u_IFU/u_IFU_PC/pc [10]),
    .i1(\u_IFU/jump_addr [10]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[10]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b11  (
    .i0(\u_IFU/u_IFU_PC/pc [11]),
    .i1(\u_IFU/jump_addr [11]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[11]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b12  (
    .i0(\u_IFU/u_IFU_PC/pc [12]),
    .i1(\u_IFU/jump_addr [12]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[12]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b13  (
    .i0(\u_IFU/u_IFU_PC/pc [13]),
    .i1(\u_IFU/jump_addr [13]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[13]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b14  (
    .i0(\u_IFU/u_IFU_PC/pc [14]),
    .i1(\u_IFU/jump_addr [14]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[14]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b15  (
    .i0(\u_IFU/u_IFU_PC/pc [15]),
    .i1(\u_IFU/jump_addr [15]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[15]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b16  (
    .i0(\u_IFU/u_IFU_PC/pc [16]),
    .i1(\u_IFU/jump_addr [16]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[16]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b17  (
    .i0(\u_IFU/u_IFU_PC/pc [17]),
    .i1(\u_IFU/jump_addr [17]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[17]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b18  (
    .i0(\u_IFU/u_IFU_PC/pc [18]),
    .i1(\u_IFU/jump_addr [18]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[18]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b19  (
    .i0(\u_IFU/u_IFU_PC/pc [19]),
    .i1(\u_IFU/jump_addr [19]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[19]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b2  (
    .i0(\u_IFU/u_IFU_PC/pc [2]),
    .i1(\u_IFU/jump_addr [2]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[2]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b20  (
    .i0(\u_IFU/u_IFU_PC/pc [20]),
    .i1(\u_IFU/jump_addr [20]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[20]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b21  (
    .i0(\u_IFU/u_IFU_PC/pc [21]),
    .i1(\u_IFU/jump_addr [21]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[21]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b22  (
    .i0(\u_IFU/u_IFU_PC/pc [22]),
    .i1(\u_IFU/jump_addr [22]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[22]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b23  (
    .i0(\u_IFU/u_IFU_PC/pc [23]),
    .i1(\u_IFU/jump_addr [23]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[23]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b24  (
    .i0(\u_IFU/u_IFU_PC/pc [24]),
    .i1(\u_IFU/jump_addr [24]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[24]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b25  (
    .i0(\u_IFU/u_IFU_PC/pc [25]),
    .i1(\u_IFU/jump_addr [25]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[25]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b26  (
    .i0(\u_IFU/u_IFU_PC/pc [26]),
    .i1(\u_IFU/jump_addr [26]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[26]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b27  (
    .i0(\u_IFU/u_IFU_PC/pc [27]),
    .i1(\u_IFU/jump_addr [27]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[27]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b28  (
    .i0(\u_IFU/u_IFU_PC/pc [28]),
    .i1(\u_IFU/jump_addr [28]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[28]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b29  (
    .i0(\u_IFU/u_IFU_PC/pc [29]),
    .i1(\u_IFU/jump_addr [29]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[29]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b3  (
    .i0(\u_IFU/u_IFU_PC/pc [3]),
    .i1(\u_IFU/jump_addr [3]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[3]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b30  (
    .i0(\u_IFU/u_IFU_PC/pc [30]),
    .i1(\u_IFU/jump_addr [30]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[30]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b31  (
    .i0(\u_IFU/u_IFU_PC/pc [31]),
    .i1(\u_IFU/jump_addr [31]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[31]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b4  (
    .i0(\u_IFU/u_IFU_PC/pc [4]),
    .i1(\u_IFU/jump_addr [4]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[4]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b5  (
    .i0(\u_IFU/u_IFU_PC/pc [5]),
    .i1(\u_IFU/jump_addr [5]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[5]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b6  (
    .i0(\u_IFU/u_IFU_PC/pc [6]),
    .i1(\u_IFU/jump_addr [6]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[6]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b7  (
    .i0(\u_IFU/u_IFU_PC/pc [7]),
    .i1(\u_IFU/jump_addr [7]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[7]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b8  (
    .i0(\u_IFU/u_IFU_PC/pc [8]),
    .i1(\u_IFU/jump_addr [8]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[8]));  // ../RTL/core/ifu_pc.v(41)
  binary_mux_s1_w1 \u_IFU/u_IFU_PC/mux4_b9  (
    .i0(\u_IFU/u_IFU_PC/pc [9]),
    .i1(\u_IFU/jump_addr [9]),
    .sel(\u_IFU/jump_flag ),
    .o(o_ribm_addr0[9]));  // ../RTL/core/ifu_pc.v(41)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [0]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b1  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [1]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b10  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [10]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b11  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [11]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b12  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [12]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b13  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [13]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b14  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [14]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b15  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [15]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b16  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [16]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b17  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [17]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b18  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [18]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b19  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [19]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b2  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [2]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b20  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [20]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b21  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [21]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b22  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [22]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b23  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [23]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b24  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [24]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b25  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [25]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b26  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [26]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b27  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [27]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b28  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [28]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b29  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [29]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b3  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [3]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b30  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [30]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b31  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [31]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b4  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [4]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b5  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [5]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b6  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [6]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b7  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [7]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b8  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [8]));  // ../RTL/core/ifu_pc.v(26)
  AL_DFF_X \u_IFU/u_IFU_PC/reg0_b9  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU/u_IFU_PC/pc [9]));  // ../RTL/core/ifu_pc.v(26)
  or \u_IFU/u_IFU_PC/u3  (\u_IFU/u_IFU_PC/n1 , \u_IFU/pc_vld , \u_IFU/jump_flag );  // ../RTL/core/ifu_pc.v(31)
  not \u_IFU/u_IFU_PC/u5  (\u_IFU/u_IFU_PC/n7 , ifu_fetch_vld);  // ../RTL/core/ifu_pc.v(34)
  and \u_IFU/u_IFU_PC/u6  (\u_IFU/u_IFU_PC/n8 , \u_IFU/fifo_cnt [0], \u_IFU/u_IFU_PC/n7 );  // ../RTL/core/ifu_pc.v(34)
  and \u_IFU2BPU/u13  (\u_IFU2BPU/n2 , ctrl2bpu_wait, \u_IFU2BPU/fifo_full );  // ../RTL/core/ifu2bpu.v(60)
  not \u_IFU2BPU/u14  (bpu2ifu_vld, \u_IFU2BPU/n2 );  // ../RTL/core/ifu2bpu.v(60)
  not \u_IFU2BPU/u4  (ifu2bpu_data_vld, \u_IFU2BPU/fifo_empty );  // ../RTL/core/ifu2bpu.v(52)
  and \u_IFU2BPU/u5  (\u_IFU2BPU/n0 , n1, ifu2bpu_data_vld);  // ../RTL/core/ifu2bpu.v(52)
  add_pu4_pu4_o4 \u_IFU2BPU/u_SYNC_FIFO/add0  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/hptr ),
    .i1(4'b0001),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n2 ));  // ../RTL/core/fifos.v(40)
  add_pu4_pu4_o4 \u_IFU2BPU/u_SYNC_FIFO/add1  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/eptr ),
    .i1(4'b0001),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n5 ));  // ../RTL/core/fifos.v(42)
  add_pu4_pu4_o4 \u_IFU2BPU/u_SYNC_FIFO/add2  (
    .i0(\u_IFU2BPU/fifo_cnt [3:0]),
    .i1(4'b0001),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n10 ));  // ../RTL/core/fifos.v(64)
  EG_LOGIC_DRAM #(
    .ADDR_WIDTH_R(3),
    .ADDR_WIDTH_W(3),
    .DATA_DEPTH_R(8),
    .DATA_DEPTH_W(8),
    .DATA_WIDTH_R(64),
    .DATA_WIDTH_W(64))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units  (
    .di({i_ribm_rdata0,ifu_iaddr}),
    .raddr(\u_IFU2BPU/u_SYNC_FIFO/eptr [2:0]),
    .waddr(\u_IFU2BPU/u_SYNC_FIFO/hptr [2:0]),
    .wclk(i_clk),
    .we(\u_IFU2BPU/u_SYNC_FIFO/n19 ),
    .do({ifu2bpu_data,ifu2bpu_iaddr}));
  eq_w4 \u_IFU2BPU/u_SYNC_FIFO/eq0  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/hptr ),
    .i1(4'b0111),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n0 ));  // ../RTL/core/fifos.v(40)
  eq_w4 \u_IFU2BPU/u_SYNC_FIFO/eq1  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/eptr ),
    .i1(4'b0111),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n3 ));  // ../RTL/core/fifos.v(42)
  eq_w4 \u_IFU2BPU/u_SYNC_FIFO/eq2  (
    .i0(\u_IFU2BPU/fifo_cnt [3:0]),
    .i1(4'b1000),
    .o(\u_IFU2BPU/fifo_full ));  // ../RTL/core/fifos.v(44)
  eq_w4 \u_IFU2BPU/u_SYNC_FIFO/eq3  (
    .i0(\u_IFU2BPU/fifo_cnt [3:0]),
    .i1(4'b0000),
    .o(\u_IFU2BPU/fifo_empty ));  // ../RTL/core/fifos.v(45)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux0_b0  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n2 [0]),
    .i1(1'b0),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n0 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/hptr_1 [0]));  // ../RTL/core/fifos.v(40)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux0_b1  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n2 [1]),
    .i1(1'b0),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n0 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/hptr_1 [1]));  // ../RTL/core/fifos.v(40)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux0_b2  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n2 [2]),
    .i1(1'b0),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n0 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/hptr_1 [2]));  // ../RTL/core/fifos.v(40)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux0_b3  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n2 [3]),
    .i1(1'b0),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n0 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/hptr_1 [3]));  // ../RTL/core/fifos.v(40)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux1_b0  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n5 [0]),
    .i1(1'b0),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n3 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/eptr_1 [0]));  // ../RTL/core/fifos.v(42)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux1_b1  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n5 [1]),
    .i1(1'b0),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n3 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/eptr_1 [1]));  // ../RTL/core/fifos.v(42)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux1_b2  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n5 [2]),
    .i1(1'b0),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n3 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/eptr_1 [2]));  // ../RTL/core/fifos.v(42)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux1_b3  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n5 [3]),
    .i1(1'b0),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n3 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/eptr_1 [3]));  // ../RTL/core/fifos.v(42)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux2_b0  (
    .i0(\u_IFU2BPU/fifo_cnt [0]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/n13 [0]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n12 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n14 [0]));  // ../RTL/core/fifos.v(66)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux2_b1  (
    .i0(\u_IFU2BPU/fifo_cnt [1]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/n13 [1]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n12 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n14 [1]));  // ../RTL/core/fifos.v(66)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux2_b2  (
    .i0(\u_IFU2BPU/fifo_cnt [2]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/n13 [2]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n12 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n14 [2]));  // ../RTL/core/fifos.v(66)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux2_b3  (
    .i0(\u_IFU2BPU/fifo_cnt [3]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/n13 [3]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n12 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n14 [3]));  // ../RTL/core/fifos.v(66)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux3_b0  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n14 [0]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/n10 [0]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n9 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n15 [0]));  // ../RTL/core/fifos.v(63)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux3_b1  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n14 [1]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/n10 [1]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n9 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n15 [1]));  // ../RTL/core/fifos.v(63)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux3_b2  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n14 [2]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/n10 [2]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n9 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n15 [2]));  // ../RTL/core/fifos.v(63)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux3_b3  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n14 [3]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/n10 [3]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n9 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n15 [3]));  // ../RTL/core/fifos.v(63)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux4_b0  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n15 [0]),
    .i1(\u_IFU2BPU/fifo_cnt [0]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n7 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n16 [0]));  // ../RTL/core/fifos.v(60)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux4_b1  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n15 [1]),
    .i1(\u_IFU2BPU/fifo_cnt [1]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n7 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n16 [1]));  // ../RTL/core/fifos.v(60)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux4_b2  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n15 [2]),
    .i1(\u_IFU2BPU/fifo_cnt [2]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n7 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n16 [2]));  // ../RTL/core/fifos.v(60)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux4_b3  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n15 [3]),
    .i1(\u_IFU2BPU/fifo_cnt [3]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n7 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n16 [3]));  // ../RTL/core/fifos.v(60)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux5_b0  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/hptr [0]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/hptr_1 [0]),
    .sel(ifu_data_vld),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n20 [0]));  // ../RTL/core/fifos.v(71)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux5_b1  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/hptr [1]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/hptr_1 [1]),
    .sel(ifu_data_vld),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n20 [1]));  // ../RTL/core/fifos.v(71)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux5_b2  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/hptr [2]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/hptr_1 [2]),
    .sel(ifu_data_vld),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n20 [2]));  // ../RTL/core/fifos.v(71)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux5_b3  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/hptr [3]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/hptr_1 [3]),
    .sel(ifu_data_vld),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n20 [3]));  // ../RTL/core/fifos.v(71)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux6_b0  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/eptr [0]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/eptr_1 [0]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n12 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n21 [0]));  // ../RTL/core/fifos.v(75)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux6_b1  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/eptr [1]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/eptr_1 [1]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n12 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n21 [1]));  // ../RTL/core/fifos.v(75)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux6_b2  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/eptr [2]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/eptr_1 [2]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n12 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n21 [2]));  // ../RTL/core/fifos.v(75)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux6_b3  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/eptr [3]),
    .i1(\u_IFU2BPU/u_SYNC_FIFO/eptr_1 [3]),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/n12 ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n21 [3]));  // ../RTL/core/fifos.v(75)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux7_b0  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n20 [0]),
    .i1(1'b0),
    .sel(n0),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n22 [0]));  // ../RTL/core/fifos.v(53)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux7_b1  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n20 [1]),
    .i1(1'b0),
    .sel(n0),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n22 [1]));  // ../RTL/core/fifos.v(53)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux7_b2  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n20 [2]),
    .i1(1'b0),
    .sel(n0),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n22 [2]));  // ../RTL/core/fifos.v(53)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux7_b3  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n20 [3]),
    .i1(1'b0),
    .sel(n0),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n22 [3]));  // ../RTL/core/fifos.v(53)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux8_b0  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n21 [0]),
    .i1(1'b0),
    .sel(n0),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n23 [0]));  // ../RTL/core/fifos.v(53)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux8_b1  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n21 [1]),
    .i1(1'b0),
    .sel(n0),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n23 [1]));  // ../RTL/core/fifos.v(53)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux8_b2  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n21 [2]),
    .i1(1'b0),
    .sel(n0),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n23 [2]));  // ../RTL/core/fifos.v(53)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux8_b3  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n21 [3]),
    .i1(1'b0),
    .sel(n0),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n23 [3]));  // ../RTL/core/fifos.v(53)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux9_b0  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n16 [0]),
    .i1(1'b0),
    .sel(n0),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n24 [0]));  // ../RTL/core/fifos.v(53)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux9_b1  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n16 [1]),
    .i1(1'b0),
    .sel(n0),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n24 [1]));  // ../RTL/core/fifos.v(53)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux9_b2  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n16 [2]),
    .i1(1'b0),
    .sel(n0),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n24 [2]));  // ../RTL/core/fifos.v(53)
  binary_mux_s1_w1 \u_IFU2BPU/u_SYNC_FIFO/mux9_b3  (
    .i0(\u_IFU2BPU/u_SYNC_FIFO/n16 [3]),
    .i1(1'b0),
    .sel(n0),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n24 [3]));  // ../RTL/core/fifos.v(53)
  AL_DFF_X \u_IFU2BPU/u_SYNC_FIFO/reg0_b0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n23 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU2BPU/u_SYNC_FIFO/eptr [0]));  // ../RTL/core/fifos.v(48)
  AL_DFF_X \u_IFU2BPU/u_SYNC_FIFO/reg0_b1  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n23 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU2BPU/u_SYNC_FIFO/eptr [1]));  // ../RTL/core/fifos.v(48)
  AL_DFF_X \u_IFU2BPU/u_SYNC_FIFO/reg0_b2  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n23 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU2BPU/u_SYNC_FIFO/eptr [2]));  // ../RTL/core/fifos.v(48)
  AL_DFF_X \u_IFU2BPU/u_SYNC_FIFO/reg0_b3  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n23 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU2BPU/u_SYNC_FIFO/eptr [3]));  // ../RTL/core/fifos.v(48)
  AL_DFF_X \u_IFU2BPU/u_SYNC_FIFO/reg1_b0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n24 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU2BPU/fifo_cnt [0]));  // ../RTL/core/fifos.v(48)
  AL_DFF_X \u_IFU2BPU/u_SYNC_FIFO/reg1_b1  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n24 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU2BPU/fifo_cnt [1]));  // ../RTL/core/fifos.v(48)
  AL_DFF_X \u_IFU2BPU/u_SYNC_FIFO/reg1_b2  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n24 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU2BPU/fifo_cnt [2]));  // ../RTL/core/fifos.v(48)
  AL_DFF_X \u_IFU2BPU/u_SYNC_FIFO/reg1_b3  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n24 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU2BPU/fifo_cnt [3]));  // ../RTL/core/fifos.v(48)
  AL_DFF_X \u_IFU2BPU/u_SYNC_FIFO/reg2_b0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n22 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU2BPU/u_SYNC_FIFO/hptr [0]));  // ../RTL/core/fifos.v(48)
  AL_DFF_X \u_IFU2BPU/u_SYNC_FIFO/reg2_b1  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n22 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU2BPU/u_SYNC_FIFO/hptr [1]));  // ../RTL/core/fifos.v(48)
  AL_DFF_X \u_IFU2BPU/u_SYNC_FIFO/reg2_b2  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n22 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU2BPU/u_SYNC_FIFO/hptr [2]));  // ../RTL/core/fifos.v(48)
  AL_DFF_X \u_IFU2BPU/u_SYNC_FIFO/reg2_b3  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n22 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_IFU2BPU/u_SYNC_FIFO/hptr [3]));  // ../RTL/core/fifos.v(48)
  add_pu4_mu4_o4 \u_IFU2BPU/u_SYNC_FIFO/sub0  (
    .i0(\u_IFU2BPU/fifo_cnt [3:0]),
    .i1(4'b0001),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n13 [3:0]));  // ../RTL/core/fifos.v(67)
  AL_MUX \u_IFU2BPU/u_SYNC_FIFO/u11  (
    .i0(1'b0),
    .i1(ifu_data_vld),
    .sel(\u_IFU2BPU/u_SYNC_FIFO/u11_sel_is_0_o ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n18 ));
  and \u_IFU2BPU/u_SYNC_FIFO/u11_sel_is_0  (\u_IFU2BPU/u_SYNC_FIFO/u11_sel_is_0_o , i_rstn, n0_neg);
  not \u_IFU2BPU/u_SYNC_FIFO/u2  (\u_IFU2BPU/u_SYNC_FIFO/n17 , \u_IFU2BPU/u_SYNC_FIFO/hptr [3]);  // ../RTL/core/fifos.v(72)
  and \u_IFU2BPU/u_SYNC_FIFO/u4  (\u_IFU2BPU/u_SYNC_FIFO/n7 , ifu_data_vld, \u_IFU2BPU/n0 );  // ../RTL/core/fifos.v(60)
  not \u_IFU2BPU/u_SYNC_FIFO/u5  (\u_IFU2BPU/u_SYNC_FIFO/n8 , \u_IFU2BPU/fifo_full );  // ../RTL/core/fifos.v(63)
  and \u_IFU2BPU/u_SYNC_FIFO/u6  (\u_IFU2BPU/u_SYNC_FIFO/n9 , ifu_data_vld, \u_IFU2BPU/u_SYNC_FIFO/n8 );  // ../RTL/core/fifos.v(63)
  and \u_IFU2BPU/u_SYNC_FIFO/u8  (\u_IFU2BPU/u_SYNC_FIFO/n12 , \u_IFU2BPU/n0 , ifu2bpu_data_vld);  // ../RTL/core/fifos.v(66)
  and \u_IFU2BPU/u_SYNC_FIFO/u9  (\u_IFU2BPU/u_SYNC_FIFO/n19 , \u_IFU2BPU/u_SYNC_FIFO/n17 , \u_IFU2BPU/u_SYNC_FIFO/n18 );  // ../RTL/core/fifos.v(72)
  eq_w5 \u_PIPE_CTRL/eq0  (
    .i0(ctrl2bpu_rs1idx),
    .i1(ctrl2exu_rdidx0),
    .o(\u_PIPE_CTRL/n0 ));  // ../RTL/core/pipe_ctrl.v(42)
  eq_w5 \u_PIPE_CTRL/eq1  (
    .i0(ctrl2bpu_rs1idx),
    .i1(ctrl2exu_rdidx1),
    .o(\u_PIPE_CTRL/n2 ));  // ../RTL/core/pipe_ctrl.v(43)
  eq_w5 \u_PIPE_CTRL/eq2  (
    .i0(ctrl2bpu_rs1idx),
    .i1(ctrl2exu_rdidx2),
    .o(\u_PIPE_CTRL/n5 ));  // ../RTL/core/pipe_ctrl.v(44)
  eq_w5 \u_PIPE_CTRL/eq3  (
    .i0(ctrl2bpu_rs2idx),
    .i1(ctrl2exu_rdidx0),
    .o(\u_PIPE_CTRL/n8 ));  // ../RTL/core/pipe_ctrl.v(46)
  eq_w5 \u_PIPE_CTRL/eq4  (
    .i0(ctrl2bpu_rs2idx),
    .i1(ctrl2exu_rdidx1),
    .o(\u_PIPE_CTRL/n10 ));  // ../RTL/core/pipe_ctrl.v(47)
  eq_w5 \u_PIPE_CTRL/eq5  (
    .i0(ctrl2bpu_rs2idx),
    .i1(ctrl2exu_rdidx2),
    .o(\u_PIPE_CTRL/n13 ));  // ../RTL/core/pipe_ctrl.v(48)
  binary_mux_s1_w1 \u_PIPE_CTRL/mux0_b0  (
    .i0(1'b0),
    .i1(\u_PIPE_CTRL/n7 [0]),
    .sel(ctrl2bpu_rs1ren),
    .o(\u_PIPE_CTRL/rs1_match ));  // ../RTL/core/pipe_ctrl.v(41)
  binary_mux_s1_w1 \u_PIPE_CTRL/mux1_b0  (
    .i0(1'b0),
    .i1(\u_PIPE_CTRL/n15 [0]),
    .sel(ctrl2bpu_rs2ren),
    .o(\u_PIPE_CTRL/rs2_match ));  // ../RTL/core/pipe_ctrl.v(45)
  and \u_PIPE_CTRL/u1  (\u_PIPE_CTRL/n1 [0], ctrl2exu_rdwen0, \u_PIPE_CTRL/n0 );  // ../RTL/core/pipe_ctrl.v(42)
  or \u_PIPE_CTRL/u10  (\u_PIPE_CTRL/read_after_write , \u_PIPE_CTRL/rs1_match , \u_PIPE_CTRL/rs2_match );  // ../RTL/core/pipe_ctrl.v(51)
  or \u_PIPE_CTRL/u11  (\u_PIPE_CTRL/n16 , ctrl2exu_resource_match, \u_PIPE_CTRL/read_after_write );  // ../RTL/core/pipe_ctrl.v(54)
  or \u_PIPE_CTRL/u12  (ctrl2bpu_wait, \u_PIPE_CTRL/n16 , ctrl2wb_match);  // ../RTL/core/pipe_ctrl.v(54)
  or \u_PIPE_CTRL/u14  (ctrl2dis_wait, ctrl2exu_resource_match, ctrl2wb_match);  // ../RTL/core/pipe_ctrl.v(57)
  or \u_PIPE_CTRL/u15  (\u_PIPE_CTRL/n15 [0], \u_PIPE_CTRL/n12 [0], \u_PIPE_CTRL/n14 [0]);  // ../RTL/core/pipe_ctrl.v(46)
  AL_MUX \u_PIPE_CTRL/u16  (
    .i0(\u_PIPE_CTRL/read_after_write ),
    .i1(1'b0),
    .sel(ctrl2dis_wait),
    .o(ctrl2dis_flush));  // ../RTL/core/pipe_ctrl.v(61)
  and \u_PIPE_CTRL/u2  (\u_PIPE_CTRL/n3 [0], ctrl2exu_rdwen1, \u_PIPE_CTRL/n2 );  // ../RTL/core/pipe_ctrl.v(43)
  or \u_PIPE_CTRL/u3  (\u_PIPE_CTRL/n4 [0], \u_PIPE_CTRL/n1 [0], \u_PIPE_CTRL/n3 [0]);  // ../RTL/core/pipe_ctrl.v(42)
  and \u_PIPE_CTRL/u4  (\u_PIPE_CTRL/n6 [0], ctrl2exu_rdwen2, \u_PIPE_CTRL/n5 );  // ../RTL/core/pipe_ctrl.v(44)
  or \u_PIPE_CTRL/u5  (\u_PIPE_CTRL/n7 [0], \u_PIPE_CTRL/n4 [0], \u_PIPE_CTRL/n6 [0]);  // ../RTL/core/pipe_ctrl.v(42)
  and \u_PIPE_CTRL/u6  (\u_PIPE_CTRL/n9 [0], ctrl2exu_rdwen0, \u_PIPE_CTRL/n8 );  // ../RTL/core/pipe_ctrl.v(46)
  and \u_PIPE_CTRL/u7  (\u_PIPE_CTRL/n11 [0], ctrl2exu_rdwen1, \u_PIPE_CTRL/n10 );  // ../RTL/core/pipe_ctrl.v(47)
  or \u_PIPE_CTRL/u8  (\u_PIPE_CTRL/n12 [0], \u_PIPE_CTRL/n9 [0], \u_PIPE_CTRL/n11 [0]);  // ../RTL/core/pipe_ctrl.v(46)
  and \u_PIPE_CTRL/u9  (\u_PIPE_CTRL/n14 [0], ctrl2exu_rdwen2, \u_PIPE_CTRL/n13 );  // ../RTL/core/pipe_ctrl.v(48)
  and \u_WB/mux10_b0_sel_is_2  (\u_WB/mux10_b0_sel_is_2_o , i_rstn, \u_WB/n1 );
  binary_mux_s1_w1 \u_WB/mux12_b0  (
    .i0(\u_WB/rdidx0 [0]),
    .i1(\u_WB/rdidx1 [0]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n34 [0]));  // ../RTL/core/wb.v(89)
  binary_mux_s1_w1 \u_WB/mux12_b1  (
    .i0(\u_WB/rdidx0 [1]),
    .i1(\u_WB/rdidx1 [1]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n34 [1]));  // ../RTL/core/wb.v(89)
  binary_mux_s1_w1 \u_WB/mux12_b2  (
    .i0(\u_WB/rdidx0 [2]),
    .i1(\u_WB/rdidx1 [2]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n34 [2]));  // ../RTL/core/wb.v(89)
  binary_mux_s1_w1 \u_WB/mux12_b3  (
    .i0(\u_WB/rdidx0 [3]),
    .i1(\u_WB/rdidx1 [3]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n34 [3]));  // ../RTL/core/wb.v(89)
  binary_mux_s1_w1 \u_WB/mux12_b4  (
    .i0(\u_WB/rdidx0 [4]),
    .i1(\u_WB/rdidx1 [4]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n34 [4]));  // ../RTL/core/wb.v(89)
  binary_mux_s1_w1 \u_WB/mux13_b0  (
    .i0(\u_WB/n34 [0]),
    .i1(\u_WB/rdidx2 [0]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdidx[0]));  // ../RTL/core/wb.v(89)
  binary_mux_s1_w1 \u_WB/mux13_b1  (
    .i0(\u_WB/n34 [1]),
    .i1(\u_WB/rdidx2 [1]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdidx[1]));  // ../RTL/core/wb.v(89)
  binary_mux_s1_w1 \u_WB/mux13_b2  (
    .i0(\u_WB/n34 [2]),
    .i1(\u_WB/rdidx2 [2]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdidx[2]));  // ../RTL/core/wb.v(89)
  binary_mux_s1_w1 \u_WB/mux13_b3  (
    .i0(\u_WB/n34 [3]),
    .i1(\u_WB/rdidx2 [3]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdidx[3]));  // ../RTL/core/wb.v(89)
  binary_mux_s1_w1 \u_WB/mux13_b4  (
    .i0(\u_WB/n34 [4]),
    .i1(\u_WB/rdidx2 [4]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdidx[4]));  // ../RTL/core/wb.v(89)
  binary_mux_s1_w1 \u_WB/mux14_b0  (
    .i0(\u_WB/rdwdata0 [0]),
    .i1(\u_WB/rdwdata1 [0]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [0]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b1  (
    .i0(\u_WB/rdwdata0 [1]),
    .i1(\u_WB/rdwdata1 [1]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [1]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b10  (
    .i0(\u_WB/rdwdata0 [10]),
    .i1(\u_WB/rdwdata1 [10]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [10]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b11  (
    .i0(\u_WB/rdwdata0 [11]),
    .i1(\u_WB/rdwdata1 [11]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [11]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b12  (
    .i0(\u_WB/rdwdata0 [12]),
    .i1(\u_WB/rdwdata1 [12]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [12]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b13  (
    .i0(\u_WB/rdwdata0 [13]),
    .i1(\u_WB/rdwdata1 [13]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [13]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b14  (
    .i0(\u_WB/rdwdata0 [14]),
    .i1(\u_WB/rdwdata1 [14]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [14]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b15  (
    .i0(\u_WB/rdwdata0 [15]),
    .i1(\u_WB/rdwdata1 [15]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [15]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b16  (
    .i0(\u_WB/rdwdata0 [16]),
    .i1(\u_WB/rdwdata1 [16]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [16]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b17  (
    .i0(\u_WB/rdwdata0 [17]),
    .i1(\u_WB/rdwdata1 [17]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [17]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b18  (
    .i0(\u_WB/rdwdata0 [18]),
    .i1(\u_WB/rdwdata1 [18]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [18]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b19  (
    .i0(\u_WB/rdwdata0 [19]),
    .i1(\u_WB/rdwdata1 [19]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [19]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b2  (
    .i0(\u_WB/rdwdata0 [2]),
    .i1(\u_WB/rdwdata1 [2]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [2]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b20  (
    .i0(\u_WB/rdwdata0 [20]),
    .i1(\u_WB/rdwdata1 [20]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [20]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b21  (
    .i0(\u_WB/rdwdata0 [21]),
    .i1(\u_WB/rdwdata1 [21]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [21]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b22  (
    .i0(\u_WB/rdwdata0 [22]),
    .i1(\u_WB/rdwdata1 [22]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [22]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b23  (
    .i0(\u_WB/rdwdata0 [23]),
    .i1(\u_WB/rdwdata1 [23]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [23]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b24  (
    .i0(\u_WB/rdwdata0 [24]),
    .i1(\u_WB/rdwdata1 [24]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [24]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b25  (
    .i0(\u_WB/rdwdata0 [25]),
    .i1(\u_WB/rdwdata1 [25]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [25]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b26  (
    .i0(\u_WB/rdwdata0 [26]),
    .i1(\u_WB/rdwdata1 [26]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [26]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b27  (
    .i0(\u_WB/rdwdata0 [27]),
    .i1(\u_WB/rdwdata1 [27]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [27]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b28  (
    .i0(\u_WB/rdwdata0 [28]),
    .i1(\u_WB/rdwdata1 [28]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [28]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b29  (
    .i0(\u_WB/rdwdata0 [29]),
    .i1(\u_WB/rdwdata1 [29]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [29]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b3  (
    .i0(\u_WB/rdwdata0 [3]),
    .i1(\u_WB/rdwdata1 [3]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [3]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b30  (
    .i0(\u_WB/rdwdata0 [30]),
    .i1(\u_WB/rdwdata1 [30]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [30]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b31  (
    .i0(\u_WB/rdwdata0 [31]),
    .i1(\u_WB/rdwdata1 [31]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [31]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b4  (
    .i0(\u_WB/rdwdata0 [4]),
    .i1(\u_WB/rdwdata1 [4]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [4]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b5  (
    .i0(\u_WB/rdwdata0 [5]),
    .i1(\u_WB/rdwdata1 [5]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [5]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b6  (
    .i0(\u_WB/rdwdata0 [6]),
    .i1(\u_WB/rdwdata1 [6]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [6]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b7  (
    .i0(\u_WB/rdwdata0 [7]),
    .i1(\u_WB/rdwdata1 [7]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [7]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b8  (
    .i0(\u_WB/rdwdata0 [8]),
    .i1(\u_WB/rdwdata1 [8]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [8]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux14_b9  (
    .i0(\u_WB/rdwdata0 [9]),
    .i1(\u_WB/rdwdata1 [9]),
    .sel(\u_WB/rdwen1 ),
    .o(\u_WB/n35 [9]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b0  (
    .i0(\u_WB/n35 [0]),
    .i1(\u_WB/rdwdata2 [0]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[0]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b1  (
    .i0(\u_WB/n35 [1]),
    .i1(\u_WB/rdwdata2 [1]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[1]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b10  (
    .i0(\u_WB/n35 [10]),
    .i1(\u_WB/rdwdata2 [10]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[10]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b11  (
    .i0(\u_WB/n35 [11]),
    .i1(\u_WB/rdwdata2 [11]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[11]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b12  (
    .i0(\u_WB/n35 [12]),
    .i1(\u_WB/rdwdata2 [12]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[12]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b13  (
    .i0(\u_WB/n35 [13]),
    .i1(\u_WB/rdwdata2 [13]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[13]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b14  (
    .i0(\u_WB/n35 [14]),
    .i1(\u_WB/rdwdata2 [14]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[14]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b15  (
    .i0(\u_WB/n35 [15]),
    .i1(\u_WB/rdwdata2 [15]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[15]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b16  (
    .i0(\u_WB/n35 [16]),
    .i1(\u_WB/rdwdata2 [16]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[16]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b17  (
    .i0(\u_WB/n35 [17]),
    .i1(\u_WB/rdwdata2 [17]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[17]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b18  (
    .i0(\u_WB/n35 [18]),
    .i1(\u_WB/rdwdata2 [18]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[18]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b19  (
    .i0(\u_WB/n35 [19]),
    .i1(\u_WB/rdwdata2 [19]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[19]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b2  (
    .i0(\u_WB/n35 [2]),
    .i1(\u_WB/rdwdata2 [2]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[2]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b20  (
    .i0(\u_WB/n35 [20]),
    .i1(\u_WB/rdwdata2 [20]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[20]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b21  (
    .i0(\u_WB/n35 [21]),
    .i1(\u_WB/rdwdata2 [21]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[21]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b22  (
    .i0(\u_WB/n35 [22]),
    .i1(\u_WB/rdwdata2 [22]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[22]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b23  (
    .i0(\u_WB/n35 [23]),
    .i1(\u_WB/rdwdata2 [23]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[23]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b24  (
    .i0(\u_WB/n35 [24]),
    .i1(\u_WB/rdwdata2 [24]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[24]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b25  (
    .i0(\u_WB/n35 [25]),
    .i1(\u_WB/rdwdata2 [25]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[25]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b26  (
    .i0(\u_WB/n35 [26]),
    .i1(\u_WB/rdwdata2 [26]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[26]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b27  (
    .i0(\u_WB/n35 [27]),
    .i1(\u_WB/rdwdata2 [27]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[27]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b28  (
    .i0(\u_WB/n35 [28]),
    .i1(\u_WB/rdwdata2 [28]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[28]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b29  (
    .i0(\u_WB/n35 [29]),
    .i1(\u_WB/rdwdata2 [29]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[29]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b3  (
    .i0(\u_WB/n35 [3]),
    .i1(\u_WB/rdwdata2 [3]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[3]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b30  (
    .i0(\u_WB/n35 [30]),
    .i1(\u_WB/rdwdata2 [30]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[30]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b31  (
    .i0(\u_WB/n35 [31]),
    .i1(\u_WB/rdwdata2 [31]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[31]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b4  (
    .i0(\u_WB/n35 [4]),
    .i1(\u_WB/rdwdata2 [4]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[4]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b5  (
    .i0(\u_WB/n35 [5]),
    .i1(\u_WB/rdwdata2 [5]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[5]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b6  (
    .i0(\u_WB/n35 [6]),
    .i1(\u_WB/rdwdata2 [6]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[6]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b7  (
    .i0(\u_WB/n35 [7]),
    .i1(\u_WB/rdwdata2 [7]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[7]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b8  (
    .i0(\u_WB/n35 [8]),
    .i1(\u_WB/rdwdata2 [8]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[8]));  // ../RTL/core/wb.v(90)
  binary_mux_s1_w1 \u_WB/mux15_b9  (
    .i0(\u_WB/n35 [9]),
    .i1(\u_WB/rdwdata2 [9]),
    .sel(\u_WB/rdwen2 ),
    .o(wb_rdwdata[9]));  // ../RTL/core/wb.v(90)
  AL_DFF_X \u_WB/o_exu_taken_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_WB/n37 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_taken_gen));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/rdwen0_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_WB/n2 ),
    .en(\u_WB/n1 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwen0 ));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/rdwen1_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_WB/n15 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwen1 ));  // ../RTL/core/wb.v(57)
  not \u_WB/rdwen2_inv  (\u_WB/rdwen2_neg , \u_WB/rdwen2 );
  AL_DFF_X \u_WB/rdwen2_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_WB/n16 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwen2 ));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg0_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx0[0]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx0 [0]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg0_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx0[1]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx0 [1]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg0_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx0[2]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx0 [2]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg0_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx0[3]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx0 [3]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg0_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx0[4]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx0 [4]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg1_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx1[0]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx1 [0]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg1_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx1[1]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx1 [1]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg1_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx1[2]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx1 [2]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg1_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx1[3]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx1 [3]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg1_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx1[4]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx1 [4]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg2_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx2[0]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx2 [0]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg2_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx2[1]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx2 [1]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg2_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx2[2]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx2 [2]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg2_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx2[3]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx2 [3]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg2_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdidx2[4]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdidx2 [4]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[0]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [0]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[1]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [1]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[10]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [10]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[11]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [11]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[12]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [12]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[13]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [13]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[14]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [14]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[15]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [15]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[16]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [16]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[17]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [17]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[18]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [18]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[19]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [19]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[2]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [2]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[20]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [20]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[21]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [21]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[22]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [22]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[23]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [23]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[24]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [24]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[25]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [25]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[26]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [26]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[27]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [27]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[28]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [28]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[29]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [29]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[3]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [3]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[30]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [30]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[31]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [31]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[4]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [4]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[5]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [5]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[6]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [6]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[7]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [7]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[8]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [8]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg3_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata0[9]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata0 [9]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[0]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [0]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[1]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [1]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[10]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [10]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[11]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [11]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[12]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [12]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[13]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [13]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[14]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [14]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[15]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [15]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[16]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [16]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[17]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [17]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[18]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [18]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[19]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [19]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[2]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [2]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[20]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [20]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[21]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [21]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[22]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [22]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[23]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [23]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[24]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [24]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[25]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [25]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[26]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [26]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[27]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [27]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[28]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [28]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[29]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [29]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[3]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [3]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[30]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [30]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[31]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [31]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[4]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [4]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[5]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [5]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[6]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [6]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[7]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [7]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[8]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [8]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg4_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata1[9]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata1 [9]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[0]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [0]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[1]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [1]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[10]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [10]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[11]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [11]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[12]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [12]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[13]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [13]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[14]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [14]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[15]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [15]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[16]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [16]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[17]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [17]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[18]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [18]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[19]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [19]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[2]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [2]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[20]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [20]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[21]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [21]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[22]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [22]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[23]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [23]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[24]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [24]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[25]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [25]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[26]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [26]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[27]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [27]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[28]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [28]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[29]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [29]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[3]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [3]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[30]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [30]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[31]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [31]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[4]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [4]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[5]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [5]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[6]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [6]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[7]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [7]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[8]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [8]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg5_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_rdwdata2[9]),
    .en(\u_WB/mux10_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_WB/rdwdata2 [9]));  // ../RTL/core/wb.v(57)
  AL_DFF_X \u_WB/reg6_b0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[0]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b1  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[1]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b10  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[10]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b11  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[11]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b12  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[12]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b13  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[13]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b14  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[14]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b15  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[15]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b16  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[16]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b17  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[17]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b18  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[18]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b19  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[19]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b2  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[2]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b20  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[20]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b21  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[21]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b22  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[22]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b23  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[23]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b24  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[24]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b25  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[25]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b26  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[26]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b27  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[27]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b28  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[28]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b29  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[29]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b3  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[3]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b30  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[30]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b31  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[31]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b4  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[4]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b5  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[5]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b6  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[6]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b7  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[7]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b8  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[8]));  // ../RTL/core/wb.v(94)
  AL_DFF_X \u_WB/reg6_b9  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(exu_jaddr[9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(exu_jaddr_gen[9]));  // ../RTL/core/wb.v(94)
  AL_MUX \u_WB/u10  (
    .i0(exu_rdwen2),
    .i1(1'b0),
    .sel(\u_WB/n7 ),
    .o(\u_WB/n8 ));  // ../RTL/core/wb.v(65)
  and \u_WB/u13_sel_is_2  (\u_WB/u13_sel_is_2_o , \u_WB/rdwen2_neg , \u_WB/rdwen1 );
  AL_MUX \u_WB/u14  (
    .i0(\u_WB/rdwen2 ),
    .i1(1'b0),
    .sel(\u_WB/u14_sel_is_3_o ),
    .o(\u_WB/n12 ));
  and \u_WB/u14_sel_is_3  (\u_WB/u14_sel_is_3_o , ctrl2wb_match, \u_WB/rdwen2 );
  AL_MUX \u_WB/u15  (
    .i0(\u_WB/rdwen1 ),
    .i1(1'b0),
    .sel(\u_WB/u15_sel_is_3_o ),
    .o(\u_WB/n13 ));
  and \u_WB/u15_sel_is_3  (\u_WB/u15_sel_is_3_o , ctrl2wb_match, \u_WB/u13_sel_is_2_o );
  AL_MUX \u_WB/u17  (
    .i0(\u_WB/n13 ),
    .i1(\u_WB/n5 ),
    .sel(\u_WB/n1 ),
    .o(\u_WB/n15 ));  // ../RTL/core/wb.v(62)
  AL_MUX \u_WB/u18  (
    .i0(\u_WB/n12 ),
    .i1(\u_WB/n8 ),
    .sel(\u_WB/n1 ),
    .o(\u_WB/n16 ));  // ../RTL/core/wb.v(62)
  and \u_WB/u19  (\u_WB/n29 , \u_WB/rdwen0 , \u_WB/rdwen1 );  // ../RTL/core/wb.v(86)
  not \u_WB/u2  (\u_WB/n0 , ctrl2wb_match);  // ../RTL/core/wb.v(62)
  and \u_WB/u20  (\u_WB/n30 , \u_WB/rdwen0 , \u_WB/rdwen2 );  // ../RTL/core/wb.v(86)
  or \u_WB/u21  (\u_WB/n31 , \u_WB/n29 , \u_WB/n30 );  // ../RTL/core/wb.v(86)
  and \u_WB/u22  (\u_WB/n32 , \u_WB/rdwen1 , \u_WB/rdwen2 );  // ../RTL/core/wb.v(86)
  or \u_WB/u23  (ctrl2wb_match, \u_WB/n31 , \u_WB/n32 );  // ../RTL/core/wb.v(86)
  or \u_WB/u24  (\u_WB/n33 , \u_WB/rdwen0 , \u_WB/rdwen1 );  // ../RTL/core/wb.v(87)
  or \u_WB/u25  (wb_rdwen, \u_WB/n33 , \u_WB/rdwen2 );  // ../RTL/core/wb.v(87)
  AL_MUX \u_WB/u26  (
    .i0(exu_taken),
    .i1(1'b0),
    .sel(exu_taken_gen),
    .o(\u_WB/n37 ));  // ../RTL/core/wb.v(99)
  or \u_WB/u3  (\u_WB/n1 , \u_WB/n0 , exu_taken_gen);  // ../RTL/core/wb.v(62)
  AL_MUX \u_WB/u4  (
    .i0(exu_rdwen0),
    .i1(1'b0),
    .sel(exu_taken_gen),
    .o(\u_WB/n2 ));  // ../RTL/core/wb.v(63)
  not \u_WB/u5  (\u_WB/n3 , exu_rdwen1);  // ../RTL/core/wb.v(64)
  and \u_WB/u6  (\u_WB/n4 , exu_taken_gen, \u_WB/n3 );  // ../RTL/core/wb.v(64)
  AL_MUX \u_WB/u7  (
    .i0(exu_rdwen1),
    .i1(1'b0),
    .sel(\u_WB/n4 ),
    .o(\u_WB/n5 ));  // ../RTL/core/wb.v(64)
  not \u_WB/u8  (\u_WB/n6 , exu_rdwen2);  // ../RTL/core/wb.v(65)
  and \u_WB/u9  (\u_WB/n7 , exu_taken_gen, \u_WB/n6 );  // ../RTL/core/wb.v(65)

endmodule 

module BPU  // ../RTL/core/bpu.v(14)
  (
  i_clk,
  i_data,
  i_data_vld,
  i_flush,
  i_iaddr,
  i_rd_wdata,
  i_rdidx,
  i_rdwen,
  i_rstn,
  i_stop,
  o_bpu_jaddr,
  o_bpu_rs1idx,
  o_bpu_rs1ren,
  o_bpu_rs2idx,
  o_bpu_rs2ren,
  o_bpu_taken,
  o_csr_ren,
  o_csr_zimm,
  o_csridx,
  o_decinfo,
  o_decinfo_grp,
  o_exu_op1,
  o_exu_op2,
  o_iaddr,
  o_imm,
  o_inst_vld,
  o_rdidx,
  o_rdwen,
  o_rs2rdata
  );

  input i_clk;  // ../RTL/core/bpu.v(15)
  input [31:0] i_data;  // ../RTL/core/bpu.v(24)
  input i_data_vld;  // ../RTL/core/bpu.v(22)
  input i_flush;  // ../RTL/core/bpu.v(19)
  input [31:0] i_iaddr;  // ../RTL/core/bpu.v(23)
  input [31:0] i_rd_wdata;  // ../RTL/core/bpu.v(35)
  input [4:0] i_rdidx;  // ../RTL/core/bpu.v(34)
  input i_rdwen;  // ../RTL/core/bpu.v(33)
  input i_rstn;  // ../RTL/core/bpu.v(16)
  input i_stop;  // ../RTL/core/bpu.v(18)
  output [31:0] o_bpu_jaddr;  // ../RTL/core/bpu.v(39)
  output [4:0] o_bpu_rs1idx;  // ../RTL/core/bpu.v(28)
  output o_bpu_rs1ren;  // ../RTL/core/bpu.v(27)
  output [4:0] o_bpu_rs2idx;  // ../RTL/core/bpu.v(30)
  output o_bpu_rs2ren;  // ../RTL/core/bpu.v(29)
  output o_bpu_taken;  // ../RTL/core/bpu.v(38)
  output o_csr_ren;  // ../RTL/core/bpu.v(50)
  output [31:0] o_csr_zimm;  // ../RTL/core/bpu.v(52)
  output [11:0] o_csridx;  // ../RTL/core/bpu.v(51)
  output [9:0] o_decinfo;  // ../RTL/core/bpu.v(55)
  output [5:0] o_decinfo_grp;  // ../RTL/core/bpu.v(54)
  output [31:0] o_exu_op1;  // ../RTL/core/bpu.v(43)
  output [31:0] o_exu_op2;  // ../RTL/core/bpu.v(44)
  output [31:0] o_iaddr;  // ../RTL/core/bpu.v(56)
  output [31:0] o_imm;  // ../RTL/core/bpu.v(46)
  output o_inst_vld;  // ../RTL/core/bpu.v(42)
  output [4:0] o_rdidx;  // ../RTL/core/bpu.v(48)
  output o_rdwen;  // ../RTL/core/bpu.v(47)
  output [31:0] o_rs2rdata;  // ../RTL/core/bpu.v(45)

  wire [31:0] bp_imm;  // ../RTL/core/bpu.v(105)
  wire [31:0] rs1_rdata;  // ../RTL/core/bpu.v(109)
  wire [31:0] \u_BPU_BP/n2 ;
  wire [31:0] \u_BPU_BP/n3 ;
  wire [31:0] \u_BPU_BP/n4 ;
  wire [9:0] \u_DECODE/aluinfo ;  // ../RTL/core/decode.v(261)
  wire [9:0] \u_DECODE/bjuinfo ;  // ../RTL/core/decode.v(287)
  wire [31:0] \u_DECODE/inst_opimm_imm ;  // ../RTL/core/decode.v(202)
  wire [9:0] \u_DECODE/lsuinfo ;  // ../RTL/core/decode.v(278)
  wire [31:0] \u_DECODE/n22 ;
  wire [31:0] \u_DECODE/n23 ;
  wire [31:0] \u_DECODE/n24 ;
  wire [31:0] \u_DECODE/n25 ;
  wire [31:0] \u_DECODE/n26 ;
  wire [31:0] \u_DECODE/n27 ;
  wire [31:0] \u_DECODE/n28 ;
  wire [31:0] \u_DECODE/n29 ;
  wire [31:0] \u_DECODE/n4 ;
  wire [31:0] \u_DECODE/n5 ;
  wire [31:0] \u_DECODE/n57 ;
  wire [31:0] \u_DECODE/n6 ;
  wire [9:0] \u_DECODE/n65 ;
  wire [9:0] \u_DECODE/n66 ;
  wire [9:0] \u_DECODE/n67 ;
  wire [9:0] \u_DECODE/n68 ;
  wire [9:0] \u_DECODE/n69 ;
  wire [31:0] \u_DECODE/n7 ;
  wire [9:0] \u_DECODE/n70 ;
  wire [9:0] \u_DECODE/n71 ;
  wire [9:0] \u_DECODE/n72 ;
  wire [9:0] \u_DECODE/scuinfo ;  // ../RTL/core/decode.v(320)
  wire bpu_bflag;  // ../RTL/core/bpu.v(100)
  wire inst_bxx;  // ../RTL/core/bpu.v(103)
  wire inst_jal;  // ../RTL/core/bpu.v(101)
  wire inst_jalr;  // ../RTL/core/bpu.v(102)
  wire jalr_rs1ren;  // ../RTL/core/bpu.v(162)
  wire n0;
  wire n1;
  wire rs1ren;  // ../RTL/core/bpu.v(107)
  wire rs1topc;  // ../RTL/core/bpu.v(114)
  wire rs2ren;  // ../RTL/core/bpu.v(110)
  wire rs2toimm;  // ../RTL/core/bpu.v(115)
  wire \u_BPU_BP/n0 ;
  wire \u_BPU_BP/n1 ;
  wire \u_DECODE/func7_0000000 ;  // ../RTL/core/decode.v(107)
  wire \u_DECODE/func7_0000001 ;  // ../RTL/core/decode.v(109)
  wire \u_DECODE/func7_0100000 ;  // ../RTL/core/decode.v(108)
  wire \u_DECODE/func_000 ;  // ../RTL/core/decode.v(97)
  wire \u_DECODE/func_001 ;  // ../RTL/core/decode.v(98)
  wire \u_DECODE/func_010 ;  // ../RTL/core/decode.v(99)
  wire \u_DECODE/func_011 ;  // ../RTL/core/decode.v(100)
  wire \u_DECODE/func_100 ;  // ../RTL/core/decode.v(101)
  wire \u_DECODE/func_101 ;  // ../RTL/core/decode.v(102)
  wire \u_DECODE/func_110 ;  // ../RTL/core/decode.v(103)
  wire \u_DECODE/func_111 ;  // ../RTL/core/decode.v(104)
  wire \u_DECODE/inst_add ;  // ../RTL/core/decode.v(150)
  wire \u_DECODE/inst_addi ;  // ../RTL/core/decode.v(140)
  wire \u_DECODE/inst_and ;  // ../RTL/core/decode.v(159)
  wire \u_DECODE/inst_andi ;  // ../RTL/core/decode.v(145)
  wire \u_DECODE/inst_beq ;  // ../RTL/core/decode.v(123)
  wire \u_DECODE/inst_bge ;  // ../RTL/core/decode.v(126)
  wire \u_DECODE/inst_bgeu ;  // ../RTL/core/decode.v(128)
  wire \u_DECODE/inst_blt ;  // ../RTL/core/decode.v(125)
  wire \u_DECODE/inst_bltu ;  // ../RTL/core/decode.v(127)
  wire \u_DECODE/inst_bne ;  // ../RTL/core/decode.v(124)
  wire \u_DECODE/inst_csrrc ;  // ../RTL/core/decode.v(168)
  wire \u_DECODE/inst_csrrci ;  // ../RTL/core/decode.v(171)
  wire \u_DECODE/inst_csrrs ;  // ../RTL/core/decode.v(167)
  wire \u_DECODE/inst_csrrsi ;  // ../RTL/core/decode.v(170)
  wire \u_DECODE/inst_csrrw ;  // ../RTL/core/decode.v(166)
  wire \u_DECODE/inst_csrrwi ;  // ../RTL/core/decode.v(169)
  wire \u_DECODE/inst_div ;  // ../RTL/core/decode.v(178)
  wire \u_DECODE/inst_divu ;  // ../RTL/core/decode.v(179)
  wire \u_DECODE/inst_ebreak ;  // ../RTL/core/decode.v(165)
  wire \u_DECODE/inst_ecall ;  // ../RTL/core/decode.v(164)
  wire \u_DECODE/inst_mul ;  // ../RTL/core/decode.v(174)
  wire \u_DECODE/inst_mulh ;  // ../RTL/core/decode.v(175)
  wire \u_DECODE/inst_mulhsu ;  // ../RTL/core/decode.v(176)
  wire \u_DECODE/inst_mulhu ;  // ../RTL/core/decode.v(177)
  wire \u_DECODE/inst_or ;  // ../RTL/core/decode.v(158)
  wire \u_DECODE/inst_ori ;  // ../RTL/core/decode.v(144)
  wire \u_DECODE/inst_rem ;  // ../RTL/core/decode.v(180)
  wire \u_DECODE/inst_remu ;  // ../RTL/core/decode.v(181)
  wire \u_DECODE/inst_sll ;  // ../RTL/core/decode.v(152)
  wire \u_DECODE/inst_slli ;  // ../RTL/core/decode.v(146)
  wire \u_DECODE/inst_slt ;  // ../RTL/core/decode.v(153)
  wire \u_DECODE/inst_slti ;  // ../RTL/core/decode.v(141)
  wire \u_DECODE/inst_sltiu ;  // ../RTL/core/decode.v(142)
  wire \u_DECODE/inst_sltu ;  // ../RTL/core/decode.v(154)
  wire \u_DECODE/inst_sra ;  // ../RTL/core/decode.v(157)
  wire \u_DECODE/inst_srai ;  // ../RTL/core/decode.v(148)
  wire \u_DECODE/inst_srl ;  // ../RTL/core/decode.v(156)
  wire \u_DECODE/inst_srli ;  // ../RTL/core/decode.v(147)
  wire \u_DECODE/inst_sub ;  // ../RTL/core/decode.v(151)
  wire \u_DECODE/inst_xor ;  // ../RTL/core/decode.v(155)
  wire \u_DECODE/inst_xori ;  // ../RTL/core/decode.v(143)
  wire \u_DECODE/n0 ;
  wire \u_DECODE/n1 ;
  wire \u_DECODE/n10 ;
  wire \u_DECODE/n11 ;
  wire \u_DECODE/n12 ;
  wire \u_DECODE/n13 ;
  wire \u_DECODE/n14 ;
  wire \u_DECODE/n15 ;
  wire \u_DECODE/n16 ;
  wire \u_DECODE/n17 ;
  wire \u_DECODE/n18 ;
  wire \u_DECODE/n19 ;
  wire \u_DECODE/n2 ;
  wire \u_DECODE/n20 ;
  wire \u_DECODE/n21 ;
  wire \u_DECODE/n3 ;
  wire \u_DECODE/n30 ;
  wire \u_DECODE/n31 ;
  wire \u_DECODE/n32 ;
  wire \u_DECODE/n33 ;
  wire \u_DECODE/n34 ;
  wire \u_DECODE/n35 ;
  wire \u_DECODE/n36 ;
  wire \u_DECODE/n38 ;
  wire \u_DECODE/n39 ;
  wire \u_DECODE/n40 ;
  wire \u_DECODE/n41 ;
  wire \u_DECODE/n42 ;
  wire \u_DECODE/n43 ;
  wire \u_DECODE/n44 ;
  wire \u_DECODE/n45 ;
  wire \u_DECODE/n46 ;
  wire \u_DECODE/n47 ;
  wire \u_DECODE/n48 ;
  wire \u_DECODE/n49 ;
  wire \u_DECODE/n50 ;
  wire \u_DECODE/n51 ;
  wire \u_DECODE/n52 ;
  wire \u_DECODE/n53 ;
  wire \u_DECODE/n54 ;
  wire \u_DECODE/n55 ;
  wire \u_DECODE/n56 ;
  wire \u_DECODE/n58 ;
  wire \u_DECODE/n59 ;
  wire \u_DECODE/n60 ;
  wire \u_DECODE/n61 ;
  wire \u_DECODE/n62 ;
  wire \u_DECODE/n63 ;
  wire \u_DECODE/n64 ;
  wire \u_DECODE/n8 ;
  wire \u_DECODE/n9 ;
  wire \u_DECODE/opc_load ;  // ../RTL/core/decode.v(89)
  wire \u_DECODE/opc_lui ;  // ../RTL/core/decode.v(84)
  wire \u_DECODE/opc_op ;  // ../RTL/core/decode.v(92)
  wire \u_DECODE/opc_opimm ;  // ../RTL/core/decode.v(91)
  wire \u_DECODE/opc_rv32 ;  // ../RTL/core/decode.v(67)
  wire \u_DECODE/opc_store ;  // ../RTL/core/decode.v(90)
  wire \u_DECODE/type_i_imm_000000000000 ;  // ../RTL/core/decode.v(112)
  wire \u_DECODE/type_i_imm_000000000001 ;  // ../RTL/core/decode.v(113)

  assign o_iaddr[31] = i_iaddr[31];
  assign o_iaddr[30] = i_iaddr[30];
  assign o_iaddr[29] = i_iaddr[29];
  assign o_iaddr[28] = i_iaddr[28];
  assign o_iaddr[27] = i_iaddr[27];
  assign o_iaddr[26] = i_iaddr[26];
  assign o_iaddr[25] = i_iaddr[25];
  assign o_iaddr[24] = i_iaddr[24];
  assign o_iaddr[23] = i_iaddr[23];
  assign o_iaddr[22] = i_iaddr[22];
  assign o_iaddr[21] = i_iaddr[21];
  assign o_iaddr[20] = i_iaddr[20];
  assign o_iaddr[19] = i_iaddr[19];
  assign o_iaddr[18] = i_iaddr[18];
  assign o_iaddr[17] = i_iaddr[17];
  assign o_iaddr[16] = i_iaddr[16];
  assign o_iaddr[15] = i_iaddr[15];
  assign o_iaddr[14] = i_iaddr[14];
  assign o_iaddr[13] = i_iaddr[13];
  assign o_iaddr[12] = i_iaddr[12];
  assign o_iaddr[11] = i_iaddr[11];
  assign o_iaddr[10] = i_iaddr[10];
  assign o_iaddr[9] = i_iaddr[9];
  assign o_iaddr[8] = i_iaddr[8];
  assign o_iaddr[7] = i_iaddr[7];
  assign o_iaddr[6] = i_iaddr[6];
  assign o_iaddr[5] = i_iaddr[5];
  assign o_iaddr[4] = i_iaddr[4];
  assign o_iaddr[3] = i_iaddr[3];
  assign o_iaddr[2] = i_iaddr[2];
  assign o_iaddr[1] = i_iaddr[1];
  assign o_iaddr[0] = i_iaddr[0];
  assign o_bpu_rs1idx[4] = i_data[19];
  assign o_bpu_rs1idx[3] = i_data[18];
  assign o_bpu_rs1idx[2] = i_data[17];
  assign o_bpu_rs1idx[1] = i_data[16];
  assign o_bpu_rs1idx[0] = i_data[15];
  assign o_bpu_rs2idx[4] = i_data[24];
  assign o_bpu_rs2idx[3] = i_data[23];
  assign o_bpu_rs2idx[2] = i_data[22];
  assign o_bpu_rs2idx[1] = i_data[21];
  assign o_bpu_rs2idx[0] = i_data[20];
  assign o_csr_zimm[31] = 1'b0;
  assign o_csr_zimm[30] = 1'b0;
  assign o_csr_zimm[29] = 1'b0;
  assign o_csr_zimm[28] = 1'b0;
  assign o_csr_zimm[27] = 1'b0;
  assign o_csr_zimm[26] = 1'b0;
  assign o_csr_zimm[25] = 1'b0;
  assign o_csr_zimm[24] = 1'b0;
  assign o_csr_zimm[23] = 1'b0;
  assign o_csr_zimm[22] = 1'b0;
  assign o_csr_zimm[21] = 1'b0;
  assign o_csr_zimm[20] = 1'b0;
  assign o_csr_zimm[19] = 1'b0;
  assign o_csr_zimm[18] = 1'b0;
  assign o_csr_zimm[17] = 1'b0;
  assign o_csr_zimm[16] = 1'b0;
  assign o_csr_zimm[15] = 1'b0;
  assign o_csr_zimm[14] = 1'b0;
  assign o_csr_zimm[13] = 1'b0;
  assign o_csr_zimm[12] = 1'b0;
  assign o_csr_zimm[11] = 1'b0;
  assign o_csr_zimm[10] = 1'b0;
  assign o_csr_zimm[9] = 1'b0;
  assign o_csr_zimm[8] = 1'b0;
  assign o_csr_zimm[7] = 1'b0;
  assign o_csr_zimm[6] = 1'b0;
  assign o_csr_zimm[5] = 1'b0;
  assign o_decinfo[9] = \u_DECODE/n65 [9];
  assign o_decinfo[8] = \u_DECODE/n71 [8];
  assign o_rdidx[4] = i_data[11];
  assign o_rdidx[3] = i_data[10];
  assign o_rdidx[2] = i_data[9];
  assign o_rdidx[1] = i_data[8];
  assign o_rdidx[0] = i_data[7];
  binary_mux_s1_w1 mux0_b0 (
    .i0(rs1_rdata[0]),
    .i1(o_iaddr[0]),
    .sel(rs1topc),
    .o(o_exu_op1[0]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b1 (
    .i0(rs1_rdata[1]),
    .i1(o_iaddr[1]),
    .sel(rs1topc),
    .o(o_exu_op1[1]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b10 (
    .i0(rs1_rdata[10]),
    .i1(o_iaddr[10]),
    .sel(rs1topc),
    .o(o_exu_op1[10]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b11 (
    .i0(rs1_rdata[11]),
    .i1(o_iaddr[11]),
    .sel(rs1topc),
    .o(o_exu_op1[11]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b12 (
    .i0(rs1_rdata[12]),
    .i1(o_iaddr[12]),
    .sel(rs1topc),
    .o(o_exu_op1[12]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b13 (
    .i0(rs1_rdata[13]),
    .i1(o_iaddr[13]),
    .sel(rs1topc),
    .o(o_exu_op1[13]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b14 (
    .i0(rs1_rdata[14]),
    .i1(o_iaddr[14]),
    .sel(rs1topc),
    .o(o_exu_op1[14]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b15 (
    .i0(rs1_rdata[15]),
    .i1(o_iaddr[15]),
    .sel(rs1topc),
    .o(o_exu_op1[15]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b16 (
    .i0(rs1_rdata[16]),
    .i1(o_iaddr[16]),
    .sel(rs1topc),
    .o(o_exu_op1[16]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b17 (
    .i0(rs1_rdata[17]),
    .i1(o_iaddr[17]),
    .sel(rs1topc),
    .o(o_exu_op1[17]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b18 (
    .i0(rs1_rdata[18]),
    .i1(o_iaddr[18]),
    .sel(rs1topc),
    .o(o_exu_op1[18]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b19 (
    .i0(rs1_rdata[19]),
    .i1(o_iaddr[19]),
    .sel(rs1topc),
    .o(o_exu_op1[19]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b2 (
    .i0(rs1_rdata[2]),
    .i1(o_iaddr[2]),
    .sel(rs1topc),
    .o(o_exu_op1[2]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b20 (
    .i0(rs1_rdata[20]),
    .i1(o_iaddr[20]),
    .sel(rs1topc),
    .o(o_exu_op1[20]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b21 (
    .i0(rs1_rdata[21]),
    .i1(o_iaddr[21]),
    .sel(rs1topc),
    .o(o_exu_op1[21]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b22 (
    .i0(rs1_rdata[22]),
    .i1(o_iaddr[22]),
    .sel(rs1topc),
    .o(o_exu_op1[22]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b23 (
    .i0(rs1_rdata[23]),
    .i1(o_iaddr[23]),
    .sel(rs1topc),
    .o(o_exu_op1[23]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b24 (
    .i0(rs1_rdata[24]),
    .i1(o_iaddr[24]),
    .sel(rs1topc),
    .o(o_exu_op1[24]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b25 (
    .i0(rs1_rdata[25]),
    .i1(o_iaddr[25]),
    .sel(rs1topc),
    .o(o_exu_op1[25]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b26 (
    .i0(rs1_rdata[26]),
    .i1(o_iaddr[26]),
    .sel(rs1topc),
    .o(o_exu_op1[26]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b27 (
    .i0(rs1_rdata[27]),
    .i1(o_iaddr[27]),
    .sel(rs1topc),
    .o(o_exu_op1[27]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b28 (
    .i0(rs1_rdata[28]),
    .i1(o_iaddr[28]),
    .sel(rs1topc),
    .o(o_exu_op1[28]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b29 (
    .i0(rs1_rdata[29]),
    .i1(o_iaddr[29]),
    .sel(rs1topc),
    .o(o_exu_op1[29]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b3 (
    .i0(rs1_rdata[3]),
    .i1(o_iaddr[3]),
    .sel(rs1topc),
    .o(o_exu_op1[3]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b30 (
    .i0(rs1_rdata[30]),
    .i1(o_iaddr[30]),
    .sel(rs1topc),
    .o(o_exu_op1[30]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b31 (
    .i0(rs1_rdata[31]),
    .i1(o_iaddr[31]),
    .sel(rs1topc),
    .o(o_exu_op1[31]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b4 (
    .i0(rs1_rdata[4]),
    .i1(o_iaddr[4]),
    .sel(rs1topc),
    .o(o_exu_op1[4]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b5 (
    .i0(rs1_rdata[5]),
    .i1(o_iaddr[5]),
    .sel(rs1topc),
    .o(o_exu_op1[5]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b6 (
    .i0(rs1_rdata[6]),
    .i1(o_iaddr[6]),
    .sel(rs1topc),
    .o(o_exu_op1[6]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b7 (
    .i0(rs1_rdata[7]),
    .i1(o_iaddr[7]),
    .sel(rs1topc),
    .o(o_exu_op1[7]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b8 (
    .i0(rs1_rdata[8]),
    .i1(o_iaddr[8]),
    .sel(rs1topc),
    .o(o_exu_op1[8]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux0_b9 (
    .i0(rs1_rdata[9]),
    .i1(o_iaddr[9]),
    .sel(rs1topc),
    .o(o_exu_op1[9]));  // ../RTL/core/bpu.v(152)
  binary_mux_s1_w1 mux1_b0 (
    .i0(o_rs2rdata[0]),
    .i1(o_imm[0]),
    .sel(rs2toimm),
    .o(o_exu_op2[0]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b1 (
    .i0(o_rs2rdata[1]),
    .i1(o_imm[1]),
    .sel(rs2toimm),
    .o(o_exu_op2[1]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b10 (
    .i0(o_rs2rdata[10]),
    .i1(o_imm[10]),
    .sel(rs2toimm),
    .o(o_exu_op2[10]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b11 (
    .i0(o_rs2rdata[11]),
    .i1(o_imm[11]),
    .sel(rs2toimm),
    .o(o_exu_op2[11]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b12 (
    .i0(o_rs2rdata[12]),
    .i1(o_imm[12]),
    .sel(rs2toimm),
    .o(o_exu_op2[12]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b13 (
    .i0(o_rs2rdata[13]),
    .i1(o_imm[13]),
    .sel(rs2toimm),
    .o(o_exu_op2[13]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b14 (
    .i0(o_rs2rdata[14]),
    .i1(o_imm[14]),
    .sel(rs2toimm),
    .o(o_exu_op2[14]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b15 (
    .i0(o_rs2rdata[15]),
    .i1(o_imm[15]),
    .sel(rs2toimm),
    .o(o_exu_op2[15]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b16 (
    .i0(o_rs2rdata[16]),
    .i1(o_imm[16]),
    .sel(rs2toimm),
    .o(o_exu_op2[16]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b17 (
    .i0(o_rs2rdata[17]),
    .i1(o_imm[17]),
    .sel(rs2toimm),
    .o(o_exu_op2[17]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b18 (
    .i0(o_rs2rdata[18]),
    .i1(o_imm[18]),
    .sel(rs2toimm),
    .o(o_exu_op2[18]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b19 (
    .i0(o_rs2rdata[19]),
    .i1(o_imm[19]),
    .sel(rs2toimm),
    .o(o_exu_op2[19]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b2 (
    .i0(o_rs2rdata[2]),
    .i1(o_imm[2]),
    .sel(rs2toimm),
    .o(o_exu_op2[2]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b20 (
    .i0(o_rs2rdata[20]),
    .i1(o_imm[20]),
    .sel(rs2toimm),
    .o(o_exu_op2[20]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b21 (
    .i0(o_rs2rdata[21]),
    .i1(o_imm[21]),
    .sel(rs2toimm),
    .o(o_exu_op2[21]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b22 (
    .i0(o_rs2rdata[22]),
    .i1(o_imm[22]),
    .sel(rs2toimm),
    .o(o_exu_op2[22]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b23 (
    .i0(o_rs2rdata[23]),
    .i1(o_imm[23]),
    .sel(rs2toimm),
    .o(o_exu_op2[23]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b24 (
    .i0(o_rs2rdata[24]),
    .i1(o_imm[24]),
    .sel(rs2toimm),
    .o(o_exu_op2[24]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b25 (
    .i0(o_rs2rdata[25]),
    .i1(o_imm[25]),
    .sel(rs2toimm),
    .o(o_exu_op2[25]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b26 (
    .i0(o_rs2rdata[26]),
    .i1(o_imm[26]),
    .sel(rs2toimm),
    .o(o_exu_op2[26]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b27 (
    .i0(o_rs2rdata[27]),
    .i1(o_imm[27]),
    .sel(rs2toimm),
    .o(o_exu_op2[27]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b28 (
    .i0(o_rs2rdata[28]),
    .i1(o_imm[28]),
    .sel(rs2toimm),
    .o(o_exu_op2[28]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b29 (
    .i0(o_rs2rdata[29]),
    .i1(o_imm[29]),
    .sel(rs2toimm),
    .o(o_exu_op2[29]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b3 (
    .i0(o_rs2rdata[3]),
    .i1(o_imm[3]),
    .sel(rs2toimm),
    .o(o_exu_op2[3]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b30 (
    .i0(o_rs2rdata[30]),
    .i1(o_imm[30]),
    .sel(rs2toimm),
    .o(o_exu_op2[30]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b31 (
    .i0(o_rs2rdata[31]),
    .i1(o_imm[31]),
    .sel(rs2toimm),
    .o(o_exu_op2[31]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b4 (
    .i0(o_rs2rdata[4]),
    .i1(o_imm[4]),
    .sel(rs2toimm),
    .o(o_exu_op2[4]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b5 (
    .i0(o_rs2rdata[5]),
    .i1(o_imm[5]),
    .sel(rs2toimm),
    .o(o_exu_op2[5]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b6 (
    .i0(o_rs2rdata[6]),
    .i1(o_imm[6]),
    .sel(rs2toimm),
    .o(o_exu_op2[6]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b7 (
    .i0(o_rs2rdata[7]),
    .i1(o_imm[7]),
    .sel(rs2toimm),
    .o(o_exu_op2[7]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b8 (
    .i0(o_rs2rdata[8]),
    .i1(o_imm[8]),
    .sel(rs2toimm),
    .o(o_exu_op2[8]));  // ../RTL/core/bpu.v(153)
  binary_mux_s1_w1 mux1_b9 (
    .i0(o_rs2rdata[9]),
    .i1(o_imm[9]),
    .sel(rs2toimm),
    .o(o_exu_op2[9]));  // ../RTL/core/bpu.v(153)
  ne_w5 neq0 (
    .i0(i_data[19:15]),
    .i1(5'b00000),
    .o(n1));  // ../RTL/core/bpu.v(162)
  and u12 (o_bpu_rs1ren, i_data_vld, rs1ren);  // ../RTL/core/bpu.v(157)
  and u14 (o_bpu_rs2ren, i_data_vld, rs2ren);  // ../RTL/core/bpu.v(159)
  and u16 (jalr_rs1ren, inst_jalr, n1);  // ../RTL/core/bpu.v(162)
  and u17 (bpu_bflag, inst_bxx, o_bpu_taken);  // ../RTL/core/bpu.v(184)
  not u6 (n0, i_stop);  // ../RTL/core/bpu.v(96)
  and u7 (o_inst_vld, i_data_vld, n0);  // ../RTL/core/bpu.v(96)
  add_pu32_pu32_o32 \u_BPU_BP/add0  (
    .i0(rs1_rdata),
    .i1({bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[19:1],\u_DECODE/n5 [0]}),
    .o(\u_BPU_BP/n2 ));  // ../RTL/core/bpu_bp.v(44)
  add_pu32_pu32_o32 \u_BPU_BP/add1  (
    .i0(o_iaddr),
    .i1({bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[31],bp_imm[19:1],\u_DECODE/n5 [0]}),
    .o(\u_BPU_BP/n4 ));  // ../RTL/core/bpu_bp.v(45)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b0  (
    .i0(\u_DECODE/n5 [0]),
    .i1(\u_BPU_BP/n2 [0]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [0]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b1  (
    .i0(bp_imm[1]),
    .i1(\u_BPU_BP/n2 [1]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [1]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b10  (
    .i0(bp_imm[10]),
    .i1(\u_BPU_BP/n2 [10]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [10]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b11  (
    .i0(bp_imm[11]),
    .i1(\u_BPU_BP/n2 [11]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [11]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b12  (
    .i0(bp_imm[12]),
    .i1(\u_BPU_BP/n2 [12]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [12]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b13  (
    .i0(bp_imm[13]),
    .i1(\u_BPU_BP/n2 [13]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [13]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b14  (
    .i0(bp_imm[14]),
    .i1(\u_BPU_BP/n2 [14]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [14]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b15  (
    .i0(bp_imm[15]),
    .i1(\u_BPU_BP/n2 [15]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [15]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b16  (
    .i0(bp_imm[16]),
    .i1(\u_BPU_BP/n2 [16]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [16]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b17  (
    .i0(bp_imm[17]),
    .i1(\u_BPU_BP/n2 [17]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [17]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b18  (
    .i0(bp_imm[18]),
    .i1(\u_BPU_BP/n2 [18]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [18]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b19  (
    .i0(bp_imm[19]),
    .i1(\u_BPU_BP/n2 [19]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [19]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b2  (
    .i0(bp_imm[2]),
    .i1(\u_BPU_BP/n2 [2]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [2]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b20  (
    .i0(bp_imm[31]),
    .i1(\u_BPU_BP/n2 [20]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [20]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b21  (
    .i0(bp_imm[31]),
    .i1(\u_BPU_BP/n2 [21]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [21]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b22  (
    .i0(bp_imm[31]),
    .i1(\u_BPU_BP/n2 [22]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [22]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b23  (
    .i0(bp_imm[31]),
    .i1(\u_BPU_BP/n2 [23]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [23]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b24  (
    .i0(bp_imm[31]),
    .i1(\u_BPU_BP/n2 [24]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [24]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b25  (
    .i0(bp_imm[31]),
    .i1(\u_BPU_BP/n2 [25]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [25]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b26  (
    .i0(bp_imm[31]),
    .i1(\u_BPU_BP/n2 [26]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [26]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b27  (
    .i0(bp_imm[31]),
    .i1(\u_BPU_BP/n2 [27]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [27]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b28  (
    .i0(bp_imm[31]),
    .i1(\u_BPU_BP/n2 [28]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [28]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b29  (
    .i0(bp_imm[31]),
    .i1(\u_BPU_BP/n2 [29]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [29]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b3  (
    .i0(bp_imm[3]),
    .i1(\u_BPU_BP/n2 [3]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [3]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b30  (
    .i0(bp_imm[31]),
    .i1(\u_BPU_BP/n2 [30]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [30]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b31  (
    .i0(bp_imm[31]),
    .i1(\u_BPU_BP/n2 [31]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [31]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b4  (
    .i0(bp_imm[4]),
    .i1(\u_BPU_BP/n2 [4]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [4]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b5  (
    .i0(bp_imm[5]),
    .i1(\u_BPU_BP/n2 [5]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [5]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b6  (
    .i0(bp_imm[6]),
    .i1(\u_BPU_BP/n2 [6]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [6]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b7  (
    .i0(bp_imm[7]),
    .i1(\u_BPU_BP/n2 [7]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [7]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b8  (
    .i0(bp_imm[8]),
    .i1(\u_BPU_BP/n2 [8]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [8]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux0_b9  (
    .i0(bp_imm[9]),
    .i1(\u_BPU_BP/n2 [9]),
    .sel(jalr_rs1ren),
    .o(\u_BPU_BP/n3 [9]));  // ../RTL/core/bpu_bp.v(44)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b0  (
    .i0(\u_BPU_BP/n4 [0]),
    .i1(\u_BPU_BP/n3 [0]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[0]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b1  (
    .i0(\u_BPU_BP/n4 [1]),
    .i1(\u_BPU_BP/n3 [1]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[1]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b10  (
    .i0(\u_BPU_BP/n4 [10]),
    .i1(\u_BPU_BP/n3 [10]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[10]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b11  (
    .i0(\u_BPU_BP/n4 [11]),
    .i1(\u_BPU_BP/n3 [11]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[11]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b12  (
    .i0(\u_BPU_BP/n4 [12]),
    .i1(\u_BPU_BP/n3 [12]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[12]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b13  (
    .i0(\u_BPU_BP/n4 [13]),
    .i1(\u_BPU_BP/n3 [13]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[13]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b14  (
    .i0(\u_BPU_BP/n4 [14]),
    .i1(\u_BPU_BP/n3 [14]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[14]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b15  (
    .i0(\u_BPU_BP/n4 [15]),
    .i1(\u_BPU_BP/n3 [15]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[15]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b16  (
    .i0(\u_BPU_BP/n4 [16]),
    .i1(\u_BPU_BP/n3 [16]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[16]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b17  (
    .i0(\u_BPU_BP/n4 [17]),
    .i1(\u_BPU_BP/n3 [17]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[17]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b18  (
    .i0(\u_BPU_BP/n4 [18]),
    .i1(\u_BPU_BP/n3 [18]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[18]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b19  (
    .i0(\u_BPU_BP/n4 [19]),
    .i1(\u_BPU_BP/n3 [19]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[19]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b2  (
    .i0(\u_BPU_BP/n4 [2]),
    .i1(\u_BPU_BP/n3 [2]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[2]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b20  (
    .i0(\u_BPU_BP/n4 [20]),
    .i1(\u_BPU_BP/n3 [20]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[20]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b21  (
    .i0(\u_BPU_BP/n4 [21]),
    .i1(\u_BPU_BP/n3 [21]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[21]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b22  (
    .i0(\u_BPU_BP/n4 [22]),
    .i1(\u_BPU_BP/n3 [22]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[22]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b23  (
    .i0(\u_BPU_BP/n4 [23]),
    .i1(\u_BPU_BP/n3 [23]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[23]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b24  (
    .i0(\u_BPU_BP/n4 [24]),
    .i1(\u_BPU_BP/n3 [24]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[24]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b25  (
    .i0(\u_BPU_BP/n4 [25]),
    .i1(\u_BPU_BP/n3 [25]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[25]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b26  (
    .i0(\u_BPU_BP/n4 [26]),
    .i1(\u_BPU_BP/n3 [26]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[26]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b27  (
    .i0(\u_BPU_BP/n4 [27]),
    .i1(\u_BPU_BP/n3 [27]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[27]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b28  (
    .i0(\u_BPU_BP/n4 [28]),
    .i1(\u_BPU_BP/n3 [28]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[28]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b29  (
    .i0(\u_BPU_BP/n4 [29]),
    .i1(\u_BPU_BP/n3 [29]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[29]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b3  (
    .i0(\u_BPU_BP/n4 [3]),
    .i1(\u_BPU_BP/n3 [3]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[3]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b30  (
    .i0(\u_BPU_BP/n4 [30]),
    .i1(\u_BPU_BP/n3 [30]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[30]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b31  (
    .i0(\u_BPU_BP/n4 [31]),
    .i1(\u_BPU_BP/n3 [31]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[31]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b4  (
    .i0(\u_BPU_BP/n4 [4]),
    .i1(\u_BPU_BP/n3 [4]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[4]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b5  (
    .i0(\u_BPU_BP/n4 [5]),
    .i1(\u_BPU_BP/n3 [5]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[5]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b6  (
    .i0(\u_BPU_BP/n4 [6]),
    .i1(\u_BPU_BP/n3 [6]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[6]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b7  (
    .i0(\u_BPU_BP/n4 [7]),
    .i1(\u_BPU_BP/n3 [7]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[7]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b8  (
    .i0(\u_BPU_BP/n4 [8]),
    .i1(\u_BPU_BP/n3 [8]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[8]));  // ../RTL/core/bpu_bp.v(43)
  binary_mux_s1_w1 \u_BPU_BP/mux1_b9  (
    .i0(\u_BPU_BP/n4 [9]),
    .i1(\u_BPU_BP/n3 [9]),
    .sel(inst_jalr),
    .o(o_bpu_jaddr[9]));  // ../RTL/core/bpu_bp.v(43)
  or \u_BPU_BP/u1  (\u_BPU_BP/n0 , inst_jalr, inst_jal);  // ../RTL/core/bpu_bp.v(40)
  and \u_BPU_BP/u2  (\u_BPU_BP/n1 , inst_bxx, bp_imm[31]);  // ../RTL/core/bpu_bp.v(40)
  or \u_BPU_BP/u3  (o_bpu_taken, \u_BPU_BP/n0 , \u_BPU_BP/n1 );  // ../RTL/core/bpu_bp.v(40)
  eq_w5 \u_DECODE/eq0  (
    .i0(i_data[6:2]),
    .i1(5'b11011),
    .o(\u_DECODE/n1 ));  // ../RTL/core/decode.v(55)
  eq_w5 \u_DECODE/eq1  (
    .i0(i_data[6:2]),
    .i1(5'b11001),
    .o(\u_DECODE/n2 ));  // ../RTL/core/decode.v(56)
  eq_w5 \u_DECODE/eq10  (
    .i0(i_data[6:2]),
    .i1(5'b00100),
    .o(\u_DECODE/opc_opimm ));  // ../RTL/core/decode.v(91)
  eq_w5 \u_DECODE/eq11  (
    .i0(i_data[6:2]),
    .i1(5'b01100),
    .o(\u_DECODE/opc_op ));  // ../RTL/core/decode.v(92)
  eq_w5 \u_DECODE/eq13  (
    .i0(i_data[6:2]),
    .i1(5'b11100),
    .o(o_decinfo_grp[4]));  // ../RTL/core/decode.v(94)
  eq_w3 \u_DECODE/eq14  (
    .i0(i_data[14:12]),
    .i1(3'b000),
    .o(\u_DECODE/func_000 ));  // ../RTL/core/decode.v(97)
  eq_w3 \u_DECODE/eq15  (
    .i0(i_data[14:12]),
    .i1(3'b001),
    .o(\u_DECODE/func_001 ));  // ../RTL/core/decode.v(98)
  eq_w3 \u_DECODE/eq16  (
    .i0(i_data[14:12]),
    .i1(3'b010),
    .o(\u_DECODE/func_010 ));  // ../RTL/core/decode.v(99)
  eq_w3 \u_DECODE/eq17  (
    .i0(i_data[14:12]),
    .i1(3'b011),
    .o(\u_DECODE/func_011 ));  // ../RTL/core/decode.v(100)
  eq_w3 \u_DECODE/eq18  (
    .i0(i_data[14:12]),
    .i1(3'b100),
    .o(\u_DECODE/func_100 ));  // ../RTL/core/decode.v(101)
  eq_w3 \u_DECODE/eq19  (
    .i0(i_data[14:12]),
    .i1(3'b101),
    .o(\u_DECODE/func_101 ));  // ../RTL/core/decode.v(102)
  eq_w5 \u_DECODE/eq2  (
    .i0(i_data[6:2]),
    .i1(5'b11000),
    .o(\u_DECODE/n3 ));  // ../RTL/core/decode.v(57)
  eq_w3 \u_DECODE/eq20  (
    .i0(i_data[14:12]),
    .i1(3'b110),
    .o(\u_DECODE/func_110 ));  // ../RTL/core/decode.v(103)
  eq_w3 \u_DECODE/eq21  (
    .i0(i_data[14:12]),
    .i1(3'b111),
    .o(\u_DECODE/func_111 ));  // ../RTL/core/decode.v(104)
  eq_w7 \u_DECODE/eq22  (
    .i0(i_data[31:25]),
    .i1(7'b0000000),
    .o(\u_DECODE/func7_0000000 ));  // ../RTL/core/decode.v(107)
  eq_w7 \u_DECODE/eq23  (
    .i0(i_data[31:25]),
    .i1(7'b0100000),
    .o(\u_DECODE/func7_0100000 ));  // ../RTL/core/decode.v(108)
  eq_w7 \u_DECODE/eq24  (
    .i0(i_data[31:25]),
    .i1(7'b0000001),
    .o(\u_DECODE/func7_0000001 ));  // ../RTL/core/decode.v(109)
  eq_w12 \u_DECODE/eq25  (
    .i0(i_data[31:20]),
    .i1(12'b000000000000),
    .o(\u_DECODE/type_i_imm_000000000000 ));  // ../RTL/core/decode.v(112)
  eq_w12 \u_DECODE/eq26  (
    .i0(i_data[31:20]),
    .i1(12'b000000000001),
    .o(\u_DECODE/type_i_imm_000000000001 ));  // ../RTL/core/decode.v(113)
  eq_w5 \u_DECODE/eq3  (
    .i0(i_data[6:2]),
    .i1(5'b01101),
    .o(\u_DECODE/opc_lui ));  // ../RTL/core/decode.v(84)
  eq_w5 \u_DECODE/eq4  (
    .i0(i_data[6:2]),
    .i1(5'b00101),
    .o(rs1topc));  // ../RTL/core/decode.v(85)
  eq_w5 \u_DECODE/eq8  (
    .i0(i_data[6:2]),
    .i1(5'b00000),
    .o(\u_DECODE/opc_load ));  // ../RTL/core/decode.v(89)
  eq_w5 \u_DECODE/eq9  (
    .i0(i_data[6:2]),
    .i1(5'b01000),
    .o(\u_DECODE/opc_store ));  // ../RTL/core/decode.v(90)
  binary_mux_s1_w1 \u_DECODE/mux0_b10  (
    .i0(i_data[30]),
    .i1(1'b0),
    .sel(\u_DECODE/n20 ),
    .o(\u_DECODE/inst_opimm_imm [10]));  // ../RTL/core/decode.v(202)
  binary_mux_s1_w1 \u_DECODE/mux0_b11  (
    .i0(i_data[31]),
    .i1(1'b0),
    .sel(\u_DECODE/n20 ),
    .o(\u_DECODE/inst_opimm_imm [11]));  // ../RTL/core/decode.v(202)
  binary_mux_s1_w1 \u_DECODE/mux0_b5  (
    .i0(i_data[25]),
    .i1(1'b0),
    .sel(\u_DECODE/n20 ),
    .o(\u_DECODE/inst_opimm_imm [5]));  // ../RTL/core/decode.v(202)
  binary_mux_s1_w1 \u_DECODE/mux0_b6  (
    .i0(i_data[26]),
    .i1(1'b0),
    .sel(\u_DECODE/n20 ),
    .o(\u_DECODE/inst_opimm_imm [6]));  // ../RTL/core/decode.v(202)
  binary_mux_s1_w1 \u_DECODE/mux0_b7  (
    .i0(i_data[27]),
    .i1(1'b0),
    .sel(\u_DECODE/n20 ),
    .o(\u_DECODE/inst_opimm_imm [7]));  // ../RTL/core/decode.v(202)
  binary_mux_s1_w1 \u_DECODE/mux0_b8  (
    .i0(i_data[28]),
    .i1(1'b0),
    .sel(\u_DECODE/n20 ),
    .o(\u_DECODE/inst_opimm_imm [8]));  // ../RTL/core/decode.v(202)
  binary_mux_s1_w1 \u_DECODE/mux0_b9  (
    .i0(i_data[29]),
    .i1(1'b0),
    .sel(\u_DECODE/n20 ),
    .o(\u_DECODE/inst_opimm_imm [9]));  // ../RTL/core/decode.v(202)
  ne_w5 \u_DECODE/neq0  (
    .i0(i_data[11:7]),
    .i1(5'b00000),
    .o(\u_DECODE/n30 ));  // ../RTL/core/decode.v(216)
  ne_w5 \u_DECODE/neq2  (
    .i0(i_data[24:20]),
    .i1(5'b00000),
    .o(\u_DECODE/n46 ));  // ../RTL/core/decode.v(241)
  or \u_DECODE/u100  (\u_DECODE/n6 [11], \u_DECODE/n4 [11], \u_DECODE/n5 [31]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u1000  (\u_DECODE/n22 [15], \u_DECODE/n21 , i_data[15]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1001  (\u_DECODE/n22 [16], \u_DECODE/n21 , i_data[16]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1002  (\u_DECODE/n22 [17], \u_DECODE/n21 , i_data[17]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1003  (\u_DECODE/n22 [18], \u_DECODE/n21 , i_data[18]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1004  (\u_DECODE/n22 [19], \u_DECODE/n21 , i_data[19]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1005  (\u_DECODE/n22 [20], \u_DECODE/n21 , i_data[20]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1006  (\u_DECODE/n22 [21], \u_DECODE/n21 , i_data[21]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1007  (\u_DECODE/n22 [22], \u_DECODE/n21 , i_data[22]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1008  (\u_DECODE/n22 [23], \u_DECODE/n21 , i_data[23]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1009  (\u_DECODE/n22 [24], \u_DECODE/n21 , i_data[24]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u101  (\u_DECODE/inst_divu , \u_DECODE/n15 , \u_DECODE/func7_0000001 );  // ../RTL/core/decode.v(179)
  and \u_DECODE/u1010  (\u_DECODE/n22 [25], \u_DECODE/n21 , i_data[25]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1011  (\u_DECODE/n22 [26], \u_DECODE/n21 , i_data[26]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1012  (\u_DECODE/n22 [27], \u_DECODE/n21 , i_data[27]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1013  (\u_DECODE/n22 [28], \u_DECODE/n21 , i_data[28]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1014  (\u_DECODE/n22 [29], \u_DECODE/n21 , i_data[29]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1015  (\u_DECODE/n22 [30], \u_DECODE/n21 , i_data[30]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u1016  (\u_DECODE/n22 [31], \u_DECODE/n21 , i_data[31]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u102  (\u_DECODE/n6 [10], \u_DECODE/n4 [10], \u_DECODE/n5 [10]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u1021  (\u_DECODE/n7 [1], inst_bxx, i_data[8]);  // ../RTL/core/decode.v(64)
  and \u_DECODE/u1022  (\u_DECODE/n7 [2], inst_bxx, i_data[9]);  // ../RTL/core/decode.v(64)
  and \u_DECODE/u1023  (\u_DECODE/n7 [3], inst_bxx, i_data[10]);  // ../RTL/core/decode.v(64)
  and \u_DECODE/u1024  (\u_DECODE/n7 [4], inst_bxx, i_data[11]);  // ../RTL/core/decode.v(64)
  and \u_DECODE/u1025  (\u_DECODE/n7 [5], inst_bxx, i_data[25]);  // ../RTL/core/decode.v(64)
  and \u_DECODE/u1026  (\u_DECODE/n7 [6], inst_bxx, i_data[26]);  // ../RTL/core/decode.v(64)
  and \u_DECODE/u1027  (\u_DECODE/n7 [7], inst_bxx, i_data[27]);  // ../RTL/core/decode.v(64)
  and \u_DECODE/u1028  (\u_DECODE/n7 [8], inst_bxx, i_data[28]);  // ../RTL/core/decode.v(64)
  and \u_DECODE/u1029  (\u_DECODE/n7 [9], inst_bxx, i_data[29]);  // ../RTL/core/decode.v(64)
  and \u_DECODE/u103  (\u_DECODE/inst_rem , \u_DECODE/n16 , \u_DECODE/func7_0000001 );  // ../RTL/core/decode.v(180)
  and \u_DECODE/u1030  (\u_DECODE/n7 [10], inst_bxx, i_data[30]);  // ../RTL/core/decode.v(64)
  and \u_DECODE/u1031  (\u_DECODE/n7 [11], inst_bxx, i_data[7]);  // ../RTL/core/decode.v(64)
  and \u_DECODE/u1032  (\u_DECODE/n7 [31], inst_bxx, i_data[31]);  // ../RTL/core/decode.v(64)
  or \u_DECODE/u104  (\u_DECODE/n6 [9], \u_DECODE/n4 [9], \u_DECODE/n5 [9]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u105  (\u_DECODE/inst_remu , \u_DECODE/n17 , \u_DECODE/func7_0000001 );  // ../RTL/core/decode.v(181)
  and \u_DECODE/u106  (o_decinfo_grp[3], \u_DECODE/opc_op , \u_DECODE/func7_0000001 );  // ../RTL/core/decode.v(183)
  or \u_DECODE/u11  (\u_DECODE/n69 [3], \u_DECODE/n67 [3], \u_DECODE/n68 [3]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u114  (\u_DECODE/n19 , \u_DECODE/inst_slli , \u_DECODE/inst_srli );  // ../RTL/core/decode.v(202)
  or \u_DECODE/u115  (\u_DECODE/n20 , \u_DECODE/n19 , \u_DECODE/inst_srai );  // ../RTL/core/decode.v(202)
  or \u_DECODE/u116  (\u_DECODE/n21 , \u_DECODE/opc_lui , rs1topc);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u118  (\u_DECODE/n69 [2], \u_DECODE/n67 [2], \u_DECODE/n68 [2]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u12  (o_decinfo[3], \u_DECODE/n71 [3], \u_DECODE/n72 [3]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u121  (\u_DECODE/n25 [0], \u_DECODE/opc_store , i_data[7]);  // ../RTL/core/decode.v(208)
  and \u_DECODE/u123  (\u_DECODE/n27 [0], \u_DECODE/opc_load , i_data[20]);  // ../RTL/core/decode.v(209)
  or \u_DECODE/u124  (\u_DECODE/n28 [0], \u_DECODE/n25 [0], \u_DECODE/n27 [0]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u125  (\u_DECODE/n29 [0], \u_DECODE/opc_opimm , i_data[20]);  // ../RTL/core/decode.v(210)
  or \u_DECODE/u126  (\u_DECODE/n6 [8], \u_DECODE/n4 [8], \u_DECODE/n5 [8]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u127  (\u_DECODE/n31 , \u_DECODE/n21 , \u_DECODE/n1 );  // ../RTL/core/decode.v(217)
  or \u_DECODE/u128  (\u_DECODE/n32 , \u_DECODE/n31 , \u_DECODE/n2 );  // ../RTL/core/decode.v(217)
  or \u_DECODE/u129  (\u_DECODE/n33 , \u_DECODE/n32 , \u_DECODE/opc_opimm );  // ../RTL/core/decode.v(217)
  or \u_DECODE/u130  (\u_DECODE/n34 , \u_DECODE/n33 , \u_DECODE/opc_op );  // ../RTL/core/decode.v(217)
  or \u_DECODE/u131  (\u_DECODE/n35 , \u_DECODE/n34 , o_decinfo_grp[4]);  // ../RTL/core/decode.v(217)
  or \u_DECODE/u132  (\u_DECODE/n36 , \u_DECODE/n35 , \u_DECODE/opc_load );  // ../RTL/core/decode.v(217)
  and \u_DECODE/u133  (o_rdwen, \u_DECODE/n30 , \u_DECODE/n36 );  // ../RTL/core/decode.v(216)
  or \u_DECODE/u134  (o_imm[0], \u_DECODE/n28 [0], \u_DECODE/n29 [0]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u135  (\u_DECODE/n38 , \u_DECODE/n2 , \u_DECODE/n3 );  // ../RTL/core/decode.v(229)
  or \u_DECODE/u136  (\u_DECODE/n39 , \u_DECODE/n38 , \u_DECODE/opc_load );  // ../RTL/core/decode.v(229)
  or \u_DECODE/u137  (\u_DECODE/n40 , \u_DECODE/n39 , \u_DECODE/opc_store );  // ../RTL/core/decode.v(229)
  or \u_DECODE/u138  (\u_DECODE/n41 , \u_DECODE/n40 , \u_DECODE/opc_opimm );  // ../RTL/core/decode.v(229)
  or \u_DECODE/u139  (\u_DECODE/n42 , \u_DECODE/n41 , \u_DECODE/opc_op );  // ../RTL/core/decode.v(229)
  and \u_DECODE/u14  (\u_DECODE/opc_rv32 , i_data[1], i_data[0]);  // ../RTL/core/decode.v(67)
  or \u_DECODE/u140  (\u_DECODE/n43 , \u_DECODE/n42 , \u_DECODE/inst_csrrw );  // ../RTL/core/decode.v(229)
  or \u_DECODE/u141  (\u_DECODE/n44 , \u_DECODE/n43 , \u_DECODE/inst_csrrs );  // ../RTL/core/decode.v(229)
  or \u_DECODE/u142  (\u_DECODE/n45 , \u_DECODE/n44 , \u_DECODE/inst_csrrc );  // ../RTL/core/decode.v(229)
  and \u_DECODE/u143  (rs1ren, n1, \u_DECODE/n45 );  // ../RTL/core/decode.v(228)
  or \u_DECODE/u145  (\u_DECODE/n47 , \u_DECODE/n3 , \u_DECODE/opc_store );  // ../RTL/core/decode.v(242)
  or \u_DECODE/u146  (\u_DECODE/n48 , \u_DECODE/n47 , \u_DECODE/opc_op );  // ../RTL/core/decode.v(242)
  and \u_DECODE/u147  (rs2ren, \u_DECODE/n46 , \u_DECODE/n48 );  // ../RTL/core/decode.v(241)
  or \u_DECODE/u149  (\u_DECODE/n6 [7], \u_DECODE/n4 [7], \u_DECODE/n5 [7]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u150  (\u_DECODE/n49 , \u_DECODE/n21 , \u_DECODE/opc_opimm );  // ../RTL/core/decode.v(253)
  not \u_DECODE/u151  (\u_DECODE/n50 , o_decinfo_grp[3]);  // ../RTL/core/decode.v(253)
  and \u_DECODE/u152  (\u_DECODE/n51 , \u_DECODE/opc_op , \u_DECODE/n50 );  // ../RTL/core/decode.v(253)
  and \u_DECODE/u154  (\u_DECODE/n70 [8], o_decinfo_grp[3], \u_DECODE/inst_remu );  // ../RTL/core/decode.v(340)
  or \u_DECODE/u155  (\u_DECODE/bjuinfo [1], \u_DECODE/n1 , \u_DECODE/n2 );  // ../RTL/core/decode.v(255)
  and \u_DECODE/u156  (\u_DECODE/n70 [7], o_decinfo_grp[3], \u_DECODE/inst_rem );  // ../RTL/core/decode.v(340)
  and \u_DECODE/u157  (\u_DECODE/n70 [6], o_decinfo_grp[3], \u_DECODE/inst_divu );  // ../RTL/core/decode.v(340)
  or \u_DECODE/u159  (\u_DECODE/n6 [6], \u_DECODE/n4 [6], \u_DECODE/n5 [6]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u160  (\u_DECODE/n52 , \u_DECODE/n21 , \u_DECODE/inst_add );  // ../RTL/core/decode.v(258)
  or \u_DECODE/u161  (\u_DECODE/n53 , \u_DECODE/n52 , \u_DECODE/inst_addi );  // ../RTL/core/decode.v(258)
  or \u_DECODE/u162  (\u_DECODE/n54 , \u_DECODE/n53 , \u_DECODE/opc_load );  // ../RTL/core/decode.v(258)
  or \u_DECODE/u163  (\u_DECODE/aluinfo [2], \u_DECODE/inst_sll , \u_DECODE/inst_slli );  // ../RTL/core/decode.v(270)
  and \u_DECODE/u165  (\u_DECODE/n70 [5], o_decinfo_grp[3], \u_DECODE/inst_div );  // ../RTL/core/decode.v(340)
  and \u_DECODE/u166  (\u_DECODE/n70 [4], o_decinfo_grp[3], \u_DECODE/inst_mulhu );  // ../RTL/core/decode.v(340)
  and \u_DECODE/u167  (\u_DECODE/n70 [3], o_decinfo_grp[3], \u_DECODE/inst_mulhsu );  // ../RTL/core/decode.v(340)
  and \u_DECODE/u168  (\u_DECODE/n70 [2], o_decinfo_grp[3], \u_DECODE/inst_mulh );  // ../RTL/core/decode.v(340)
  and \u_DECODE/u169  (\u_DECODE/n70 [1], o_decinfo_grp[3], \u_DECODE/inst_mul );  // ../RTL/core/decode.v(340)
  or \u_DECODE/u171  (\u_DECODE/n71 [8], \u_DECODE/n69 [8], \u_DECODE/n70 [8]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u174  (\u_DECODE/n6 [5], \u_DECODE/n4 [5], \u_DECODE/n5 [5]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u175  (\u_DECODE/n6 [4], \u_DECODE/n4 [4], \u_DECODE/n5 [4]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u176  (\u_DECODE/n55 , \u_DECODE/n49 , \u_DECODE/opc_load );  // ../RTL/core/decode.v(275)
  or \u_DECODE/u177  (rs2toimm, \u_DECODE/n55 , \u_DECODE/opc_store );  // ../RTL/core/decode.v(275)
  or \u_DECODE/u178  (\u_DECODE/n71 [5], \u_DECODE/n69 [5], \u_DECODE/n70 [5]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u179  (\u_DECODE/n71 [7], \u_DECODE/n69 [7], \u_DECODE/n70 [7]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u180  (\u_DECODE/n71 [6], \u_DECODE/n69 [6], \u_DECODE/n70 [6]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u181  (\u_DECODE/lsuinfo [2], \u_DECODE/func_000 , \u_DECODE/func_100 );  // ../RTL/core/decode.v(284)
  or \u_DECODE/u183  (\u_DECODE/n6 [3], \u_DECODE/n4 [3], \u_DECODE/n5 [3]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u184  (\u_DECODE/n71 [4], \u_DECODE/n69 [4], \u_DECODE/n70 [4]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u185  (\u_DECODE/n71 [3], \u_DECODE/n69 [3], \u_DECODE/n70 [3]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u186  (\u_DECODE/n71 [2], \u_DECODE/n69 [2], \u_DECODE/n70 [2]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u187  (\u_DECODE/n71 [1], \u_DECODE/n69 [1], \u_DECODE/n70 [1]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u191  (\u_DECODE/n72 [7], o_decinfo_grp[4], \u_DECODE/scuinfo [7]);  // ../RTL/core/decode.v(341)
  and \u_DECODE/u192  (\u_DECODE/n72 [6], o_decinfo_grp[4], i_data[14]);  // ../RTL/core/decode.v(341)
  and \u_DECODE/u193  (\u_DECODE/n72 [5], o_decinfo_grp[4], \u_DECODE/scuinfo [5]);  // ../RTL/core/decode.v(341)
  and \u_DECODE/u194  (\u_DECODE/n72 [4], o_decinfo_grp[4], \u_DECODE/n61 );  // ../RTL/core/decode.v(341)
  and \u_DECODE/u195  (\u_DECODE/n72 [3], o_decinfo_grp[4], \u_DECODE/scuinfo [3]);  // ../RTL/core/decode.v(341)
  and \u_DECODE/u196  (\u_DECODE/n72 [2], o_decinfo_grp[4], \u_DECODE/inst_ebreak );  // ../RTL/core/decode.v(341)
  and \u_DECODE/u197  (\u_DECODE/n72 [1], o_decinfo_grp[4], \u_DECODE/inst_ecall );  // ../RTL/core/decode.v(341)
  or \u_DECODE/u2  (o_decinfo[4], \u_DECODE/n71 [4], \u_DECODE/n72 [4]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u200  (\u_DECODE/n64 , i_data[13], i_data[14]);  // ../RTL/core/decode.v(313)
  and \u_DECODE/u201  (\u_DECODE/n58 , \u_DECODE/inst_csrrw , \u_DECODE/inst_csrrwi );  // ../RTL/core/decode.v(313)
  or \u_DECODE/u202  (\u_DECODE/n6 [2], \u_DECODE/n4 [2], \u_DECODE/n5 [2]);  // ../RTL/core/decode.v(62)
  AL_MUX \u_DECODE/u203  (
    .i0(1'b1),
    .i1(\u_DECODE/n30 ),
    .sel(\u_DECODE/n58 ),
    .o(\u_DECODE/n59 ));  // ../RTL/core/decode.v(313)
  and \u_DECODE/u204  (o_csr_ren, \u_DECODE/n57 [0], \u_DECODE/n59 );  // ../RTL/core/decode.v(313)
  and \u_DECODE/u205  (\u_DECODE/n5 [0], inst_jalr, i_data[20]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u206  (\u_DECODE/n60 , o_csr_ren, i_data[14]);  // ../RTL/core/decode.v(317)
  and \u_DECODE/u207  (o_csridx[0], o_csr_ren, i_data[20]);  // ../RTL/core/decode.v(315)
  or \u_DECODE/u210  (o_decinfo[7], \u_DECODE/n71 [7], \u_DECODE/n72 [7]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u211  (o_decinfo[6], \u_DECODE/n71 [6], \u_DECODE/n72 [6]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u212  (o_decinfo[5], \u_DECODE/n71 [5], \u_DECODE/n72 [5]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u213  (o_csr_zimm[0], \u_DECODE/n60 , i_data[15]);  // ../RTL/core/decode.v(317)
  or \u_DECODE/u214  (\u_DECODE/n61 , \u_DECODE/inst_csrrs , \u_DECODE/inst_csrrsi );  // ../RTL/core/decode.v(330)
  or \u_DECODE/u215  (\u_DECODE/n62 , \u_DECODE/n61 , \u_DECODE/inst_csrrc );  // ../RTL/core/decode.v(330)
  or \u_DECODE/u216  (\u_DECODE/n63 , \u_DECODE/n62 , \u_DECODE/inst_csrrci );  // ../RTL/core/decode.v(330)
  or \u_DECODE/u217  (\u_DECODE/n6 [1], \u_DECODE/n4 [1], \u_DECODE/n5 [1]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u218  (\u_DECODE/scuinfo [3], \u_DECODE/inst_csrrw , \u_DECODE/inst_csrrwi );  // ../RTL/core/decode.v(325)
  AL_MUX \u_DECODE/u219  (
    .i0(\u_DECODE/n56 ),
    .i1(n1),
    .sel(\u_DECODE/n63 ),
    .o(\u_DECODE/scuinfo [7]));  // ../RTL/core/decode.v(330)
  and \u_DECODE/u220  (\u_DECODE/n57 [0], o_decinfo_grp[4], \u_DECODE/n56 );  // ../RTL/core/decode.v(313)
  or \u_DECODE/u222  (\u_DECODE/n69 [1], \u_DECODE/n67 [1], \u_DECODE/n68 [1]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u223  (o_decinfo_grp[0], \u_DECODE/n49 , \u_DECODE/n51 );  // ../RTL/core/decode.v(258)
  or \u_DECODE/u231  (\u_DECODE/n69 [4], \u_DECODE/n67 [4], \u_DECODE/n68 [4]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u232  (\u_DECODE/n69 [5], \u_DECODE/n67 [5], \u_DECODE/n68 [5]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u233  (\u_DECODE/n69 [6], \u_DECODE/n65 [6], \u_DECODE/n68 [6]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u234  (\u_DECODE/n69 [7], \u_DECODE/n65 [7], \u_DECODE/n68 [7]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u235  (\u_DECODE/n69 [8], \u_DECODE/n65 [8], \u_DECODE/n68 [8]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u237  (\u_DECODE/n68 [1], o_decinfo_grp[2], \u_DECODE/bjuinfo [1]);  // ../RTL/core/decode.v(339)
  and \u_DECODE/u238  (\u_DECODE/n68 [2], o_decinfo_grp[2], \u_DECODE/inst_beq );  // ../RTL/core/decode.v(339)
  and \u_DECODE/u239  (\u_DECODE/n68 [3], o_decinfo_grp[2], \u_DECODE/inst_bne );  // ../RTL/core/decode.v(339)
  and \u_DECODE/u240  (\u_DECODE/n68 [4], o_decinfo_grp[2], \u_DECODE/inst_blt );  // ../RTL/core/decode.v(339)
  and \u_DECODE/u241  (\u_DECODE/n68 [5], o_decinfo_grp[2], \u_DECODE/inst_bge );  // ../RTL/core/decode.v(339)
  and \u_DECODE/u242  (\u_DECODE/n68 [6], o_decinfo_grp[2], \u_DECODE/inst_bltu );  // ../RTL/core/decode.v(339)
  and \u_DECODE/u243  (\u_DECODE/n68 [7], o_decinfo_grp[2], \u_DECODE/inst_bgeu );  // ../RTL/core/decode.v(339)
  and \u_DECODE/u244  (\u_DECODE/n68 [8], o_decinfo_grp[2], bpu_bflag);  // ../RTL/core/decode.v(339)
  or \u_DECODE/u246  (\u_DECODE/n67 [1], \u_DECODE/n65 [1], \u_DECODE/n66 [1]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u247  (\u_DECODE/n67 [2], \u_DECODE/n65 [2], \u_DECODE/n66 [2]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u248  (\u_DECODE/n67 [3], \u_DECODE/n65 [3], \u_DECODE/n66 [3]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u249  (\u_DECODE/n67 [4], \u_DECODE/n65 [4], \u_DECODE/n66 [4]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u250  (\u_DECODE/n67 [5], \u_DECODE/n65 [5], \u_DECODE/n66 [5]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u255  (o_decinfo_grp[1], \u_DECODE/opc_load , \u_DECODE/opc_store );  // ../RTL/core/decode.v(258)
  or \u_DECODE/u256  (o_decinfo_grp[2], \u_DECODE/bjuinfo [1], \u_DECODE/n3 );  // ../RTL/core/decode.v(258)
  or \u_DECODE/u257  (o_decinfo_grp[5], \u_DECODE/n54 , \u_DECODE/opc_store );  // ../RTL/core/decode.v(258)
  or \u_DECODE/u264  (\u_DECODE/scuinfo [5], \u_DECODE/inst_csrrc , \u_DECODE/inst_csrrci );  // ../RTL/core/decode.v(325)
  and \u_DECODE/u265  (o_csr_zimm[1], \u_DECODE/n60 , i_data[16]);  // ../RTL/core/decode.v(317)
  and \u_DECODE/u266  (o_csr_zimm[2], \u_DECODE/n60 , i_data[17]);  // ../RTL/core/decode.v(317)
  and \u_DECODE/u267  (o_csr_zimm[3], \u_DECODE/n60 , i_data[18]);  // ../RTL/core/decode.v(317)
  and \u_DECODE/u268  (o_csr_zimm[4], \u_DECODE/n60 , i_data[19]);  // ../RTL/core/decode.v(317)
  and \u_DECODE/u296  (o_csridx[1], o_csr_ren, i_data[21]);  // ../RTL/core/decode.v(315)
  and \u_DECODE/u297  (o_csridx[2], o_csr_ren, i_data[22]);  // ../RTL/core/decode.v(315)
  and \u_DECODE/u298  (o_csridx[3], o_csr_ren, i_data[23]);  // ../RTL/core/decode.v(315)
  and \u_DECODE/u299  (o_csridx[4], o_csr_ren, i_data[24]);  // ../RTL/core/decode.v(315)
  and \u_DECODE/u300  (o_csridx[5], o_csr_ren, i_data[25]);  // ../RTL/core/decode.v(315)
  and \u_DECODE/u301  (o_csridx[6], o_csr_ren, i_data[26]);  // ../RTL/core/decode.v(315)
  and \u_DECODE/u302  (o_csridx[7], o_csr_ren, i_data[27]);  // ../RTL/core/decode.v(315)
  and \u_DECODE/u303  (o_csridx[8], o_csr_ren, i_data[28]);  // ../RTL/core/decode.v(315)
  and \u_DECODE/u304  (o_csridx[9], o_csr_ren, i_data[29]);  // ../RTL/core/decode.v(315)
  and \u_DECODE/u305  (o_csridx[10], o_csr_ren, i_data[30]);  // ../RTL/core/decode.v(315)
  and \u_DECODE/u306  (o_csridx[11], o_csr_ren, i_data[31]);  // ../RTL/core/decode.v(315)
  and \u_DECODE/u307  (\u_DECODE/n5 [1], inst_jalr, i_data[21]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u308  (\u_DECODE/n5 [2], inst_jalr, i_data[22]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u309  (\u_DECODE/n5 [3], inst_jalr, i_data[23]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u310  (\u_DECODE/n5 [4], inst_jalr, i_data[24]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u311  (\u_DECODE/n5 [5], inst_jalr, i_data[25]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u312  (\u_DECODE/n5 [6], inst_jalr, i_data[26]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u313  (\u_DECODE/n5 [7], inst_jalr, i_data[27]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u314  (\u_DECODE/n5 [8], inst_jalr, i_data[28]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u315  (\u_DECODE/n5 [9], inst_jalr, i_data[29]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u316  (\u_DECODE/n5 [10], inst_jalr, i_data[30]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u317  (\u_DECODE/n5 [31], inst_jalr, i_data[31]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u318  (\u_DECODE/n4 [1], inst_jal, i_data[21]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u319  (\u_DECODE/n4 [2], inst_jal, i_data[22]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u32  (\u_DECODE/inst_beq , \u_DECODE/n3 , \u_DECODE/func_000 );  // ../RTL/core/decode.v(123)
  and \u_DECODE/u320  (\u_DECODE/n4 [3], inst_jal, i_data[23]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u321  (\u_DECODE/n4 [4], inst_jal, i_data[24]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u322  (\u_DECODE/n4 [5], inst_jal, i_data[25]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u323  (\u_DECODE/n4 [6], inst_jal, i_data[26]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u324  (\u_DECODE/n4 [7], inst_jal, i_data[27]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u325  (\u_DECODE/n4 [8], inst_jal, i_data[28]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u326  (\u_DECODE/n4 [9], inst_jal, i_data[29]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u327  (\u_DECODE/n4 [10], inst_jal, i_data[30]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u328  (\u_DECODE/n4 [11], inst_jal, i_data[20]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u329  (\u_DECODE/n4 [12], inst_jal, i_data[12]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u33  (\u_DECODE/inst_bne , \u_DECODE/n3 , \u_DECODE/func_001 );  // ../RTL/core/decode.v(124)
  and \u_DECODE/u330  (\u_DECODE/n4 [13], inst_jal, i_data[13]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u331  (\u_DECODE/n4 [14], inst_jal, i_data[14]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u332  (\u_DECODE/n4 [15], inst_jal, i_data[15]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u333  (\u_DECODE/n4 [16], inst_jal, i_data[16]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u334  (\u_DECODE/n4 [17], inst_jal, i_data[17]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u335  (\u_DECODE/n4 [18], inst_jal, i_data[18]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u336  (\u_DECODE/n4 [19], inst_jal, i_data[19]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u337  (\u_DECODE/n4 [31], inst_jal, i_data[31]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u338  (\u_DECODE/n56 , i_data[12], \u_DECODE/n64 );  // ../RTL/core/decode.v(313)
  and \u_DECODE/u34  (\u_DECODE/inst_blt , \u_DECODE/n3 , \u_DECODE/func_100 );  // ../RTL/core/decode.v(125)
  and \u_DECODE/u35  (\u_DECODE/inst_bge , \u_DECODE/n3 , \u_DECODE/func_101 );  // ../RTL/core/decode.v(126)
  or \u_DECODE/u355  (\u_DECODE/lsuinfo [3], \u_DECODE/func_001 , \u_DECODE/func_101 );  // ../RTL/core/decode.v(284)
  or \u_DECODE/u356  (\u_DECODE/lsuinfo [5], \u_DECODE/func_100 , \u_DECODE/func_101 );  // ../RTL/core/decode.v(284)
  or \u_DECODE/u358  (\u_DECODE/aluinfo [3], \u_DECODE/inst_srl , \u_DECODE/inst_srli );  // ../RTL/core/decode.v(270)
  or \u_DECODE/u359  (\u_DECODE/aluinfo [4], \u_DECODE/inst_sra , \u_DECODE/inst_srai );  // ../RTL/core/decode.v(270)
  and \u_DECODE/u36  (\u_DECODE/inst_bltu , \u_DECODE/n3 , \u_DECODE/func_110 );  // ../RTL/core/decode.v(127)
  or \u_DECODE/u360  (\u_DECODE/aluinfo [5], \u_DECODE/inst_xor , \u_DECODE/inst_xori );  // ../RTL/core/decode.v(270)
  or \u_DECODE/u361  (\u_DECODE/aluinfo [6], \u_DECODE/inst_and , \u_DECODE/inst_andi );  // ../RTL/core/decode.v(270)
  or \u_DECODE/u362  (\u_DECODE/aluinfo [7], \u_DECODE/inst_or , \u_DECODE/inst_ori );  // ../RTL/core/decode.v(270)
  or \u_DECODE/u363  (\u_DECODE/aluinfo [8], \u_DECODE/inst_slt , \u_DECODE/inst_slti );  // ../RTL/core/decode.v(270)
  or \u_DECODE/u364  (\u_DECODE/aluinfo [9], \u_DECODE/inst_sltu , \u_DECODE/inst_sltiu );  // ../RTL/core/decode.v(270)
  and \u_DECODE/u37  (\u_DECODE/inst_bgeu , \u_DECODE/n3 , \u_DECODE/func_111 );  // ../RTL/core/decode.v(128)
  or \u_DECODE/u377  (o_imm[1], \u_DECODE/n28 [1], \u_DECODE/n29 [1]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u378  (o_imm[2], \u_DECODE/n28 [2], \u_DECODE/n29 [2]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u379  (o_imm[3], \u_DECODE/n28 [3], \u_DECODE/n29 [3]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u380  (o_imm[4], \u_DECODE/n28 [4], \u_DECODE/n29 [4]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u381  (o_imm[5], \u_DECODE/n28 [5], \u_DECODE/n29 [5]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u382  (o_imm[6], \u_DECODE/n28 [6], \u_DECODE/n29 [6]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u383  (o_imm[7], \u_DECODE/n28 [7], \u_DECODE/n29 [7]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u384  (o_imm[8], \u_DECODE/n28 [8], \u_DECODE/n29 [8]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u385  (o_imm[9], \u_DECODE/n28 [9], \u_DECODE/n29 [9]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u386  (o_imm[10], \u_DECODE/n28 [10], \u_DECODE/n29 [10]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u387  (o_imm[11], \u_DECODE/n28 [11], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u388  (o_imm[12], \u_DECODE/n28 [12], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u389  (o_imm[13], \u_DECODE/n28 [13], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u390  (o_imm[14], \u_DECODE/n28 [14], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u391  (o_imm[15], \u_DECODE/n28 [15], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u392  (o_imm[16], \u_DECODE/n28 [16], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u393  (o_imm[17], \u_DECODE/n28 [17], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u394  (o_imm[18], \u_DECODE/n28 [18], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u395  (o_imm[19], \u_DECODE/n28 [19], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u396  (o_imm[20], \u_DECODE/n28 [20], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u397  (o_imm[21], \u_DECODE/n28 [21], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u398  (o_imm[22], \u_DECODE/n28 [22], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u399  (o_imm[23], \u_DECODE/n28 [23], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u4  (\u_DECODE/n0 , \u_DECODE/opc_rv32 , i_data_vld);  // ../RTL/core/decode.v(55)
  or \u_DECODE/u400  (o_imm[24], \u_DECODE/n28 [24], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u401  (o_imm[25], \u_DECODE/n28 [25], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u402  (o_imm[26], \u_DECODE/n28 [26], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u403  (o_imm[27], \u_DECODE/n28 [27], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u404  (o_imm[28], \u_DECODE/n28 [28], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u405  (o_imm[29], \u_DECODE/n28 [29], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u406  (o_imm[30], \u_DECODE/n28 [30], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u407  (o_imm[31], \u_DECODE/n28 [31], \u_DECODE/n29 [11]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u408  (\u_DECODE/n29 [1], \u_DECODE/opc_opimm , i_data[21]);  // ../RTL/core/decode.v(210)
  and \u_DECODE/u409  (\u_DECODE/n29 [2], \u_DECODE/opc_opimm , i_data[22]);  // ../RTL/core/decode.v(210)
  and \u_DECODE/u410  (\u_DECODE/n29 [3], \u_DECODE/opc_opimm , i_data[23]);  // ../RTL/core/decode.v(210)
  and \u_DECODE/u411  (\u_DECODE/n29 [4], \u_DECODE/opc_opimm , i_data[24]);  // ../RTL/core/decode.v(210)
  and \u_DECODE/u412  (\u_DECODE/n29 [5], \u_DECODE/opc_opimm , \u_DECODE/inst_opimm_imm [5]);  // ../RTL/core/decode.v(210)
  and \u_DECODE/u413  (\u_DECODE/n29 [6], \u_DECODE/opc_opimm , \u_DECODE/inst_opimm_imm [6]);  // ../RTL/core/decode.v(210)
  and \u_DECODE/u414  (\u_DECODE/n29 [7], \u_DECODE/opc_opimm , \u_DECODE/inst_opimm_imm [7]);  // ../RTL/core/decode.v(210)
  and \u_DECODE/u415  (\u_DECODE/n29 [8], \u_DECODE/opc_opimm , \u_DECODE/inst_opimm_imm [8]);  // ../RTL/core/decode.v(210)
  and \u_DECODE/u416  (\u_DECODE/n29 [9], \u_DECODE/opc_opimm , \u_DECODE/inst_opimm_imm [9]);  // ../RTL/core/decode.v(210)
  and \u_DECODE/u417  (\u_DECODE/n29 [10], \u_DECODE/opc_opimm , \u_DECODE/inst_opimm_imm [10]);  // ../RTL/core/decode.v(210)
  and \u_DECODE/u418  (\u_DECODE/n29 [11], \u_DECODE/opc_opimm , \u_DECODE/inst_opimm_imm [11]);  // ../RTL/core/decode.v(210)
  or \u_DECODE/u439  (\u_DECODE/n28 [1], \u_DECODE/n26 [1], \u_DECODE/n27 [1]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u440  (\u_DECODE/n28 [2], \u_DECODE/n26 [2], \u_DECODE/n27 [2]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u441  (\u_DECODE/n28 [3], \u_DECODE/n26 [3], \u_DECODE/n27 [3]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u442  (\u_DECODE/n28 [4], \u_DECODE/n26 [4], \u_DECODE/n27 [4]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u443  (\u_DECODE/n28 [5], \u_DECODE/n26 [5], \u_DECODE/n27 [5]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u444  (\u_DECODE/n28 [6], \u_DECODE/n26 [6], \u_DECODE/n27 [6]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u445  (\u_DECODE/n28 [7], \u_DECODE/n26 [7], \u_DECODE/n27 [7]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u446  (\u_DECODE/n28 [8], \u_DECODE/n26 [8], \u_DECODE/n27 [8]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u447  (\u_DECODE/n28 [9], \u_DECODE/n26 [9], \u_DECODE/n27 [9]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u448  (\u_DECODE/n28 [10], \u_DECODE/n26 [10], \u_DECODE/n27 [10]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u449  (\u_DECODE/n28 [11], \u_DECODE/n26 [11], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u450  (\u_DECODE/n28 [12], \u_DECODE/n26 [12], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u451  (\u_DECODE/n28 [13], \u_DECODE/n26 [13], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u452  (\u_DECODE/n28 [14], \u_DECODE/n26 [14], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u453  (\u_DECODE/n28 [15], \u_DECODE/n26 [15], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u454  (\u_DECODE/n28 [16], \u_DECODE/n26 [16], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u455  (\u_DECODE/n28 [17], \u_DECODE/n26 [17], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u456  (\u_DECODE/n28 [18], \u_DECODE/n26 [18], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u457  (\u_DECODE/n28 [19], \u_DECODE/n26 [19], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u458  (\u_DECODE/n28 [20], \u_DECODE/n26 [20], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u459  (\u_DECODE/n28 [21], \u_DECODE/n26 [21], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u46  (\u_DECODE/inst_addi , \u_DECODE/opc_opimm , \u_DECODE/func_000 );  // ../RTL/core/decode.v(140)
  or \u_DECODE/u460  (\u_DECODE/n28 [22], \u_DECODE/n26 [22], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u461  (\u_DECODE/n28 [23], \u_DECODE/n26 [23], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u462  (\u_DECODE/n28 [24], \u_DECODE/n26 [24], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u463  (\u_DECODE/n28 [25], \u_DECODE/n26 [25], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u464  (\u_DECODE/n28 [26], \u_DECODE/n26 [26], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u465  (\u_DECODE/n28 [27], \u_DECODE/n26 [27], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u466  (\u_DECODE/n28 [28], \u_DECODE/n26 [28], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u467  (\u_DECODE/n28 [29], \u_DECODE/n26 [29], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u468  (\u_DECODE/n28 [30], \u_DECODE/n26 [30], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u469  (\u_DECODE/n28 [31], \u_DECODE/n26 [31], \u_DECODE/n27 [11]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u47  (\u_DECODE/inst_slti , \u_DECODE/opc_opimm , \u_DECODE/func_010 );  // ../RTL/core/decode.v(141)
  and \u_DECODE/u470  (\u_DECODE/n27 [1], \u_DECODE/opc_load , i_data[21]);  // ../RTL/core/decode.v(209)
  and \u_DECODE/u471  (\u_DECODE/n27 [2], \u_DECODE/opc_load , i_data[22]);  // ../RTL/core/decode.v(209)
  and \u_DECODE/u472  (\u_DECODE/n27 [3], \u_DECODE/opc_load , i_data[23]);  // ../RTL/core/decode.v(209)
  and \u_DECODE/u473  (\u_DECODE/n27 [4], \u_DECODE/opc_load , i_data[24]);  // ../RTL/core/decode.v(209)
  and \u_DECODE/u474  (\u_DECODE/n27 [5], \u_DECODE/opc_load , i_data[25]);  // ../RTL/core/decode.v(209)
  and \u_DECODE/u475  (\u_DECODE/n27 [6], \u_DECODE/opc_load , i_data[26]);  // ../RTL/core/decode.v(209)
  and \u_DECODE/u476  (\u_DECODE/n27 [7], \u_DECODE/opc_load , i_data[27]);  // ../RTL/core/decode.v(209)
  and \u_DECODE/u477  (\u_DECODE/n27 [8], \u_DECODE/opc_load , i_data[28]);  // ../RTL/core/decode.v(209)
  and \u_DECODE/u478  (\u_DECODE/n27 [9], \u_DECODE/opc_load , i_data[29]);  // ../RTL/core/decode.v(209)
  and \u_DECODE/u479  (\u_DECODE/n27 [10], \u_DECODE/opc_load , i_data[30]);  // ../RTL/core/decode.v(209)
  and \u_DECODE/u48  (\u_DECODE/inst_sltiu , \u_DECODE/opc_opimm , \u_DECODE/func_011 );  // ../RTL/core/decode.v(142)
  and \u_DECODE/u480  (\u_DECODE/n27 [11], \u_DECODE/opc_load , i_data[31]);  // ../RTL/core/decode.v(209)
  and \u_DECODE/u49  (\u_DECODE/inst_xori , \u_DECODE/opc_opimm , \u_DECODE/func_100 );  // ../RTL/core/decode.v(143)
  AL_MUX \u_DECODE/u5  (
    .i0(1'b0),
    .i1(\u_DECODE/n1 ),
    .sel(\u_DECODE/n0 ),
    .o(inst_jal));  // ../RTL/core/decode.v(55)
  and \u_DECODE/u50  (\u_DECODE/inst_ori , \u_DECODE/opc_opimm , \u_DECODE/func_110 );  // ../RTL/core/decode.v(144)
  or \u_DECODE/u501  (\u_DECODE/n26 [1], \u_DECODE/n23 [1], \u_DECODE/n25 [1]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u502  (\u_DECODE/n26 [2], \u_DECODE/n23 [2], \u_DECODE/n25 [2]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u503  (\u_DECODE/n26 [3], \u_DECODE/n23 [3], \u_DECODE/n25 [3]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u504  (\u_DECODE/n26 [4], \u_DECODE/n23 [4], \u_DECODE/n25 [4]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u505  (\u_DECODE/n26 [5], \u_DECODE/n23 [5], \u_DECODE/n25 [5]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u506  (\u_DECODE/n26 [6], \u_DECODE/n23 [6], \u_DECODE/n25 [6]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u507  (\u_DECODE/n26 [7], \u_DECODE/n23 [7], \u_DECODE/n25 [7]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u508  (\u_DECODE/n26 [8], \u_DECODE/n23 [8], \u_DECODE/n25 [8]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u509  (\u_DECODE/n26 [9], \u_DECODE/n23 [9], \u_DECODE/n25 [9]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u51  (\u_DECODE/inst_andi , \u_DECODE/opc_opimm , \u_DECODE/func_111 );  // ../RTL/core/decode.v(145)
  or \u_DECODE/u510  (\u_DECODE/n26 [10], \u_DECODE/n23 [10], \u_DECODE/n25 [10]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u511  (\u_DECODE/n26 [11], \u_DECODE/n23 [11], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u512  (\u_DECODE/n26 [12], \u_DECODE/n24 [12], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u513  (\u_DECODE/n26 [13], \u_DECODE/n24 [13], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u514  (\u_DECODE/n26 [14], \u_DECODE/n24 [14], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u515  (\u_DECODE/n26 [15], \u_DECODE/n24 [15], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u516  (\u_DECODE/n26 [16], \u_DECODE/n24 [16], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u517  (\u_DECODE/n26 [17], \u_DECODE/n24 [17], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u518  (\u_DECODE/n26 [18], \u_DECODE/n24 [18], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u519  (\u_DECODE/n26 [19], \u_DECODE/n24 [19], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u52  (\u_DECODE/n8 , \u_DECODE/opc_opimm , \u_DECODE/func_001 );  // ../RTL/core/decode.v(146)
  or \u_DECODE/u520  (\u_DECODE/n26 [20], \u_DECODE/n24 [20], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u521  (\u_DECODE/n26 [21], \u_DECODE/n24 [21], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u522  (\u_DECODE/n26 [22], \u_DECODE/n24 [22], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u523  (\u_DECODE/n26 [23], \u_DECODE/n24 [23], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u524  (\u_DECODE/n26 [24], \u_DECODE/n24 [24], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u525  (\u_DECODE/n26 [25], \u_DECODE/n24 [25], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u526  (\u_DECODE/n26 [26], \u_DECODE/n24 [26], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u527  (\u_DECODE/n26 [27], \u_DECODE/n24 [27], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u528  (\u_DECODE/n26 [28], \u_DECODE/n24 [28], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u529  (\u_DECODE/n26 [29], \u_DECODE/n24 [29], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u53  (\u_DECODE/inst_slli , \u_DECODE/n8 , \u_DECODE/func7_0000000 );  // ../RTL/core/decode.v(146)
  or \u_DECODE/u530  (\u_DECODE/n26 [30], \u_DECODE/n24 [30], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u531  (\u_DECODE/n26 [31], \u_DECODE/n24 [31], \u_DECODE/n25 [11]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u532  (\u_DECODE/n25 [1], \u_DECODE/opc_store , i_data[8]);  // ../RTL/core/decode.v(208)
  and \u_DECODE/u533  (\u_DECODE/n25 [2], \u_DECODE/opc_store , i_data[9]);  // ../RTL/core/decode.v(208)
  and \u_DECODE/u534  (\u_DECODE/n25 [3], \u_DECODE/opc_store , i_data[10]);  // ../RTL/core/decode.v(208)
  and \u_DECODE/u535  (\u_DECODE/n25 [4], \u_DECODE/opc_store , i_data[11]);  // ../RTL/core/decode.v(208)
  and \u_DECODE/u536  (\u_DECODE/n25 [5], \u_DECODE/opc_store , i_data[25]);  // ../RTL/core/decode.v(208)
  and \u_DECODE/u537  (\u_DECODE/n25 [6], \u_DECODE/opc_store , i_data[26]);  // ../RTL/core/decode.v(208)
  and \u_DECODE/u538  (\u_DECODE/n25 [7], \u_DECODE/opc_store , i_data[27]);  // ../RTL/core/decode.v(208)
  and \u_DECODE/u539  (\u_DECODE/n25 [8], \u_DECODE/opc_store , i_data[28]);  // ../RTL/core/decode.v(208)
  and \u_DECODE/u54  (\u_DECODE/n9 , \u_DECODE/opc_opimm , \u_DECODE/func_101 );  // ../RTL/core/decode.v(147)
  and \u_DECODE/u540  (\u_DECODE/n25 [9], \u_DECODE/opc_store , i_data[29]);  // ../RTL/core/decode.v(208)
  and \u_DECODE/u541  (\u_DECODE/n25 [10], \u_DECODE/opc_store , i_data[30]);  // ../RTL/core/decode.v(208)
  and \u_DECODE/u542  (\u_DECODE/n25 [11], \u_DECODE/opc_store , i_data[31]);  // ../RTL/core/decode.v(208)
  and \u_DECODE/u55  (\u_DECODE/inst_srli , \u_DECODE/n9 , \u_DECODE/func7_0000000 );  // ../RTL/core/decode.v(147)
  or \u_DECODE/u56  (\u_DECODE/n6 [31], \u_DECODE/n4 [31], \u_DECODE/n5 [31]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u57  (\u_DECODE/inst_srai , \u_DECODE/n9 , \u_DECODE/func7_0100000 );  // ../RTL/core/decode.v(148)
  or \u_DECODE/u574  (\u_DECODE/n24 [12], \u_DECODE/n22 [12], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u575  (\u_DECODE/n24 [13], \u_DECODE/n22 [13], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u576  (\u_DECODE/n24 [14], \u_DECODE/n22 [14], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u577  (\u_DECODE/n24 [15], \u_DECODE/n22 [15], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u578  (\u_DECODE/n24 [16], \u_DECODE/n22 [16], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u579  (\u_DECODE/n24 [17], \u_DECODE/n22 [17], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u58  (\u_DECODE/n10 , \u_DECODE/opc_op , \u_DECODE/func_000 );  // ../RTL/core/decode.v(150)
  or \u_DECODE/u580  (\u_DECODE/n24 [18], \u_DECODE/n22 [18], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u581  (\u_DECODE/n24 [19], \u_DECODE/n22 [19], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u582  (\u_DECODE/n24 [20], \u_DECODE/n22 [20], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u583  (\u_DECODE/n24 [21], \u_DECODE/n22 [21], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u584  (\u_DECODE/n24 [22], \u_DECODE/n22 [22], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u585  (\u_DECODE/n24 [23], \u_DECODE/n22 [23], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u586  (\u_DECODE/n24 [24], \u_DECODE/n22 [24], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u587  (\u_DECODE/n24 [25], \u_DECODE/n22 [25], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u588  (\u_DECODE/n24 [26], \u_DECODE/n22 [26], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u589  (\u_DECODE/n24 [27], \u_DECODE/n22 [27], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u59  (\u_DECODE/inst_add , \u_DECODE/n10 , \u_DECODE/func7_0000000 );  // ../RTL/core/decode.v(150)
  or \u_DECODE/u590  (\u_DECODE/n24 [28], \u_DECODE/n22 [28], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u591  (\u_DECODE/n24 [29], \u_DECODE/n22 [29], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u592  (\u_DECODE/n24 [30], \u_DECODE/n22 [30], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u593  (\u_DECODE/n24 [31], \u_DECODE/n22 [31], \u_DECODE/n23 [12]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u594  (\u_DECODE/n66 [1], o_decinfo_grp[1], \u_DECODE/opc_store );  // ../RTL/core/decode.v(337)
  and \u_DECODE/u595  (\u_DECODE/n66 [2], o_decinfo_grp[1], \u_DECODE/lsuinfo [2]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u596  (\u_DECODE/n66 [3], o_decinfo_grp[1], \u_DECODE/lsuinfo [3]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u597  (\u_DECODE/n66 [4], o_decinfo_grp[1], \u_DECODE/func_010 );  // ../RTL/core/decode.v(337)
  and \u_DECODE/u598  (\u_DECODE/n66 [5], o_decinfo_grp[1], \u_DECODE/lsuinfo [5]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u6  (o_decinfo[2], \u_DECODE/n71 [2], \u_DECODE/n72 [2]);  // ../RTL/core/decode.v(337)
  or \u_DECODE/u60  (\u_DECODE/n6 [19], \u_DECODE/n4 [19], \u_DECODE/n5 [31]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u604  (\u_DECODE/n65 [1], o_decinfo_grp[0], \u_DECODE/inst_sub );  // ../RTL/core/decode.v(337)
  and \u_DECODE/u605  (\u_DECODE/n65 [2], o_decinfo_grp[0], \u_DECODE/aluinfo [2]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u606  (\u_DECODE/n65 [3], o_decinfo_grp[0], \u_DECODE/aluinfo [3]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u607  (\u_DECODE/n65 [4], o_decinfo_grp[0], \u_DECODE/aluinfo [4]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u608  (\u_DECODE/n65 [5], o_decinfo_grp[0], \u_DECODE/aluinfo [5]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u609  (\u_DECODE/n65 [6], o_decinfo_grp[0], \u_DECODE/aluinfo [6]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u61  (\u_DECODE/inst_sub , \u_DECODE/n10 , \u_DECODE/func7_0100000 );  // ../RTL/core/decode.v(151)
  and \u_DECODE/u610  (\u_DECODE/n65 [7], o_decinfo_grp[0], \u_DECODE/aluinfo [7]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u611  (\u_DECODE/n65 [8], o_decinfo_grp[0], \u_DECODE/aluinfo [8]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u612  (\u_DECODE/n65 [9], o_decinfo_grp[0], \u_DECODE/aluinfo [9]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u62  (\u_DECODE/n11 , \u_DECODE/opc_op , \u_DECODE/func_001 );  // ../RTL/core/decode.v(152)
  and \u_DECODE/u63  (\u_DECODE/inst_sll , \u_DECODE/n11 , \u_DECODE/func7_0000000 );  // ../RTL/core/decode.v(152)
  and \u_DECODE/u64  (\u_DECODE/n12 , \u_DECODE/opc_op , \u_DECODE/func_010 );  // ../RTL/core/decode.v(153)
  and \u_DECODE/u65  (\u_DECODE/inst_slt , \u_DECODE/n12 , \u_DECODE/func7_0000000 );  // ../RTL/core/decode.v(153)
  and \u_DECODE/u66  (\u_DECODE/n13 , \u_DECODE/opc_op , \u_DECODE/func_011 );  // ../RTL/core/decode.v(154)
  and \u_DECODE/u67  (\u_DECODE/inst_sltu , \u_DECODE/n13 , \u_DECODE/func7_0000000 );  // ../RTL/core/decode.v(154)
  and \u_DECODE/u68  (\u_DECODE/n14 , \u_DECODE/opc_op , \u_DECODE/func_100 );  // ../RTL/core/decode.v(155)
  and \u_DECODE/u69  (\u_DECODE/inst_xor , \u_DECODE/n14 , \u_DECODE/func7_0000000 );  // ../RTL/core/decode.v(155)
  AL_MUX \u_DECODE/u7  (
    .i0(1'b0),
    .i1(\u_DECODE/n2 ),
    .sel(\u_DECODE/n0 ),
    .o(inst_jalr));  // ../RTL/core/decode.v(56)
  and \u_DECODE/u70  (\u_DECODE/n15 , \u_DECODE/opc_op , \u_DECODE/func_101 );  // ../RTL/core/decode.v(156)
  and \u_DECODE/u71  (\u_DECODE/inst_srl , \u_DECODE/n15 , \u_DECODE/func7_0000000 );  // ../RTL/core/decode.v(156)
  or \u_DECODE/u72  (\u_DECODE/n6 [18], \u_DECODE/n4 [18], \u_DECODE/n5 [31]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u73  (\u_DECODE/inst_sra , \u_DECODE/n15 , \u_DECODE/func7_0100000 );  // ../RTL/core/decode.v(157)
  and \u_DECODE/u74  (\u_DECODE/n16 , \u_DECODE/opc_op , \u_DECODE/func_110 );  // ../RTL/core/decode.v(158)
  and \u_DECODE/u75  (\u_DECODE/inst_or , \u_DECODE/n16 , \u_DECODE/func7_0000000 );  // ../RTL/core/decode.v(158)
  and \u_DECODE/u76  (\u_DECODE/n17 , \u_DECODE/opc_op , \u_DECODE/func_111 );  // ../RTL/core/decode.v(159)
  and \u_DECODE/u77  (\u_DECODE/inst_and , \u_DECODE/n17 , \u_DECODE/func7_0000000 );  // ../RTL/core/decode.v(159)
  or \u_DECODE/u8  (o_decinfo[1], \u_DECODE/n71 [1], \u_DECODE/n72 [1]);  // ../RTL/core/decode.v(337)
  and \u_DECODE/u80  (\u_DECODE/n18 , o_decinfo_grp[4], \u_DECODE/func_000 );  // ../RTL/core/decode.v(164)
  and \u_DECODE/u81  (\u_DECODE/inst_ecall , \u_DECODE/n18 , \u_DECODE/type_i_imm_000000000000 );  // ../RTL/core/decode.v(164)
  or \u_DECODE/u82  (\u_DECODE/n6 [17], \u_DECODE/n4 [17], \u_DECODE/n5 [31]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u83  (\u_DECODE/inst_ebreak , \u_DECODE/n18 , \u_DECODE/type_i_imm_000000000001 );  // ../RTL/core/decode.v(165)
  and \u_DECODE/u84  (\u_DECODE/inst_csrrw , o_decinfo_grp[4], \u_DECODE/func_001 );  // ../RTL/core/decode.v(166)
  and \u_DECODE/u85  (\u_DECODE/inst_csrrs , o_decinfo_grp[4], \u_DECODE/func_010 );  // ../RTL/core/decode.v(167)
  and \u_DECODE/u86  (\u_DECODE/inst_csrrc , o_decinfo_grp[4], \u_DECODE/func_011 );  // ../RTL/core/decode.v(168)
  and \u_DECODE/u87  (\u_DECODE/inst_csrrwi , o_decinfo_grp[4], \u_DECODE/func_101 );  // ../RTL/core/decode.v(169)
  and \u_DECODE/u88  (\u_DECODE/inst_csrrsi , o_decinfo_grp[4], \u_DECODE/func_110 );  // ../RTL/core/decode.v(170)
  and \u_DECODE/u89  (\u_DECODE/inst_csrrci , o_decinfo_grp[4], \u_DECODE/func_111 );  // ../RTL/core/decode.v(171)
  AL_MUX \u_DECODE/u9  (
    .i0(1'b0),
    .i1(\u_DECODE/n3 ),
    .sel(\u_DECODE/n0 ),
    .o(inst_bxx));  // ../RTL/core/decode.v(57)
  or \u_DECODE/u90  (\u_DECODE/n6 [16], \u_DECODE/n4 [16], \u_DECODE/n5 [31]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u91  (\u_DECODE/inst_mul , \u_DECODE/n10 , \u_DECODE/func7_0000001 );  // ../RTL/core/decode.v(174)
  or \u_DECODE/u92  (\u_DECODE/n6 [15], \u_DECODE/n4 [15], \u_DECODE/n5 [31]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u923  (bp_imm[1], \u_DECODE/n6 [1], \u_DECODE/n7 [1]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u924  (bp_imm[2], \u_DECODE/n6 [2], \u_DECODE/n7 [2]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u925  (bp_imm[3], \u_DECODE/n6 [3], \u_DECODE/n7 [3]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u926  (bp_imm[4], \u_DECODE/n6 [4], \u_DECODE/n7 [4]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u927  (bp_imm[5], \u_DECODE/n6 [5], \u_DECODE/n7 [5]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u928  (bp_imm[6], \u_DECODE/n6 [6], \u_DECODE/n7 [6]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u929  (bp_imm[7], \u_DECODE/n6 [7], \u_DECODE/n7 [7]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u93  (\u_DECODE/inst_mulh , \u_DECODE/n11 , \u_DECODE/func7_0000001 );  // ../RTL/core/decode.v(175)
  or \u_DECODE/u930  (bp_imm[8], \u_DECODE/n6 [8], \u_DECODE/n7 [8]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u931  (bp_imm[9], \u_DECODE/n6 [9], \u_DECODE/n7 [9]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u932  (bp_imm[10], \u_DECODE/n6 [10], \u_DECODE/n7 [10]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u933  (bp_imm[11], \u_DECODE/n6 [11], \u_DECODE/n7 [11]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u934  (bp_imm[12], \u_DECODE/n6 [12], \u_DECODE/n7 [31]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u935  (bp_imm[13], \u_DECODE/n6 [13], \u_DECODE/n7 [31]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u936  (bp_imm[14], \u_DECODE/n6 [14], \u_DECODE/n7 [31]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u937  (bp_imm[15], \u_DECODE/n6 [15], \u_DECODE/n7 [31]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u938  (bp_imm[16], \u_DECODE/n6 [16], \u_DECODE/n7 [31]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u939  (bp_imm[17], \u_DECODE/n6 [17], \u_DECODE/n7 [31]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u94  (\u_DECODE/n6 [14], \u_DECODE/n4 [14], \u_DECODE/n5 [31]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u940  (bp_imm[18], \u_DECODE/n6 [18], \u_DECODE/n7 [31]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u941  (bp_imm[19], \u_DECODE/n6 [19], \u_DECODE/n7 [31]);  // ../RTL/core/decode.v(62)
  or \u_DECODE/u942  (bp_imm[31], \u_DECODE/n6 [31], \u_DECODE/n7 [31]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u95  (\u_DECODE/inst_mulhsu , \u_DECODE/n12 , \u_DECODE/func7_0000001 );  // ../RTL/core/decode.v(176)
  and \u_DECODE/u954  (\u_DECODE/n23 [1], \u_DECODE/n3 , i_data[8]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u955  (\u_DECODE/n23 [2], \u_DECODE/n3 , i_data[9]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u956  (\u_DECODE/n23 [3], \u_DECODE/n3 , i_data[10]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u957  (\u_DECODE/n23 [4], \u_DECODE/n3 , i_data[11]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u958  (\u_DECODE/n23 [5], \u_DECODE/n3 , i_data[25]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u959  (\u_DECODE/n23 [6], \u_DECODE/n3 , i_data[26]);  // ../RTL/core/decode.v(206)
  or \u_DECODE/u96  (\u_DECODE/n6 [13], \u_DECODE/n4 [13], \u_DECODE/n5 [31]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u960  (\u_DECODE/n23 [7], \u_DECODE/n3 , i_data[27]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u961  (\u_DECODE/n23 [8], \u_DECODE/n3 , i_data[28]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u962  (\u_DECODE/n23 [9], \u_DECODE/n3 , i_data[29]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u963  (\u_DECODE/n23 [10], \u_DECODE/n3 , i_data[30]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u964  (\u_DECODE/n23 [11], \u_DECODE/n3 , i_data[7]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u965  (\u_DECODE/n23 [12], \u_DECODE/n3 , i_data[31]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u97  (\u_DECODE/inst_mulhu , \u_DECODE/n13 , \u_DECODE/func7_0000001 );  // ../RTL/core/decode.v(177)
  or \u_DECODE/u98  (\u_DECODE/n6 [12], \u_DECODE/n4 [12], \u_DECODE/n5 [31]);  // ../RTL/core/decode.v(62)
  and \u_DECODE/u99  (\u_DECODE/inst_div , \u_DECODE/n14 , \u_DECODE/func7_0000001 );  // ../RTL/core/decode.v(178)
  and \u_DECODE/u997  (\u_DECODE/n22 [12], \u_DECODE/n21 , i_data[12]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u998  (\u_DECODE/n22 [13], \u_DECODE/n21 , i_data[13]);  // ../RTL/core/decode.v(206)
  and \u_DECODE/u999  (\u_DECODE/n22 [14], \u_DECODE/n21 , i_data[14]);  // ../RTL/core/decode.v(206)
  REGFILE u_REGFILE (
    .i_clk(i_clk),
    .i_rd_wdata(i_rd_wdata),
    .i_rdidx(i_rdidx),
    .i_rdwen(i_rdwen),
    .i_rs1idx(i_data[19:15]),
    .i_rs1ren(rs1ren),
    .i_rs2idx(i_data[24:20]),
    .i_rs2ren(rs2ren),
    .i_rstn(1'b0),
    .o_rs1_rdata(rs1_rdata),
    .o_rs2_rdata(o_rs2rdata));  // ../RTL/core/bpu.v(186)

endmodule 

module CSR_REGFILE  // ../RTL/core/csr_regfile.v(21)
  (
  i_clk,
  i_csr_ren,
  i_csr_ridx,
  i_csr_wdata,
  i_csr_wen,
  i_csr_widx,
  i_rstn,
  o_csr_rdata
  );

  input i_clk;  // ../RTL/core/csr_regfile.v(22)
  input i_csr_ren;  // ../RTL/core/csr_regfile.v(26)
  input [11:0] i_csr_ridx;  // ../RTL/core/csr_regfile.v(27)
  input [31:0] i_csr_wdata;  // ../RTL/core/csr_regfile.v(32)
  input i_csr_wen;  // ../RTL/core/csr_regfile.v(30)
  input [11:0] i_csr_widx;  // ../RTL/core/csr_regfile.v(31)
  input i_rstn;  // ../RTL/core/csr_regfile.v(23)
  output [31:0] o_csr_rdata;  // ../RTL/core/csr_regfile.v(28)

  wire [31:0] fctrl;  // ../RTL/core/csr_regfile.v(128)
  wire [31:0] fop1;  // ../RTL/core/csr_regfile.v(129)
  wire [31:0] fop2;  // ../RTL/core/csr_regfile.v(130)
  wire [31:0] fres;  // ../RTL/core/csr_regfile.v(134)
  wire [31:0] fres0_add;  // ../RTL/core/csr_regfile.v(131)
  wire [31:0] fres0_mul;  // ../RTL/core/csr_regfile.v(133)
  wire [31:0] fres0_sub;  // ../RTL/core/csr_regfile.v(132)
  wire [31:2] mtvec_base;  // ../RTL/core/csr_regfile.v(60)
  wire [1:0] mtvec_mode;  // ../RTL/core/csr_regfile.v(61)
  wire  \mux17_oh_b0/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b0/B6 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b0/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b0/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b0/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b1/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b1/B6 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b1/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b1/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b1/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b10/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b10/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b10/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b10/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b11/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b11/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b11/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b11/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b12/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b12/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b12/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b12/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b13/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b13/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b13/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b13/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b14/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b14/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b14/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b14/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b15/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b15/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b15/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b15/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b16/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b16/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b16/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b16/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b17/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b17/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b17/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b17/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b18/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b18/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b18/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b18/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b19/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b19/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b19/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b19/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b2/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b2/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b2/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b2/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b20/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b20/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b20/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b20/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b21/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b21/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b21/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b21/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b22/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b22/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b22/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b22/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b23/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b23/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b23/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b23/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b24/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b24/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b24/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b24/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b25/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b25/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b25/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b25/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b26/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b26/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b26/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b26/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b27/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b27/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b27/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b27/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b28/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b28/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b28/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b28/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b29/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b29/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b29/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b29/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b3/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b3/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b3/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b3/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b30/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b30/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b30/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b30/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b31/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b31/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b31/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b31/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b4/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b4/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b4/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b4/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b5/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b5/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b5/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b5/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b6/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b6/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b6/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b6/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b7/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b7/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b7/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b7/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b8/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b8/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b8/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b8/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b9/B2 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b9/B7 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b9/B8 ;  // ../RTL/core/csr_regfile.v(170)
  wire  \mux17_oh_b9/B9 ;  // ../RTL/core/csr_regfile.v(170)
  wire [31:0] n39;
  wire \mux17_oh_b0/or_B6_B7_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b0/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b0/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b1/or_B6_B7_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b1/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b1/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b10/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b10/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b11/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b11/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b12/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b12/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b13/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b13/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b14/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b14/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b15/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b15/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b16/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b16/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b17/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b17/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b18/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b18/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b19/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b19/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b2/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b2/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b20/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b20/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b21/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b21/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b22/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b22/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b23/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b23/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b24/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b24/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b25/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b25/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b26/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b26/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b27/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b27/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b28/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b28/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b29/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b29/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b3/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b3/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b30/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b30/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b31/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b31/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b4/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b4/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b5/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b5/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b6/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b6/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b7/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b7/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b8/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b8/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b9/or_B8_or_B9_B10_o_o ;  // ../RTL/core/csr_regfile.v(170)
  wire \mux17_oh_b9/or_or_B5_or_B6_B7_o__o ;  // ../RTL/core/csr_regfile.v(170)
  wire n0;
  wire n1;
  wire n10;
  wire n11;
  wire n13;
  wire n14;
  wire n16;
  wire n17;
  wire n19;
  wire n22;
  wire n26;
  wire n27;
  wire n28;
  wire n29;

  eq_w12 eq0 (
    .i0(i_csr_widx),
    .i1(12'b001100000101),
    .o(n0));  // ../RTL/core/csr_regfile.v(68)
  eq_w12 eq13 (
    .i0(i_csr_ridx),
    .i1(12'b001100010000),
    .o(n26));  // ../RTL/core/csr_regfile.v(177)
  eq_w12 eq14 (
    .i0(i_csr_ridx),
    .i1(12'b001100010001),
    .o(n27));  // ../RTL/core/csr_regfile.v(178)
  eq_w12 eq15 (
    .i0(i_csr_ridx),
    .i1(12'b001100010010),
    .o(n28));  // ../RTL/core/csr_regfile.v(179)
  eq_w12 eq16 (
    .i0(i_csr_ridx),
    .i1(12'b001100010011),
    .o(n29));  // ../RTL/core/csr_regfile.v(180)
  eq_w12 eq4 (
    .i0(i_csr_widx),
    .i1(12'b001100010000),
    .o(n10));  // ../RTL/core/csr_regfile.v(144)
  eq_w12 eq5 (
    .i0(i_csr_widx),
    .i1(12'b001100010010),
    .o(n13));  // ../RTL/core/csr_regfile.v(147)
  eq_w12 eq6 (
    .i0(i_csr_widx),
    .i1(12'b001100010011),
    .o(n16));  // ../RTL/core/csr_regfile.v(150)
  eq_w12 eq9 (
    .i0(i_csr_ridx),
    .i1(12'b001100000101),
    .o(n22));  // ../RTL/core/csr_regfile.v(172)
  and \mux17_oh_b0/and_b0_2  (\mux17_oh_b0/B2 , mtvec_mode[0], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b0/and_b0_6  (\mux17_oh_b0/B6 , fctrl[0], n26);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b0/and_b0_7  (\mux17_oh_b0/B7 , fres[0], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b0/and_b0_8  (\mux17_oh_b0/B8 , fop1[0], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b0/and_b0_9  (\mux17_oh_b0/B9 , fop2[0], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b0/or_B6_B7  (\mux17_oh_b0/or_B6_B7_o , \mux17_oh_b0/B6 , \mux17_oh_b0/B7 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b0/or_B8_or_B9_B10_o  (\mux17_oh_b0/or_B8_or_B9_B10_o_o , \mux17_oh_b0/B8 , \mux17_oh_b0/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b0/or_or_B5_or_B6_B7_o_  (\mux17_oh_b0/or_or_B5_or_B6_B7_o__o , \mux17_oh_b0/or_B6_B7_o , \mux17_oh_b0/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b0/or_or_or_B0_B1_o_or_  (n39[0], \mux17_oh_b0/B2 , \mux17_oh_b0/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b1/and_b0_2  (\mux17_oh_b1/B2 , mtvec_mode[1], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b1/and_b0_6  (\mux17_oh_b1/B6 , fctrl[1], n26);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b1/and_b0_7  (\mux17_oh_b1/B7 , fres[1], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b1/and_b0_8  (\mux17_oh_b1/B8 , fop1[1], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b1/and_b0_9  (\mux17_oh_b1/B9 , fop2[1], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b1/or_B6_B7  (\mux17_oh_b1/or_B6_B7_o , \mux17_oh_b1/B6 , \mux17_oh_b1/B7 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b1/or_B8_or_B9_B10_o  (\mux17_oh_b1/or_B8_or_B9_B10_o_o , \mux17_oh_b1/B8 , \mux17_oh_b1/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b1/or_or_B5_or_B6_B7_o_  (\mux17_oh_b1/or_or_B5_or_B6_B7_o__o , \mux17_oh_b1/or_B6_B7_o , \mux17_oh_b1/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b1/or_or_or_B0_B1_o_or_  (n39[1], \mux17_oh_b1/B2 , \mux17_oh_b1/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b10/and_b0_2  (\mux17_oh_b10/B2 , mtvec_base[10], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b10/and_b0_7  (\mux17_oh_b10/B7 , fres[10], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b10/and_b0_8  (\mux17_oh_b10/B8 , fop1[10], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b10/and_b0_9  (\mux17_oh_b10/B9 , fop2[10], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b10/or_B8_or_B9_B10_o  (\mux17_oh_b10/or_B8_or_B9_B10_o_o , \mux17_oh_b10/B8 , \mux17_oh_b10/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b10/or_or_B5_or_B6_B7_o_  (\mux17_oh_b10/or_or_B5_or_B6_B7_o__o , \mux17_oh_b10/B7 , \mux17_oh_b10/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b10/or_or_or_B0_B1_o_or_  (n39[10], \mux17_oh_b10/B2 , \mux17_oh_b10/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b11/and_b0_2  (\mux17_oh_b11/B2 , mtvec_base[11], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b11/and_b0_7  (\mux17_oh_b11/B7 , fres[11], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b11/and_b0_8  (\mux17_oh_b11/B8 , fop1[11], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b11/and_b0_9  (\mux17_oh_b11/B9 , fop2[11], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b11/or_B8_or_B9_B10_o  (\mux17_oh_b11/or_B8_or_B9_B10_o_o , \mux17_oh_b11/B8 , \mux17_oh_b11/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b11/or_or_B5_or_B6_B7_o_  (\mux17_oh_b11/or_or_B5_or_B6_B7_o__o , \mux17_oh_b11/B7 , \mux17_oh_b11/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b11/or_or_or_B0_B1_o_or_  (n39[11], \mux17_oh_b11/B2 , \mux17_oh_b11/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b12/and_b0_2  (\mux17_oh_b12/B2 , mtvec_base[12], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b12/and_b0_7  (\mux17_oh_b12/B7 , fres[12], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b12/and_b0_8  (\mux17_oh_b12/B8 , fop1[12], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b12/and_b0_9  (\mux17_oh_b12/B9 , fop2[12], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b12/or_B8_or_B9_B10_o  (\mux17_oh_b12/or_B8_or_B9_B10_o_o , \mux17_oh_b12/B8 , \mux17_oh_b12/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b12/or_or_B5_or_B6_B7_o_  (\mux17_oh_b12/or_or_B5_or_B6_B7_o__o , \mux17_oh_b12/B7 , \mux17_oh_b12/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b12/or_or_or_B0_B1_o_or_  (n39[12], \mux17_oh_b12/B2 , \mux17_oh_b12/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b13/and_b0_2  (\mux17_oh_b13/B2 , mtvec_base[13], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b13/and_b0_7  (\mux17_oh_b13/B7 , fres[13], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b13/and_b0_8  (\mux17_oh_b13/B8 , fop1[13], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b13/and_b0_9  (\mux17_oh_b13/B9 , fop2[13], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b13/or_B8_or_B9_B10_o  (\mux17_oh_b13/or_B8_or_B9_B10_o_o , \mux17_oh_b13/B8 , \mux17_oh_b13/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b13/or_or_B5_or_B6_B7_o_  (\mux17_oh_b13/or_or_B5_or_B6_B7_o__o , \mux17_oh_b13/B7 , \mux17_oh_b13/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b13/or_or_or_B0_B1_o_or_  (n39[13], \mux17_oh_b13/B2 , \mux17_oh_b13/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b14/and_b0_2  (\mux17_oh_b14/B2 , mtvec_base[14], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b14/and_b0_7  (\mux17_oh_b14/B7 , fres[14], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b14/and_b0_8  (\mux17_oh_b14/B8 , fop1[14], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b14/and_b0_9  (\mux17_oh_b14/B9 , fop2[14], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b14/or_B8_or_B9_B10_o  (\mux17_oh_b14/or_B8_or_B9_B10_o_o , \mux17_oh_b14/B8 , \mux17_oh_b14/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b14/or_or_B5_or_B6_B7_o_  (\mux17_oh_b14/or_or_B5_or_B6_B7_o__o , \mux17_oh_b14/B7 , \mux17_oh_b14/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b14/or_or_or_B0_B1_o_or_  (n39[14], \mux17_oh_b14/B2 , \mux17_oh_b14/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b15/and_b0_2  (\mux17_oh_b15/B2 , mtvec_base[15], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b15/and_b0_7  (\mux17_oh_b15/B7 , fres[15], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b15/and_b0_8  (\mux17_oh_b15/B8 , fop1[15], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b15/and_b0_9  (\mux17_oh_b15/B9 , fop2[15], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b15/or_B8_or_B9_B10_o  (\mux17_oh_b15/or_B8_or_B9_B10_o_o , \mux17_oh_b15/B8 , \mux17_oh_b15/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b15/or_or_B5_or_B6_B7_o_  (\mux17_oh_b15/or_or_B5_or_B6_B7_o__o , \mux17_oh_b15/B7 , \mux17_oh_b15/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b15/or_or_or_B0_B1_o_or_  (n39[15], \mux17_oh_b15/B2 , \mux17_oh_b15/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b16/and_b0_2  (\mux17_oh_b16/B2 , mtvec_base[16], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b16/and_b0_7  (\mux17_oh_b16/B7 , fres[16], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b16/and_b0_8  (\mux17_oh_b16/B8 , fop1[16], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b16/and_b0_9  (\mux17_oh_b16/B9 , fop2[16], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b16/or_B8_or_B9_B10_o  (\mux17_oh_b16/or_B8_or_B9_B10_o_o , \mux17_oh_b16/B8 , \mux17_oh_b16/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b16/or_or_B5_or_B6_B7_o_  (\mux17_oh_b16/or_or_B5_or_B6_B7_o__o , \mux17_oh_b16/B7 , \mux17_oh_b16/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b16/or_or_or_B0_B1_o_or_  (n39[16], \mux17_oh_b16/B2 , \mux17_oh_b16/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b17/and_b0_2  (\mux17_oh_b17/B2 , mtvec_base[17], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b17/and_b0_7  (\mux17_oh_b17/B7 , fres[17], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b17/and_b0_8  (\mux17_oh_b17/B8 , fop1[17], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b17/and_b0_9  (\mux17_oh_b17/B9 , fop2[17], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b17/or_B8_or_B9_B10_o  (\mux17_oh_b17/or_B8_or_B9_B10_o_o , \mux17_oh_b17/B8 , \mux17_oh_b17/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b17/or_or_B5_or_B6_B7_o_  (\mux17_oh_b17/or_or_B5_or_B6_B7_o__o , \mux17_oh_b17/B7 , \mux17_oh_b17/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b17/or_or_or_B0_B1_o_or_  (n39[17], \mux17_oh_b17/B2 , \mux17_oh_b17/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b18/and_b0_2  (\mux17_oh_b18/B2 , mtvec_base[18], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b18/and_b0_7  (\mux17_oh_b18/B7 , fres[18], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b18/and_b0_8  (\mux17_oh_b18/B8 , fop1[18], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b18/and_b0_9  (\mux17_oh_b18/B9 , fop2[18], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b18/or_B8_or_B9_B10_o  (\mux17_oh_b18/or_B8_or_B9_B10_o_o , \mux17_oh_b18/B8 , \mux17_oh_b18/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b18/or_or_B5_or_B6_B7_o_  (\mux17_oh_b18/or_or_B5_or_B6_B7_o__o , \mux17_oh_b18/B7 , \mux17_oh_b18/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b18/or_or_or_B0_B1_o_or_  (n39[18], \mux17_oh_b18/B2 , \mux17_oh_b18/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b19/and_b0_2  (\mux17_oh_b19/B2 , mtvec_base[19], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b19/and_b0_7  (\mux17_oh_b19/B7 , fres[19], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b19/and_b0_8  (\mux17_oh_b19/B8 , fop1[19], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b19/and_b0_9  (\mux17_oh_b19/B9 , fop2[19], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b19/or_B8_or_B9_B10_o  (\mux17_oh_b19/or_B8_or_B9_B10_o_o , \mux17_oh_b19/B8 , \mux17_oh_b19/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b19/or_or_B5_or_B6_B7_o_  (\mux17_oh_b19/or_or_B5_or_B6_B7_o__o , \mux17_oh_b19/B7 , \mux17_oh_b19/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b19/or_or_or_B0_B1_o_or_  (n39[19], \mux17_oh_b19/B2 , \mux17_oh_b19/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b2/and_b0_2  (\mux17_oh_b2/B2 , mtvec_base[2], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b2/and_b0_7  (\mux17_oh_b2/B7 , fres[2], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b2/and_b0_8  (\mux17_oh_b2/B8 , fop1[2], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b2/and_b0_9  (\mux17_oh_b2/B9 , fop2[2], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b2/or_B8_or_B9_B10_o  (\mux17_oh_b2/or_B8_or_B9_B10_o_o , \mux17_oh_b2/B8 , \mux17_oh_b2/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b2/or_or_B5_or_B6_B7_o_  (\mux17_oh_b2/or_or_B5_or_B6_B7_o__o , \mux17_oh_b2/B7 , \mux17_oh_b2/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b2/or_or_or_B0_B1_o_or_  (n39[2], \mux17_oh_b2/B2 , \mux17_oh_b2/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b20/and_b0_2  (\mux17_oh_b20/B2 , mtvec_base[20], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b20/and_b0_7  (\mux17_oh_b20/B7 , fres[20], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b20/and_b0_8  (\mux17_oh_b20/B8 , fop1[20], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b20/and_b0_9  (\mux17_oh_b20/B9 , fop2[20], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b20/or_B8_or_B9_B10_o  (\mux17_oh_b20/or_B8_or_B9_B10_o_o , \mux17_oh_b20/B8 , \mux17_oh_b20/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b20/or_or_B5_or_B6_B7_o_  (\mux17_oh_b20/or_or_B5_or_B6_B7_o__o , \mux17_oh_b20/B7 , \mux17_oh_b20/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b20/or_or_or_B0_B1_o_or_  (n39[20], \mux17_oh_b20/B2 , \mux17_oh_b20/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b21/and_b0_2  (\mux17_oh_b21/B2 , mtvec_base[21], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b21/and_b0_7  (\mux17_oh_b21/B7 , fres[21], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b21/and_b0_8  (\mux17_oh_b21/B8 , fop1[21], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b21/and_b0_9  (\mux17_oh_b21/B9 , fop2[21], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b21/or_B8_or_B9_B10_o  (\mux17_oh_b21/or_B8_or_B9_B10_o_o , \mux17_oh_b21/B8 , \mux17_oh_b21/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b21/or_or_B5_or_B6_B7_o_  (\mux17_oh_b21/or_or_B5_or_B6_B7_o__o , \mux17_oh_b21/B7 , \mux17_oh_b21/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b21/or_or_or_B0_B1_o_or_  (n39[21], \mux17_oh_b21/B2 , \mux17_oh_b21/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b22/and_b0_2  (\mux17_oh_b22/B2 , mtvec_base[22], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b22/and_b0_7  (\mux17_oh_b22/B7 , fres[22], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b22/and_b0_8  (\mux17_oh_b22/B8 , fop1[22], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b22/and_b0_9  (\mux17_oh_b22/B9 , fop2[22], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b22/or_B8_or_B9_B10_o  (\mux17_oh_b22/or_B8_or_B9_B10_o_o , \mux17_oh_b22/B8 , \mux17_oh_b22/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b22/or_or_B5_or_B6_B7_o_  (\mux17_oh_b22/or_or_B5_or_B6_B7_o__o , \mux17_oh_b22/B7 , \mux17_oh_b22/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b22/or_or_or_B0_B1_o_or_  (n39[22], \mux17_oh_b22/B2 , \mux17_oh_b22/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b23/and_b0_2  (\mux17_oh_b23/B2 , mtvec_base[23], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b23/and_b0_7  (\mux17_oh_b23/B7 , fres[23], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b23/and_b0_8  (\mux17_oh_b23/B8 , fop1[23], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b23/and_b0_9  (\mux17_oh_b23/B9 , fop2[23], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b23/or_B8_or_B9_B10_o  (\mux17_oh_b23/or_B8_or_B9_B10_o_o , \mux17_oh_b23/B8 , \mux17_oh_b23/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b23/or_or_B5_or_B6_B7_o_  (\mux17_oh_b23/or_or_B5_or_B6_B7_o__o , \mux17_oh_b23/B7 , \mux17_oh_b23/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b23/or_or_or_B0_B1_o_or_  (n39[23], \mux17_oh_b23/B2 , \mux17_oh_b23/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b24/and_b0_2  (\mux17_oh_b24/B2 , mtvec_base[24], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b24/and_b0_7  (\mux17_oh_b24/B7 , fres[24], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b24/and_b0_8  (\mux17_oh_b24/B8 , fop1[24], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b24/and_b0_9  (\mux17_oh_b24/B9 , fop2[24], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b24/or_B8_or_B9_B10_o  (\mux17_oh_b24/or_B8_or_B9_B10_o_o , \mux17_oh_b24/B8 , \mux17_oh_b24/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b24/or_or_B5_or_B6_B7_o_  (\mux17_oh_b24/or_or_B5_or_B6_B7_o__o , \mux17_oh_b24/B7 , \mux17_oh_b24/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b24/or_or_or_B0_B1_o_or_  (n39[24], \mux17_oh_b24/B2 , \mux17_oh_b24/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b25/and_b0_2  (\mux17_oh_b25/B2 , mtvec_base[25], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b25/and_b0_7  (\mux17_oh_b25/B7 , fres[25], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b25/and_b0_8  (\mux17_oh_b25/B8 , fop1[25], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b25/and_b0_9  (\mux17_oh_b25/B9 , fop2[25], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b25/or_B8_or_B9_B10_o  (\mux17_oh_b25/or_B8_or_B9_B10_o_o , \mux17_oh_b25/B8 , \mux17_oh_b25/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b25/or_or_B5_or_B6_B7_o_  (\mux17_oh_b25/or_or_B5_or_B6_B7_o__o , \mux17_oh_b25/B7 , \mux17_oh_b25/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b25/or_or_or_B0_B1_o_or_  (n39[25], \mux17_oh_b25/B2 , \mux17_oh_b25/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b26/and_b0_2  (\mux17_oh_b26/B2 , mtvec_base[26], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b26/and_b0_7  (\mux17_oh_b26/B7 , fres[26], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b26/and_b0_8  (\mux17_oh_b26/B8 , fop1[26], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b26/and_b0_9  (\mux17_oh_b26/B9 , fop2[26], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b26/or_B8_or_B9_B10_o  (\mux17_oh_b26/or_B8_or_B9_B10_o_o , \mux17_oh_b26/B8 , \mux17_oh_b26/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b26/or_or_B5_or_B6_B7_o_  (\mux17_oh_b26/or_or_B5_or_B6_B7_o__o , \mux17_oh_b26/B7 , \mux17_oh_b26/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b26/or_or_or_B0_B1_o_or_  (n39[26], \mux17_oh_b26/B2 , \mux17_oh_b26/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b27/and_b0_2  (\mux17_oh_b27/B2 , mtvec_base[27], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b27/and_b0_7  (\mux17_oh_b27/B7 , fres[27], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b27/and_b0_8  (\mux17_oh_b27/B8 , fop1[27], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b27/and_b0_9  (\mux17_oh_b27/B9 , fop2[27], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b27/or_B8_or_B9_B10_o  (\mux17_oh_b27/or_B8_or_B9_B10_o_o , \mux17_oh_b27/B8 , \mux17_oh_b27/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b27/or_or_B5_or_B6_B7_o_  (\mux17_oh_b27/or_or_B5_or_B6_B7_o__o , \mux17_oh_b27/B7 , \mux17_oh_b27/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b27/or_or_or_B0_B1_o_or_  (n39[27], \mux17_oh_b27/B2 , \mux17_oh_b27/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b28/and_b0_2  (\mux17_oh_b28/B2 , mtvec_base[28], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b28/and_b0_7  (\mux17_oh_b28/B7 , fres[28], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b28/and_b0_8  (\mux17_oh_b28/B8 , fop1[28], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b28/and_b0_9  (\mux17_oh_b28/B9 , fop2[28], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b28/or_B8_or_B9_B10_o  (\mux17_oh_b28/or_B8_or_B9_B10_o_o , \mux17_oh_b28/B8 , \mux17_oh_b28/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b28/or_or_B5_or_B6_B7_o_  (\mux17_oh_b28/or_or_B5_or_B6_B7_o__o , \mux17_oh_b28/B7 , \mux17_oh_b28/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b28/or_or_or_B0_B1_o_or_  (n39[28], \mux17_oh_b28/B2 , \mux17_oh_b28/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b29/and_b0_2  (\mux17_oh_b29/B2 , mtvec_base[29], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b29/and_b0_7  (\mux17_oh_b29/B7 , fres[29], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b29/and_b0_8  (\mux17_oh_b29/B8 , fop1[29], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b29/and_b0_9  (\mux17_oh_b29/B9 , fop2[29], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b29/or_B8_or_B9_B10_o  (\mux17_oh_b29/or_B8_or_B9_B10_o_o , \mux17_oh_b29/B8 , \mux17_oh_b29/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b29/or_or_B5_or_B6_B7_o_  (\mux17_oh_b29/or_or_B5_or_B6_B7_o__o , \mux17_oh_b29/B7 , \mux17_oh_b29/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b29/or_or_or_B0_B1_o_or_  (n39[29], \mux17_oh_b29/B2 , \mux17_oh_b29/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b3/and_b0_2  (\mux17_oh_b3/B2 , mtvec_base[3], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b3/and_b0_7  (\mux17_oh_b3/B7 , fres[3], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b3/and_b0_8  (\mux17_oh_b3/B8 , fop1[3], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b3/and_b0_9  (\mux17_oh_b3/B9 , fop2[3], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b3/or_B8_or_B9_B10_o  (\mux17_oh_b3/or_B8_or_B9_B10_o_o , \mux17_oh_b3/B8 , \mux17_oh_b3/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b3/or_or_B5_or_B6_B7_o_  (\mux17_oh_b3/or_or_B5_or_B6_B7_o__o , \mux17_oh_b3/B7 , \mux17_oh_b3/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b3/or_or_or_B0_B1_o_or_  (n39[3], \mux17_oh_b3/B2 , \mux17_oh_b3/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b30/and_b0_2  (\mux17_oh_b30/B2 , mtvec_base[30], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b30/and_b0_7  (\mux17_oh_b30/B7 , fres[30], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b30/and_b0_8  (\mux17_oh_b30/B8 , fop1[30], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b30/and_b0_9  (\mux17_oh_b30/B9 , fop2[30], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b30/or_B8_or_B9_B10_o  (\mux17_oh_b30/or_B8_or_B9_B10_o_o , \mux17_oh_b30/B8 , \mux17_oh_b30/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b30/or_or_B5_or_B6_B7_o_  (\mux17_oh_b30/or_or_B5_or_B6_B7_o__o , \mux17_oh_b30/B7 , \mux17_oh_b30/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b30/or_or_or_B0_B1_o_or_  (n39[30], \mux17_oh_b30/B2 , \mux17_oh_b30/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b31/and_b0_2  (\mux17_oh_b31/B2 , mtvec_base[31], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b31/and_b0_7  (\mux17_oh_b31/B7 , fres[31], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b31/and_b0_8  (\mux17_oh_b31/B8 , fop1[31], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b31/and_b0_9  (\mux17_oh_b31/B9 , fop2[31], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b31/or_B8_or_B9_B10_o  (\mux17_oh_b31/or_B8_or_B9_B10_o_o , \mux17_oh_b31/B8 , \mux17_oh_b31/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b31/or_or_B5_or_B6_B7_o_  (\mux17_oh_b31/or_or_B5_or_B6_B7_o__o , \mux17_oh_b31/B7 , \mux17_oh_b31/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b31/or_or_or_B0_B1_o_or_  (n39[31], \mux17_oh_b31/B2 , \mux17_oh_b31/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b4/and_b0_2  (\mux17_oh_b4/B2 , mtvec_base[4], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b4/and_b0_7  (\mux17_oh_b4/B7 , fres[4], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b4/and_b0_8  (\mux17_oh_b4/B8 , fop1[4], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b4/and_b0_9  (\mux17_oh_b4/B9 , fop2[4], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b4/or_B8_or_B9_B10_o  (\mux17_oh_b4/or_B8_or_B9_B10_o_o , \mux17_oh_b4/B8 , \mux17_oh_b4/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b4/or_or_B5_or_B6_B7_o_  (\mux17_oh_b4/or_or_B5_or_B6_B7_o__o , \mux17_oh_b4/B7 , \mux17_oh_b4/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b4/or_or_or_B0_B1_o_or_  (n39[4], \mux17_oh_b4/B2 , \mux17_oh_b4/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b5/and_b0_2  (\mux17_oh_b5/B2 , mtvec_base[5], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b5/and_b0_7  (\mux17_oh_b5/B7 , fres[5], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b5/and_b0_8  (\mux17_oh_b5/B8 , fop1[5], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b5/and_b0_9  (\mux17_oh_b5/B9 , fop2[5], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b5/or_B8_or_B9_B10_o  (\mux17_oh_b5/or_B8_or_B9_B10_o_o , \mux17_oh_b5/B8 , \mux17_oh_b5/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b5/or_or_B5_or_B6_B7_o_  (\mux17_oh_b5/or_or_B5_or_B6_B7_o__o , \mux17_oh_b5/B7 , \mux17_oh_b5/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b5/or_or_or_B0_B1_o_or_  (n39[5], \mux17_oh_b5/B2 , \mux17_oh_b5/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b6/and_b0_2  (\mux17_oh_b6/B2 , mtvec_base[6], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b6/and_b0_7  (\mux17_oh_b6/B7 , fres[6], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b6/and_b0_8  (\mux17_oh_b6/B8 , fop1[6], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b6/and_b0_9  (\mux17_oh_b6/B9 , fop2[6], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b6/or_B8_or_B9_B10_o  (\mux17_oh_b6/or_B8_or_B9_B10_o_o , \mux17_oh_b6/B8 , \mux17_oh_b6/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b6/or_or_B5_or_B6_B7_o_  (\mux17_oh_b6/or_or_B5_or_B6_B7_o__o , \mux17_oh_b6/B7 , \mux17_oh_b6/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b6/or_or_or_B0_B1_o_or_  (n39[6], \mux17_oh_b6/B2 , \mux17_oh_b6/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b7/and_b0_2  (\mux17_oh_b7/B2 , mtvec_base[7], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b7/and_b0_7  (\mux17_oh_b7/B7 , fres[7], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b7/and_b0_8  (\mux17_oh_b7/B8 , fop1[7], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b7/and_b0_9  (\mux17_oh_b7/B9 , fop2[7], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b7/or_B8_or_B9_B10_o  (\mux17_oh_b7/or_B8_or_B9_B10_o_o , \mux17_oh_b7/B8 , \mux17_oh_b7/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b7/or_or_B5_or_B6_B7_o_  (\mux17_oh_b7/or_or_B5_or_B6_B7_o__o , \mux17_oh_b7/B7 , \mux17_oh_b7/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b7/or_or_or_B0_B1_o_or_  (n39[7], \mux17_oh_b7/B2 , \mux17_oh_b7/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b8/and_b0_2  (\mux17_oh_b8/B2 , mtvec_base[8], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b8/and_b0_7  (\mux17_oh_b8/B7 , fres[8], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b8/and_b0_8  (\mux17_oh_b8/B8 , fop1[8], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b8/and_b0_9  (\mux17_oh_b8/B9 , fop2[8], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b8/or_B8_or_B9_B10_o  (\mux17_oh_b8/or_B8_or_B9_B10_o_o , \mux17_oh_b8/B8 , \mux17_oh_b8/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b8/or_or_B5_or_B6_B7_o_  (\mux17_oh_b8/or_or_B5_or_B6_B7_o__o , \mux17_oh_b8/B7 , \mux17_oh_b8/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b8/or_or_or_B0_B1_o_or_  (n39[8], \mux17_oh_b8/B2 , \mux17_oh_b8/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b9/and_b0_2  (\mux17_oh_b9/B2 , mtvec_base[9], n22);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b9/and_b0_7  (\mux17_oh_b9/B7 , fres[9], n27);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b9/and_b0_8  (\mux17_oh_b9/B8 , fop1[9], n28);  // ../RTL/core/csr_regfile.v(170)
  and \mux17_oh_b9/and_b0_9  (\mux17_oh_b9/B9 , fop2[9], n29);  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b9/or_B8_or_B9_B10_o  (\mux17_oh_b9/or_B8_or_B9_B10_o_o , \mux17_oh_b9/B8 , \mux17_oh_b9/B9 );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b9/or_or_B5_or_B6_B7_o_  (\mux17_oh_b9/or_or_B5_or_B6_B7_o__o , \mux17_oh_b9/B7 , \mux17_oh_b9/or_B8_or_B9_B10_o_o );  // ../RTL/core/csr_regfile.v(170)
  or \mux17_oh_b9/or_or_or_B0_B1_o_or_  (n39[9], \mux17_oh_b9/B2 , \mux17_oh_b9/or_or_B5_or_B6_B7_o__o );  // ../RTL/core/csr_regfile.v(170)
  binary_mux_s1_w1 mux18_b0 (
    .i0(n39[0]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[0]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b1 (
    .i0(n39[1]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[1]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b10 (
    .i0(n39[10]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[10]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b11 (
    .i0(n39[11]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[11]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b12 (
    .i0(n39[12]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[12]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b13 (
    .i0(n39[13]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[13]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b14 (
    .i0(n39[14]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[14]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b15 (
    .i0(n39[15]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[15]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b16 (
    .i0(n39[16]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[16]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b17 (
    .i0(n39[17]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[17]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b18 (
    .i0(n39[18]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[18]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b19 (
    .i0(n39[19]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[19]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b2 (
    .i0(n39[2]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[2]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b20 (
    .i0(n39[20]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[20]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b21 (
    .i0(n39[21]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[21]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b22 (
    .i0(n39[22]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[22]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b23 (
    .i0(n39[23]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[23]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b24 (
    .i0(n39[24]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[24]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b25 (
    .i0(n39[25]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[25]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b26 (
    .i0(n39[26]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[26]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b27 (
    .i0(n39[27]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[27]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b28 (
    .i0(n39[28]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[28]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b29 (
    .i0(n39[29]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[29]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b3 (
    .i0(n39[3]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[3]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b30 (
    .i0(n39[30]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[30]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b31 (
    .i0(n39[31]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[31]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b4 (
    .i0(n39[4]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[4]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b5 (
    .i0(n39[5]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[5]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b6 (
    .i0(n39[6]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[6]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b7 (
    .i0(n39[7]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[7]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b8 (
    .i0(n39[8]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[8]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s1_w1 mux18_b9 (
    .i0(n39[9]),
    .i1(1'b0),
    .sel(n19),
    .o(o_csr_rdata[9]));  // ../RTL/core/csr_regfile.v(169)
  binary_mux_s2_w1 mux4_oh_b0 (
    .i0(fres0_add[0]),
    .i1(fres0_sub[0]),
    .i2(fres0_mul[0]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[0]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b1 (
    .i0(fres0_add[1]),
    .i1(fres0_sub[1]),
    .i2(fres0_mul[1]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[1]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b10 (
    .i0(fres0_add[10]),
    .i1(fres0_sub[10]),
    .i2(fres0_mul[10]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[10]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b11 (
    .i0(fres0_add[11]),
    .i1(fres0_sub[11]),
    .i2(fres0_mul[11]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[11]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b12 (
    .i0(fres0_add[12]),
    .i1(fres0_sub[12]),
    .i2(fres0_mul[12]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[12]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b13 (
    .i0(fres0_add[13]),
    .i1(fres0_sub[13]),
    .i2(fres0_mul[13]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[13]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b14 (
    .i0(fres0_add[14]),
    .i1(fres0_sub[14]),
    .i2(fres0_mul[14]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[14]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b15 (
    .i0(fres0_add[15]),
    .i1(fres0_sub[15]),
    .i2(fres0_mul[15]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[15]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b16 (
    .i0(fres0_add[16]),
    .i1(fres0_sub[16]),
    .i2(fres0_mul[16]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[16]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b17 (
    .i0(fres0_add[17]),
    .i1(fres0_sub[17]),
    .i2(fres0_mul[17]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[17]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b18 (
    .i0(fres0_add[18]),
    .i1(fres0_sub[18]),
    .i2(fres0_mul[18]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[18]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b19 (
    .i0(fres0_add[19]),
    .i1(fres0_sub[19]),
    .i2(fres0_mul[19]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[19]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b2 (
    .i0(fres0_add[2]),
    .i1(fres0_sub[2]),
    .i2(fres0_mul[2]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[2]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b20 (
    .i0(fres0_add[20]),
    .i1(fres0_sub[20]),
    .i2(fres0_mul[20]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[20]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b21 (
    .i0(fres0_add[21]),
    .i1(fres0_sub[21]),
    .i2(fres0_mul[21]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[21]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b22 (
    .i0(fres0_add[22]),
    .i1(fres0_sub[22]),
    .i2(fres0_mul[22]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[22]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b23 (
    .i0(fres0_add[23]),
    .i1(fres0_sub[23]),
    .i2(fres0_mul[23]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[23]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b24 (
    .i0(fres0_add[24]),
    .i1(fres0_sub[24]),
    .i2(fres0_mul[24]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[24]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b25 (
    .i0(fres0_add[25]),
    .i1(fres0_sub[25]),
    .i2(fres0_mul[25]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[25]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b26 (
    .i0(fres0_add[26]),
    .i1(fres0_sub[26]),
    .i2(fres0_mul[26]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[26]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b27 (
    .i0(fres0_add[27]),
    .i1(fres0_sub[27]),
    .i2(fres0_mul[27]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[27]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b28 (
    .i0(fres0_add[28]),
    .i1(fres0_sub[28]),
    .i2(fres0_mul[28]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[28]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b29 (
    .i0(fres0_add[29]),
    .i1(fres0_sub[29]),
    .i2(fres0_mul[29]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[29]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b3 (
    .i0(fres0_add[3]),
    .i1(fres0_sub[3]),
    .i2(fres0_mul[3]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[3]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b30 (
    .i0(fres0_add[30]),
    .i1(fres0_sub[30]),
    .i2(fres0_mul[30]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[30]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b31 (
    .i0(fres0_add[31]),
    .i1(fres0_sub[31]),
    .i2(fres0_mul[31]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[31]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b4 (
    .i0(fres0_add[4]),
    .i1(fres0_sub[4]),
    .i2(fres0_mul[4]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[4]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b5 (
    .i0(fres0_add[5]),
    .i1(fres0_sub[5]),
    .i2(fres0_mul[5]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[5]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b6 (
    .i0(fres0_add[6]),
    .i1(fres0_sub[6]),
    .i2(fres0_mul[6]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[6]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b7 (
    .i0(fres0_add[7]),
    .i1(fres0_sub[7]),
    .i2(fres0_mul[7]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[7]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b8 (
    .i0(fres0_add[8]),
    .i1(fres0_sub[8]),
    .i2(fres0_mul[8]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[8]));  // ../RTL/core/csr_regfile.v(134)
  binary_mux_s2_w1 mux4_oh_b9 (
    .i0(fres0_add[9]),
    .i1(fres0_sub[9]),
    .i2(fres0_mul[9]),
    .i3(1'b0),
    .sel(fctrl[1:0]),
    .o(fres[9]));  // ../RTL/core/csr_regfile.v(134)
  AL_DFF_0 reg0_b0 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[0]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_mode[0]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg0_b1 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[1]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_mode[1]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_X reg1_b0 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[0]),
    .en(n11),
    .sr(1'b0),
    .ss(1'b0),
    .q(fctrl[0]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg1_b1 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[1]),
    .en(n11),
    .sr(1'b0),
    .ss(1'b0),
    .q(fctrl[1]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b0 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[0]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[0]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b1 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[1]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[1]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b10 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[10]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[10]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b11 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[11]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[11]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b12 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[12]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[12]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b13 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[13]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[13]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b14 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[14]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[14]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b15 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[15]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[15]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b16 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[16]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[16]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b17 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[17]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[17]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b18 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[18]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[18]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b19 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[19]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[19]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b2 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[2]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[2]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b20 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[20]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[20]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b21 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[21]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[21]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b22 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[22]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[22]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b23 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[23]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[23]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b24 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[24]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[24]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b25 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[25]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[25]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b26 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[26]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[26]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b27 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[27]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[27]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b28 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[28]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[28]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b29 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[29]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[29]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b3 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[3]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[3]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b30 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[30]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[30]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b31 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[31]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[31]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b4 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[4]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[4]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b5 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[5]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[5]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b6 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[6]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[6]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b7 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[7]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[7]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b8 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[8]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[8]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg2_b9 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[9]),
    .en(n14),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop1[9]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b0 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[0]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[0]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b1 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[1]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[1]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b10 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[10]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[10]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b11 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[11]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[11]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b12 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[12]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[12]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b13 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[13]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[13]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b14 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[14]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[14]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b15 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[15]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[15]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b16 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[16]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[16]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b17 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[17]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[17]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b18 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[18]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[18]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b19 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[19]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[19]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b2 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[2]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[2]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b20 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[20]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[20]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b21 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[21]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[21]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b22 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[22]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[22]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b23 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[23]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[23]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b24 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[24]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[24]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b25 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[25]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[25]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b26 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[26]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[26]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b27 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[27]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[27]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b28 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[28]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[28]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b29 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[29]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[29]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b3 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[3]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[3]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b30 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[30]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[30]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b31 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[31]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[31]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b4 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[4]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[4]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b5 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[5]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[5]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b6 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[6]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[6]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b7 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[7]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[7]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b8 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[8]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[8]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_X reg3_b9 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[9]),
    .en(n17),
    .sr(1'b0),
    .ss(1'b0),
    .q(fop2[9]));  // ../RTL/core/csr_regfile.v(139)
  AL_DFF_0 reg4_b0 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[2]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[2]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b1 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[3]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[3]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b10 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[12]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[12]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b11 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[13]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[13]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b12 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[14]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[14]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b13 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[15]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[15]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b14 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[16]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[16]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b15 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[17]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[17]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b16 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[18]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[18]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b17 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[19]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[19]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b18 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[20]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[20]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b19 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[21]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[21]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b2 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[4]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[4]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b20 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[22]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[22]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b21 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[23]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[23]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b22 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[24]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[24]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b23 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[25]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[25]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b24 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[26]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[26]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b25 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[27]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[27]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b26 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[28]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[28]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b27 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[29]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[29]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b28 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[30]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[30]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b29 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[31]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[31]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b3 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[5]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[5]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b4 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[6]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[6]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b5 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[7]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[7]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b6 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[8]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[8]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b7 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[9]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[9]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b8 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[10]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[10]));  // ../RTL/core/csr_regfile.v(64)
  AL_DFF_0 reg4_b9 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(i_csr_wdata[11]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mtvec_base[11]));  // ../RTL/core/csr_regfile.v(64)
  and u13 (n11, i_csr_wen, n10);  // ../RTL/core/csr_regfile.v(144)
  and u14 (n14, i_csr_wen, n13);  // ../RTL/core/csr_regfile.v(147)
  and u15 (n17, i_csr_wen, n16);  // ../RTL/core/csr_regfile.v(150)
  not u17 (n19, i_csr_ren);  // ../RTL/core/csr_regfile.v(169)
  and u9 (n1, i_csr_wen, n0);  // ../RTL/core/csr_regfile.v(68)
  FPU32 u_FPU1 (
    .i_clk(i_clk),
    .i_op1(fop1),
    .i_op2(fop2),
    .i_rsn(1'b0),
    .o_addres(fres0_add),
    .o_mulres(fres0_mul),
    .o_subres(fres0_sub));  // ../RTL/core/csr_regfile.v(157)

endmodule 

module EXU  // ../RTL/core/exu.v(14)
  (
  i_clk,
  i_csr_rdata,
  i_csr_zimm,
  i_csridx,
  i_decinfo,
  i_decinfo_grp,
  i_exu_op1,
  i_exu_op2,
  i_iaddr,
  i_imm,
  i_rdidx,
  i_rdwen,
  i_ribm_gnt,
  i_ribm_rdata,
  i_ribm_rsp,
  i_rs2rdata,
  i_rstn,
  i_vld,
  o_csr_wdata,
  o_csr_wen,
  o_csridx,
  o_exu_jaddr,
  o_exu_rdidx0,
  o_exu_rdidx1,
  o_exu_rdidx2,
  o_exu_rdwen0,
  o_exu_rdwen1,
  o_exu_rdwen2,
  o_exu_resource_match,
  o_exu_taken,
  o_lsu_working,
  o_mdu_working,
  o_rdidx0,
  o_rdidx1,
  o_rdidx2,
  o_rdwdata0,
  o_rdwdata1,
  o_rdwdata2,
  o_rdwen0,
  o_rdwen1,
  o_rdwen2,
  o_ribm_addr,
  o_ribm_mask,
  o_ribm_rdy,
  o_ribm_req,
  o_ribm_wdata,
  o_ribm_wrcs
  );

  input i_clk;  // ../RTL/core/exu.v(15)
  input [31:0] i_csr_rdata;  // ../RTL/core/exu.v(29)
  input [31:0] i_csr_zimm;  // ../RTL/core/exu.v(30)
  input [11:0] i_csridx;  // ../RTL/core/exu.v(28)
  input [9:0] i_decinfo;  // ../RTL/core/exu.v(33)
  input [5:0] i_decinfo_grp;  // ../RTL/core/exu.v(32)
  input [31:0] i_exu_op1;  // ../RTL/core/exu.v(21)
  input [31:0] i_exu_op2;  // ../RTL/core/exu.v(22)
  input [31:0] i_iaddr;  // ../RTL/core/exu.v(34)
  input [31:0] i_imm;  // ../RTL/core/exu.v(24)
  input [4:0] i_rdidx;  // ../RTL/core/exu.v(26)
  input i_rdwen;  // ../RTL/core/exu.v(25)
  input i_ribm_gnt;  // ../RTL/core/exu.v(76)
  input [31:0] i_ribm_rdata;  // ../RTL/core/exu.v(74)
  input i_ribm_rsp;  // ../RTL/core/exu.v(77)
  input [31:0] i_rs2rdata;  // ../RTL/core/exu.v(23)
  input i_rstn;  // ../RTL/core/exu.v(16)
  input i_vld;  // ../RTL/core/exu.v(18)
  output [31:0] o_csr_wdata;  // ../RTL/core/exu.v(62)
  output o_csr_wen;  // ../RTL/core/exu.v(60)
  output [11:0] o_csridx;  // ../RTL/core/exu.v(61)
  output [31:0] o_exu_jaddr;  // ../RTL/core/exu.v(66)
  output [4:0] o_exu_rdidx0;  // ../RTL/core/exu.v(39)
  output [4:0] o_exu_rdidx1;  // ../RTL/core/exu.v(41)
  output [4:0] o_exu_rdidx2;  // ../RTL/core/exu.v(43)
  output o_exu_rdwen0;  // ../RTL/core/exu.v(38)
  output o_exu_rdwen1;  // ../RTL/core/exu.v(40)
  output o_exu_rdwen2;  // ../RTL/core/exu.v(42)
  output o_exu_resource_match;  // ../RTL/core/exu.v(44)
  output o_exu_taken;  // ../RTL/core/exu.v(65)
  output o_lsu_working;  // ../RTL/core/exu.v(55)
  output o_mdu_working;  // ../RTL/core/exu.v(51)
  output [4:0] o_rdidx0;  // ../RTL/core/exu.v(49)
  output [4:0] o_rdidx1;  // ../RTL/core/exu.v(53)
  output [4:0] o_rdidx2;  // ../RTL/core/exu.v(57)
  output [31:0] o_rdwdata0;  // ../RTL/core/exu.v(50)
  output [31:0] o_rdwdata1;  // ../RTL/core/exu.v(54)
  output [31:0] o_rdwdata2;  // ../RTL/core/exu.v(58)
  output o_rdwen0;  // ../RTL/core/exu.v(48)
  output o_rdwen1;  // ../RTL/core/exu.v(52)
  output o_rdwen2;  // ../RTL/core/exu.v(56)
  output [31:0] o_ribm_addr;  // ../RTL/core/exu.v(70)
  output [3:0] o_ribm_mask;  // ../RTL/core/exu.v(72)
  output o_ribm_rdy;  // ../RTL/core/exu.v(78)
  output o_ribm_req;  // ../RTL/core/exu.v(75)
  output [31:0] o_ribm_wdata;  // ../RTL/core/exu.v(73)
  output o_ribm_wrcs;  // ../RTL/core/exu.v(71)

  wire [31:0] alu2lsu_result;  // ../RTL/core/exu.v(90)
  wire [31:0] alu_rdwdata;  // ../RTL/core/exu.v(89)
  wire [31:0] bju_rdwdata;  // ../RTL/core/exu.v(109)
  wire [31:0] n2;
  wire [31:0] n3;
  wire [31:0] \u_EXU_ALU/alu_and ;  // ../RTL/core/exu_alu.v(51)
  wire [31:0] \u_EXU_ALU/alu_or ;  // ../RTL/core/exu_alu.v(53)
  wire [31:0] \u_EXU_ALU/alu_sll ;  // ../RTL/core/exu_alu.v(43)
  wire [31:0] \u_EXU_ALU/alu_slt ;  // ../RTL/core/exu_alu.v(55)
  wire [31:0] \u_EXU_ALU/alu_sltu ;  // ../RTL/core/exu_alu.v(57)
  wire [31:0] \u_EXU_ALU/alu_sra ;  // ../RTL/core/exu_alu.v(47)
  wire [31:0] \u_EXU_ALU/alu_srl ;  // ../RTL/core/exu_alu.v(45)
  wire [31:0] \u_EXU_ALU/alu_sub ;  // ../RTL/core/exu_alu.v(41)
  wire [31:0] \u_EXU_ALU/alu_xor ;  // ../RTL/core/exu_alu.v(49)
  wire [31:0] \u_EXU_ALU/n0 ;
  wire [31:0] \u_EXU_ALU/n132 ;
  wire [31:0] \u_EXU_ALU/n133 ;
  wire [31:0] \u_EXU_ALU/n135 ;
  wire [31:0] \u_EXU_ALU/n168 ;
  wire [31:0] \u_EXU_ALU/n201 ;
  wire [31:0] \u_EXU_ALU/n233 ;
  wire [31:0] \u_EXU_ALU/n303 ;
  wire [31:0] \u_EXU_ALU/n304 ;
  wire [31:0] \u_EXU_ALU/n305 ;
  wire [31:0] \u_EXU_ALU/n306 ;
  wire [31:0] \u_EXU_ALU/n307 ;
  wire [31:0] \u_EXU_ALU/n308 ;
  wire [31:0] \u_EXU_ALU/n309 ;
  wire [31:0] \u_EXU_ALU/n310 ;
  wire [31:0] \u_EXU_ALU/n33 ;
  wire [31:0] \u_EXU_ALU/n66 ;
  wire [31:0] \u_EXU_ALU/n99 ;
  wire [31:0] \u_EXU_BJU/bxx_nxtpc ;  // ../RTL/core/exu_bju.v(57)
  wire [63:0] \u_EXU_LSU/access2_data ;  // ../RTL/core/exu_lsu.v(209)
  wire [31:0] \u_EXU_LSU/access_data ;  // ../RTL/core/exu_lsu.v(210)
  wire [1:0] \u_EXU_LSU/align_mode_reg ;  // ../RTL/core/exu_lsu.v(98)
  wire [9:0] \u_EXU_LSU/lsuinfo ;  // ../RTL/core/exu_lsu.v(94)
  wire [31:0] \u_EXU_LSU/n136 ;
  wire [31:0] \u_EXU_LSU/n137 ;
  wire [15:0] \u_EXU_LSU/n138 ;
  wire [23:0] \u_EXU_LSU/n139 ;
  wire [31:0] \u_EXU_LSU/n140 ;
  wire [31:0] \u_EXU_LSU/n141 ;
  wire [31:0] \u_EXU_LSU/n49 ;
  wire [31:0] \u_EXU_LSU/n50 ;
  wire [31:0] \u_EXU_LSU/n52 ;
  wire [31:0] \u_EXU_LSU/n53 ;
  wire [31:0] \u_EXU_LSU/n54 ;
  wire [31:0] \u_EXU_LSU/n55 ;
  wire [29:0] \u_EXU_LSU/n59 ;
  wire [3:0] \u_EXU_LSU/n60 ;
  wire [3:0] \u_EXU_LSU/n61 ;
  wire [3:0] \u_EXU_LSU/n62 ;
  wire [3:0] \u_EXU_LSU/n63 ;
  wire [3:0] \u_EXU_LSU/n64 ;
  wire [3:0] \u_EXU_LSU/n65 ;
  wire [3:0] \u_EXU_LSU/n66 ;
  wire [31:0] \u_EXU_LSU/n67 ;
  wire [31:0] \u_EXU_LSU/n72 ;
  wire [3:0] \u_EXU_LSU/n73 ;
  wire [31:0] \u_EXU_LSU/n74 ;
  wire [31:0] \u_EXU_LSU/n76 ;
  wire [3:0] \u_EXU_LSU/n78 ;
  wire [31:0] \u_EXU_LSU/n79 ;
  wire [31:0] \u_EXU_LSU/overleft_buffer ;  // ../RTL/core/exu_lsu.v(100)
  wire [31:0] \u_EXU_LSU/rs2rdata_reg ;  // ../RTL/core/exu_lsu.v(99)
  wire [31:0] \u_EXU_SCU/csr_rc ;  // ../RTL/core/exu_scu.v(49)
  wire [31:0] \u_EXU_SCU/csr_rs ;  // ../RTL/core/exu_scu.v(48)
  wire [31:0] \u_EXU_SCU/csr_rw ;  // ../RTL/core/exu_scu.v(47)
  wire [31:0] \u_EXU_SCU/n0 ;
  wire [31:0] \u_EXU_SCU/n1 ;
  wire [31:0] \u_EXU_SCU/n2 ;
  wire [31:0] \u_EXU_SCU/n3 ;
  wire [31:0] \u_EXU_SCU/n4 ;
  wire \alu2lsu_result[1]_neg ;
  wire bju_rdwen;  // ../RTL/core/exu.v(108)
  wire \i_decinfo[2]_neg ;
  wire \i_decinfo[3]_neg ;
  wire \i_decinfo[4]_neg ;
  wire \i_exu_op2[4]_neg ;
  wire lsu_flush;  // ../RTL/core/exu.v(209)
  wire mdu_flush;  // ../RTL/core/exu.v(172)
  wire n0;
  wire n1;
  wire n4;
  wire n5;
  wire n6;
  wire n7;
  wire n8;
  wire n9;
  wire \u_EXU_ALU/n100 ;
  wire \u_EXU_ALU/n101 ;
  wire \u_EXU_ALU/n102 ;
  wire \u_EXU_ALU/n103 ;
  wire \u_EXU_ALU/n104 ;
  wire \u_EXU_ALU/n105 ;
  wire \u_EXU_ALU/n106 ;
  wire \u_EXU_ALU/n107 ;
  wire \u_EXU_ALU/n108 ;
  wire \u_EXU_ALU/n109 ;
  wire \u_EXU_ALU/n110 ;
  wire \u_EXU_ALU/n111 ;
  wire \u_EXU_ALU/n112 ;
  wire \u_EXU_ALU/n113 ;
  wire \u_EXU_ALU/n114 ;
  wire \u_EXU_ALU/n115 ;
  wire \u_EXU_ALU/n116 ;
  wire \u_EXU_ALU/n117 ;
  wire \u_EXU_ALU/n118 ;
  wire \u_EXU_ALU/n119 ;
  wire \u_EXU_ALU/n120 ;
  wire \u_EXU_ALU/n121 ;
  wire \u_EXU_ALU/n122 ;
  wire \u_EXU_ALU/n123 ;
  wire \u_EXU_ALU/n124 ;
  wire \u_EXU_ALU/n125 ;
  wire \u_EXU_ALU/n126 ;
  wire \u_EXU_ALU/n127 ;
  wire \u_EXU_ALU/n128 ;
  wire \u_EXU_ALU/n129 ;
  wire \u_EXU_ALU/n130 ;
  wire \u_EXU_ALU/n131 ;
  wire \u_EXU_ALU/n134 ;
  wire \u_EXU_ALU/n136 ;
  wire \u_EXU_ALU/n137 ;
  wire \u_EXU_ALU/n138 ;
  wire \u_EXU_ALU/n139 ;
  wire \u_EXU_ALU/n140 ;
  wire \u_EXU_ALU/n141 ;
  wire \u_EXU_ALU/n142 ;
  wire \u_EXU_ALU/n143 ;
  wire \u_EXU_ALU/n144 ;
  wire \u_EXU_ALU/n145 ;
  wire \u_EXU_ALU/n146 ;
  wire \u_EXU_ALU/n147 ;
  wire \u_EXU_ALU/n148 ;
  wire \u_EXU_ALU/n149 ;
  wire \u_EXU_ALU/n150 ;
  wire \u_EXU_ALU/n151 ;
  wire \u_EXU_ALU/n152 ;
  wire \u_EXU_ALU/n153 ;
  wire \u_EXU_ALU/n154 ;
  wire \u_EXU_ALU/n155 ;
  wire \u_EXU_ALU/n156 ;
  wire \u_EXU_ALU/n157 ;
  wire \u_EXU_ALU/n158 ;
  wire \u_EXU_ALU/n159 ;
  wire \u_EXU_ALU/n160 ;
  wire \u_EXU_ALU/n161 ;
  wire \u_EXU_ALU/n162 ;
  wire \u_EXU_ALU/n163 ;
  wire \u_EXU_ALU/n164 ;
  wire \u_EXU_ALU/n165 ;
  wire \u_EXU_ALU/n166 ;
  wire \u_EXU_ALU/n167 ;
  wire \u_EXU_ALU/n169 ;
  wire \u_EXU_ALU/n170 ;
  wire \u_EXU_ALU/n171 ;
  wire \u_EXU_ALU/n172 ;
  wire \u_EXU_ALU/n173 ;
  wire \u_EXU_ALU/n174 ;
  wire \u_EXU_ALU/n175 ;
  wire \u_EXU_ALU/n176 ;
  wire \u_EXU_ALU/n177 ;
  wire \u_EXU_ALU/n178 ;
  wire \u_EXU_ALU/n179 ;
  wire \u_EXU_ALU/n179_neg ;
  wire \u_EXU_ALU/n180 ;
  wire \u_EXU_ALU/n181 ;
  wire \u_EXU_ALU/n182 ;
  wire \u_EXU_ALU/n183 ;
  wire \u_EXU_ALU/n184 ;
  wire \u_EXU_ALU/n185 ;
  wire \u_EXU_ALU/n186 ;
  wire \u_EXU_ALU/n187 ;
  wire \u_EXU_ALU/n188 ;
  wire \u_EXU_ALU/n189 ;
  wire \u_EXU_ALU/n190 ;
  wire \u_EXU_ALU/n191 ;
  wire \u_EXU_ALU/n192 ;
  wire \u_EXU_ALU/n193 ;
  wire \u_EXU_ALU/n194 ;
  wire \u_EXU_ALU/n195 ;
  wire \u_EXU_ALU/n196 ;
  wire \u_EXU_ALU/n197 ;
  wire \u_EXU_ALU/n198 ;
  wire \u_EXU_ALU/n199 ;
  wire \u_EXU_ALU/n200 ;
  wire \u_EXU_ALU/n202 ;
  wire \u_EXU_ALU/n203 ;
  wire \u_EXU_ALU/n204 ;
  wire \u_EXU_ALU/n205 ;
  wire \u_EXU_ALU/n222 ;
  wire \u_EXU_ALU/n223 ;
  wire \u_EXU_ALU/n224 ;
  wire \u_EXU_ALU/n225 ;
  wire \u_EXU_ALU/n226 ;
  wire \u_EXU_ALU/n227 ;
  wire \u_EXU_ALU/n228 ;
  wire \u_EXU_ALU/n229 ;
  wire \u_EXU_ALU/n230 ;
  wire \u_EXU_ALU/n231 ;
  wire \u_EXU_ALU/n232 ;
  wire \u_EXU_ALU/n234 ;
  wire \u_EXU_ALU/n235 ;
  wire \u_EXU_ALU/n236 ;
  wire \u_EXU_ALU/n237 ;
  wire \u_EXU_ALU/n238 ;
  wire \u_EXU_ALU/n239 ;
  wire \u_EXU_ALU/n240 ;
  wire \u_EXU_ALU/n241 ;
  wire \u_EXU_ALU/n242 ;
  wire \u_EXU_ALU/n243 ;
  wire \u_EXU_ALU/n244 ;
  wire \u_EXU_ALU/n245 ;
  wire \u_EXU_ALU/n246 ;
  wire \u_EXU_ALU/n247 ;
  wire \u_EXU_ALU/n248 ;
  wire \u_EXU_ALU/n249 ;
  wire \u_EXU_ALU/n250 ;
  wire \u_EXU_ALU/n251 ;
  wire \u_EXU_ALU/n252 ;
  wire \u_EXU_ALU/n253 ;
  wire \u_EXU_ALU/n254 ;
  wire \u_EXU_ALU/n255 ;
  wire \u_EXU_ALU/n256 ;
  wire \u_EXU_ALU/n257 ;
  wire \u_EXU_ALU/n258 ;
  wire \u_EXU_ALU/n259 ;
  wire \u_EXU_ALU/n260 ;
  wire \u_EXU_ALU/n261 ;
  wire \u_EXU_ALU/n262 ;
  wire \u_EXU_ALU/n263 ;
  wire \u_EXU_ALU/n264 ;
  wire \u_EXU_ALU/n265 ;
  wire \u_EXU_ALU/n266 ;
  wire \u_EXU_ALU/n267 ;
  wire \u_EXU_ALU/n268 ;
  wire \u_EXU_ALU/n269 ;
  wire \u_EXU_ALU/n27 ;
  wire \u_EXU_ALU/n270 ;
  wire \u_EXU_ALU/n271 ;
  wire \u_EXU_ALU/n272 ;
  wire \u_EXU_ALU/n273 ;
  wire \u_EXU_ALU/n274 ;
  wire \u_EXU_ALU/n275 ;
  wire \u_EXU_ALU/n276 ;
  wire \u_EXU_ALU/n277 ;
  wire \u_EXU_ALU/n278 ;
  wire \u_EXU_ALU/n279 ;
  wire \u_EXU_ALU/n28 ;
  wire \u_EXU_ALU/n280 ;
  wire \u_EXU_ALU/n281 ;
  wire \u_EXU_ALU/n281_neg ;
  wire \u_EXU_ALU/n282 ;
  wire \u_EXU_ALU/n283 ;
  wire \u_EXU_ALU/n284 ;
  wire \u_EXU_ALU/n285 ;
  wire \u_EXU_ALU/n286 ;
  wire \u_EXU_ALU/n287 ;
  wire \u_EXU_ALU/n288 ;
  wire \u_EXU_ALU/n289 ;
  wire \u_EXU_ALU/n29 ;
  wire \u_EXU_ALU/n290 ;
  wire \u_EXU_ALU/n291 ;
  wire \u_EXU_ALU/n292 ;
  wire \u_EXU_ALU/n293 ;
  wire \u_EXU_ALU/n297 ;
  wire \u_EXU_ALU/n298 ;
  wire \u_EXU_ALU/n299 ;
  wire \u_EXU_ALU/n30 ;
  wire \u_EXU_ALU/n300 ;
  wire \u_EXU_ALU/n301 ;
  wire \u_EXU_ALU/n302 ;
  wire \u_EXU_ALU/n31 ;
  wire \u_EXU_ALU/n311 ;
  wire \u_EXU_ALU/n312 ;
  wire \u_EXU_ALU/n313 ;
  wire \u_EXU_ALU/n314 ;
  wire \u_EXU_ALU/n315 ;
  wire \u_EXU_ALU/n316 ;
  wire \u_EXU_ALU/n317 ;
  wire \u_EXU_ALU/n318 ;
  wire \u_EXU_ALU/n319 ;
  wire \u_EXU_ALU/n32 ;
  wire \u_EXU_ALU/n320 ;
  wire \u_EXU_ALU/n321 ;
  wire \u_EXU_ALU/n322 ;
  wire \u_EXU_ALU/n323 ;
  wire \u_EXU_ALU/n324 ;
  wire \u_EXU_ALU/n325 ;
  wire \u_EXU_ALU/n326 ;
  wire \u_EXU_ALU/n327 ;
  wire \u_EXU_ALU/n328 ;
  wire \u_EXU_ALU/n329 ;
  wire \u_EXU_ALU/n330 ;
  wire \u_EXU_ALU/n331 ;
  wire \u_EXU_ALU/n332 ;
  wire \u_EXU_ALU/n333 ;
  wire \u_EXU_ALU/n334 ;
  wire \u_EXU_ALU/n335 ;
  wire \u_EXU_ALU/n336 ;
  wire \u_EXU_ALU/n337 ;
  wire \u_EXU_ALU/n338 ;
  wire \u_EXU_ALU/n339 ;
  wire \u_EXU_ALU/n34 ;
  wire \u_EXU_ALU/n340 ;
  wire \u_EXU_ALU/n341 ;
  wire \u_EXU_ALU/n342 ;
  wire \u_EXU_ALU/n343 ;
  wire \u_EXU_ALU/n344 ;
  wire \u_EXU_ALU/n345 ;
  wire \u_EXU_ALU/n346 ;
  wire \u_EXU_ALU/n347 ;
  wire \u_EXU_ALU/n348 ;
  wire \u_EXU_ALU/n349 ;
  wire \u_EXU_ALU/n35 ;
  wire \u_EXU_ALU/n350 ;
  wire \u_EXU_ALU/n351 ;
  wire \u_EXU_ALU/n352 ;
  wire \u_EXU_ALU/n353 ;
  wire \u_EXU_ALU/n354 ;
  wire \u_EXU_ALU/n355 ;
  wire \u_EXU_ALU/n356 ;
  wire \u_EXU_ALU/n357 ;
  wire \u_EXU_ALU/n358 ;
  wire \u_EXU_ALU/n359 ;
  wire \u_EXU_ALU/n36 ;
  wire \u_EXU_ALU/n360 ;
  wire \u_EXU_ALU/n361 ;
  wire \u_EXU_ALU/n362 ;
  wire \u_EXU_ALU/n363 ;
  wire \u_EXU_ALU/n364 ;
  wire \u_EXU_ALU/n365 ;
  wire \u_EXU_ALU/n366 ;
  wire \u_EXU_ALU/n367 ;
  wire \u_EXU_ALU/n368 ;
  wire \u_EXU_ALU/n369 ;
  wire \u_EXU_ALU/n37 ;
  wire \u_EXU_ALU/n370 ;
  wire \u_EXU_ALU/n371 ;
  wire \u_EXU_ALU/n372 ;
  wire \u_EXU_ALU/n373 ;
  wire \u_EXU_ALU/n374 ;
  wire \u_EXU_ALU/n375 ;
  wire \u_EXU_ALU/n376 ;
  wire \u_EXU_ALU/n377 ;
  wire \u_EXU_ALU/n378 ;
  wire \u_EXU_ALU/n379 ;
  wire \u_EXU_ALU/n38 ;
  wire \u_EXU_ALU/n380 ;
  wire \u_EXU_ALU/n381 ;
  wire \u_EXU_ALU/n382 ;
  wire \u_EXU_ALU/n383 ;
  wire \u_EXU_ALU/n384 ;
  wire \u_EXU_ALU/n385 ;
  wire \u_EXU_ALU/n386 ;
  wire \u_EXU_ALU/n387 ;
  wire \u_EXU_ALU/n388 ;
  wire \u_EXU_ALU/n389 ;
  wire \u_EXU_ALU/n39 ;
  wire \u_EXU_ALU/n390 ;
  wire \u_EXU_ALU/n391 ;
  wire \u_EXU_ALU/n392 ;
  wire \u_EXU_ALU/n393 ;
  wire \u_EXU_ALU/n394 ;
  wire \u_EXU_ALU/n395 ;
  wire \u_EXU_ALU/n396 ;
  wire \u_EXU_ALU/n397 ;
  wire \u_EXU_ALU/n398 ;
  wire \u_EXU_ALU/n399 ;
  wire \u_EXU_ALU/n40 ;
  wire \u_EXU_ALU/n400 ;
  wire \u_EXU_ALU/n401 ;
  wire \u_EXU_ALU/n402 ;
  wire \u_EXU_ALU/n403 ;
  wire \u_EXU_ALU/n404 ;
  wire \u_EXU_ALU/n405 ;
  wire \u_EXU_ALU/n406 ;
  wire \u_EXU_ALU/n407 ;
  wire \u_EXU_ALU/n408 ;
  wire \u_EXU_ALU/n409 ;
  wire \u_EXU_ALU/n41 ;
  wire \u_EXU_ALU/n410 ;
  wire \u_EXU_ALU/n411 ;
  wire \u_EXU_ALU/n412 ;
  wire \u_EXU_ALU/n413 ;
  wire \u_EXU_ALU/n414 ;
  wire \u_EXU_ALU/n415 ;
  wire \u_EXU_ALU/n416 ;
  wire \u_EXU_ALU/n417 ;
  wire \u_EXU_ALU/n418 ;
  wire \u_EXU_ALU/n419 ;
  wire \u_EXU_ALU/n42 ;
  wire \u_EXU_ALU/n420 ;
  wire \u_EXU_ALU/n421 ;
  wire \u_EXU_ALU/n422 ;
  wire \u_EXU_ALU/n423 ;
  wire \u_EXU_ALU/n424 ;
  wire \u_EXU_ALU/n425 ;
  wire \u_EXU_ALU/n426 ;
  wire \u_EXU_ALU/n427 ;
  wire \u_EXU_ALU/n428 ;
  wire \u_EXU_ALU/n429 ;
  wire \u_EXU_ALU/n43 ;
  wire \u_EXU_ALU/n430 ;
  wire \u_EXU_ALU/n431 ;
  wire \u_EXU_ALU/n432 ;
  wire \u_EXU_ALU/n44 ;
  wire \u_EXU_ALU/n449 ;
  wire \u_EXU_ALU/n45 ;
  wire \u_EXU_ALU/n450 ;
  wire \u_EXU_ALU/n451 ;
  wire \u_EXU_ALU/n452 ;
  wire \u_EXU_ALU/n453 ;
  wire \u_EXU_ALU/n454 ;
  wire \u_EXU_ALU/n455 ;
  wire \u_EXU_ALU/n456 ;
  wire \u_EXU_ALU/n457 ;
  wire \u_EXU_ALU/n458 ;
  wire \u_EXU_ALU/n459 ;
  wire \u_EXU_ALU/n46 ;
  wire \u_EXU_ALU/n460 ;
  wire \u_EXU_ALU/n461 ;
  wire \u_EXU_ALU/n47 ;
  wire \u_EXU_ALU/n48 ;
  wire \u_EXU_ALU/n49 ;
  wire \u_EXU_ALU/n50 ;
  wire \u_EXU_ALU/n51 ;
  wire \u_EXU_ALU/n52 ;
  wire \u_EXU_ALU/n53 ;
  wire \u_EXU_ALU/n54 ;
  wire \u_EXU_ALU/n55 ;
  wire \u_EXU_ALU/n56 ;
  wire \u_EXU_ALU/n57 ;
  wire \u_EXU_ALU/n58 ;
  wire \u_EXU_ALU/n59 ;
  wire \u_EXU_ALU/n60 ;
  wire \u_EXU_ALU/n61 ;
  wire \u_EXU_ALU/n62 ;
  wire \u_EXU_ALU/n63 ;
  wire \u_EXU_ALU/n64 ;
  wire \u_EXU_ALU/n65 ;
  wire \u_EXU_ALU/n67 ;
  wire \u_EXU_ALU/n68 ;
  wire \u_EXU_ALU/n69 ;
  wire \u_EXU_ALU/n70 ;
  wire \u_EXU_ALU/n71 ;
  wire \u_EXU_ALU/n72 ;
  wire \u_EXU_ALU/n73 ;
  wire \u_EXU_ALU/n74 ;
  wire \u_EXU_ALU/n75 ;
  wire \u_EXU_ALU/n76 ;
  wire \u_EXU_ALU/n77 ;
  wire \u_EXU_ALU/n78 ;
  wire \u_EXU_ALU/n79 ;
  wire \u_EXU_ALU/n80 ;
  wire \u_EXU_ALU/n81 ;
  wire \u_EXU_ALU/n82 ;
  wire \u_EXU_ALU/n83 ;
  wire \u_EXU_ALU/n84 ;
  wire \u_EXU_ALU/n85 ;
  wire \u_EXU_ALU/n86 ;
  wire \u_EXU_ALU/n87 ;
  wire \u_EXU_ALU/n88 ;
  wire \u_EXU_ALU/n89 ;
  wire \u_EXU_ALU/n90 ;
  wire \u_EXU_ALU/n91 ;
  wire \u_EXU_ALU/n92 ;
  wire \u_EXU_ALU/n93 ;
  wire \u_EXU_ALU/n94 ;
  wire \u_EXU_ALU/n95 ;
  wire \u_EXU_ALU/n96 ;
  wire \u_EXU_ALU/n97 ;
  wire \u_EXU_ALU/n98 ;
  wire \u_EXU_ALU/u1029_sel_is_0_o ;
  wire \u_EXU_ALU/u750_sel_is_0_o ;
  wire \u_EXU_BJU/bxx_beq ;  // ../RTL/core/exu_bju.v(42)
  wire \u_EXU_BJU/bxx_bge ;  // ../RTL/core/exu_bju.v(45)
  wire \u_EXU_BJU/bxx_bgeu ;  // ../RTL/core/exu_bju.v(47)
  wire \u_EXU_BJU/bxx_blt ;  // ../RTL/core/exu_bju.v(44)
  wire \u_EXU_BJU/bxx_bltu ;  // ../RTL/core/exu_bju.v(46)
  wire \u_EXU_BJU/bxx_bne ;  // ../RTL/core/exu_bju.v(43)
  wire \u_EXU_BJU/judgeflag ;  // ../RTL/core/exu_bju.v(49)
  wire \u_EXU_BJU/n0 ;
  wire \u_EXU_BJU/n1 ;
  wire \u_EXU_BJU/n10 ;
  wire \u_EXU_BJU/n3 ;
  wire \u_EXU_BJU/n5 ;
  wire \u_EXU_BJU/n6 ;
  wire \u_EXU_BJU/n7 ;
  wire \u_EXU_BJU/n8 ;
  wire \u_EXU_BJU/n9 ;
  wire \u_EXU_LSU/access2_once ;  // ../RTL/core/exu_lsu.v(96)
  wire \u_EXU_LSU/access2_vld ;  // ../RTL/core/exu_lsu.v(95)
  wire \u_EXU_LSU/handshake_once ;  // ../RTL/core/exu_lsu.v(152)
  wire \u_EXU_LSU/handshake_rdy ;  // ../RTL/core/exu_lsu.v(66)
  wire \u_EXU_LSU/handshake_rdy_last ;  // ../RTL/core/exu_lsu.v(69)
  wire \u_EXU_LSU/lsu_finish ;  // ../RTL/core/exu_lsu.v(103)
  wire \u_EXU_LSU/lsu_finish_neg ;
  wire \u_EXU_LSU/lsu_vld ;  // ../RTL/core/exu_lsu.v(101)
  wire \u_EXU_LSU/lsu_vld_neg ;
  wire \u_EXU_LSU/lsuinfo[2]_neg ;
  wire \u_EXU_LSU/lsuinfo[3]_neg ;
  wire \u_EXU_LSU/lsuinfo[4]_neg ;
  wire \u_EXU_LSU/lsuinfo[5]_neg ;
  wire \u_EXU_LSU/mux10_b2_sel_is_2_o ;
  wire \u_EXU_LSU/mux11_b0_sel_is_2_o ;
  wire \u_EXU_LSU/mux12_b1_sel_is_1_o ;
  wire \u_EXU_LSU/mux12_b2_sel_is_3_o ;
  wire \u_EXU_LSU/mux13_b0_sel_is_0_o ;
  wire \u_EXU_LSU/mux14_b0_sel_is_0_o ;
  wire \u_EXU_LSU/mux14_b0_sel_is_2_o ;
  wire \u_EXU_LSU/mux14_b0_sel_is_2_o_neg ;
  wire \u_EXU_LSU/mux14_b1_sel_is_0_o ;
  wire \u_EXU_LSU/mux16_b0_sel_is_0_o ;
  wire \u_EXU_LSU/mux16_b3_sel_is_2_o ;
  wire \u_EXU_LSU/mux1_b0_sel_is_2_o ;
  wire \u_EXU_LSU/mux20_b0_sel_is_0_o ;
  wire \u_EXU_LSU/mux27_b16_sel_is_1_o ;
  wire \u_EXU_LSU/mux32_b0_sel_is_0_o ;
  wire \u_EXU_LSU/mux6_b0_sel_is_2_o ;
  wire \u_EXU_LSU/n0 ;
  wire \u_EXU_LSU/n1 ;
  wire \u_EXU_LSU/n10 ;
  wire \u_EXU_LSU/n100 ;
  wire \u_EXU_LSU/n101 ;
  wire \u_EXU_LSU/n102 ;
  wire \u_EXU_LSU/n11 ;
  wire \u_EXU_LSU/n12 ;
  wire \u_EXU_LSU/n13 ;
  wire \u_EXU_LSU/n13_neg ;
  wire \u_EXU_LSU/n142 ;
  wire \u_EXU_LSU/n143 ;
  wire \u_EXU_LSU/n144 ;
  wire \u_EXU_LSU/n145 ;
  wire \u_EXU_LSU/n146 ;
  wire \u_EXU_LSU/n147 ;
  wire \u_EXU_LSU/n148 ;
  wire \u_EXU_LSU/n149 ;
  wire \u_EXU_LSU/n150 ;
  wire \u_EXU_LSU/n151 ;
  wire \u_EXU_LSU/n152 ;
  wire \u_EXU_LSU/n153 ;
  wire \u_EXU_LSU/n154 ;
  wire \u_EXU_LSU/n155 ;
  wire \u_EXU_LSU/n156 ;
  wire \u_EXU_LSU/n157 ;
  wire \u_EXU_LSU/n158 ;
  wire \u_EXU_LSU/n159 ;
  wire \u_EXU_LSU/n16 ;
  wire \u_EXU_LSU/n160 ;
  wire \u_EXU_LSU/n161 ;
  wire \u_EXU_LSU/n162 ;
  wire \u_EXU_LSU/n163 ;
  wire \u_EXU_LSU/n164 ;
  wire \u_EXU_LSU/n165 ;
  wire \u_EXU_LSU/n166 ;
  wire \u_EXU_LSU/n167 ;
  wire \u_EXU_LSU/n168 ;
  wire \u_EXU_LSU/n169 ;
  wire \u_EXU_LSU/n170 ;
  wire \u_EXU_LSU/n171 ;
  wire \u_EXU_LSU/n172 ;
  wire \u_EXU_LSU/n173 ;
  wire \u_EXU_LSU/n174 ;
  wire \u_EXU_LSU/n175 ;
  wire \u_EXU_LSU/n176 ;
  wire \u_EXU_LSU/n177 ;
  wire \u_EXU_LSU/n178 ;
  wire \u_EXU_LSU/n179 ;
  wire \u_EXU_LSU/n18 ;
  wire \u_EXU_LSU/n180 ;
  wire \u_EXU_LSU/n181 ;
  wire \u_EXU_LSU/n182 ;
  wire \u_EXU_LSU/n183 ;
  wire \u_EXU_LSU/n184 ;
  wire \u_EXU_LSU/n185 ;
  wire \u_EXU_LSU/n186 ;
  wire \u_EXU_LSU/n187 ;
  wire \u_EXU_LSU/n188 ;
  wire \u_EXU_LSU/n189 ;
  wire \u_EXU_LSU/n19 ;
  wire \u_EXU_LSU/n190 ;
  wire \u_EXU_LSU/n191 ;
  wire \u_EXU_LSU/n192 ;
  wire \u_EXU_LSU/n193 ;
  wire \u_EXU_LSU/n194 ;
  wire \u_EXU_LSU/n195 ;
  wire \u_EXU_LSU/n196 ;
  wire \u_EXU_LSU/n197 ;
  wire \u_EXU_LSU/n198 ;
  wire \u_EXU_LSU/n199 ;
  wire \u_EXU_LSU/n20 ;
  wire \u_EXU_LSU/n200 ;
  wire \u_EXU_LSU/n201 ;
  wire \u_EXU_LSU/n202 ;
  wire \u_EXU_LSU/n203 ;
  wire \u_EXU_LSU/n204 ;
  wire \u_EXU_LSU/n205 ;
  wire \u_EXU_LSU/n206 ;
  wire \u_EXU_LSU/n207 ;
  wire \u_EXU_LSU/n208 ;
  wire \u_EXU_LSU/n209 ;
  wire \u_EXU_LSU/n210 ;
  wire \u_EXU_LSU/n211 ;
  wire \u_EXU_LSU/n212 ;
  wire \u_EXU_LSU/n213 ;
  wire \u_EXU_LSU/n214 ;
  wire \u_EXU_LSU/n215 ;
  wire \u_EXU_LSU/n216 ;
  wire \u_EXU_LSU/n217 ;
  wire \u_EXU_LSU/n218 ;
  wire \u_EXU_LSU/n219 ;
  wire \u_EXU_LSU/n220 ;
  wire \u_EXU_LSU/n221 ;
  wire \u_EXU_LSU/n222 ;
  wire \u_EXU_LSU/n223 ;
  wire \u_EXU_LSU/n224 ;
  wire \u_EXU_LSU/n225 ;
  wire \u_EXU_LSU/n226 ;
  wire \u_EXU_LSU/n227 ;
  wire \u_EXU_LSU/n228 ;
  wire \u_EXU_LSU/n229 ;
  wire \u_EXU_LSU/n23 ;
  wire \u_EXU_LSU/n25 ;
  wire \u_EXU_LSU/n250 ;
  wire \u_EXU_LSU/n252 ;
  wire \u_EXU_LSU/n253 ;
  wire \u_EXU_LSU/n254 ;
  wire \u_EXU_LSU/n255 ;
  wire \u_EXU_LSU/n256 ;
  wire \u_EXU_LSU/n257 ;
  wire \u_EXU_LSU/n258 ;
  wire \u_EXU_LSU/n259 ;
  wire \u_EXU_LSU/n26 ;
  wire \u_EXU_LSU/n260 ;
  wire \u_EXU_LSU/n261 ;
  wire \u_EXU_LSU/n262 ;
  wire \u_EXU_LSU/n263 ;
  wire \u_EXU_LSU/n264 ;
  wire \u_EXU_LSU/n265 ;
  wire \u_EXU_LSU/n266 ;
  wire \u_EXU_LSU/n267 ;
  wire \u_EXU_LSU/n268 ;
  wire \u_EXU_LSU/n269 ;
  wire \u_EXU_LSU/n270 ;
  wire \u_EXU_LSU/n271 ;
  wire \u_EXU_LSU/n272 ;
  wire \u_EXU_LSU/n273 ;
  wire \u_EXU_LSU/n274 ;
  wire \u_EXU_LSU/n275 ;
  wire \u_EXU_LSU/n276 ;
  wire \u_EXU_LSU/n277 ;
  wire \u_EXU_LSU/n278 ;
  wire \u_EXU_LSU/n279 ;
  wire \u_EXU_LSU/n280 ;
  wire \u_EXU_LSU/n281 ;
  wire \u_EXU_LSU/n282 ;
  wire \u_EXU_LSU/n283 ;
  wire \u_EXU_LSU/n284 ;
  wire \u_EXU_LSU/n3 ;
  wire \u_EXU_LSU/n30 ;
  wire \u_EXU_LSU/n37 ;
  wire \u_EXU_LSU/n38 ;
  wire \u_EXU_LSU/n39 ;
  wire \u_EXU_LSU/n4 ;
  wire \u_EXU_LSU/n40 ;
  wire \u_EXU_LSU/n41 ;
  wire \u_EXU_LSU/n42 ;
  wire \u_EXU_LSU/n43 ;
  wire \u_EXU_LSU/n44 ;
  wire \u_EXU_LSU/n45 ;
  wire \u_EXU_LSU/n46 ;
  wire \u_EXU_LSU/n47 ;
  wire \u_EXU_LSU/n48 ;
  wire \u_EXU_LSU/n5 ;
  wire \u_EXU_LSU/n56 ;
  wire \u_EXU_LSU/n57 ;
  wire \u_EXU_LSU/n58 ;
  wire \u_EXU_LSU/n58_neg ;
  wire \u_EXU_LSU/n66[1]_neg ;
  wire \u_EXU_LSU/n68 ;
  wire \u_EXU_LSU/n69 ;
  wire \u_EXU_LSU/n7 ;
  wire \u_EXU_LSU/n70 ;
  wire \u_EXU_LSU/n75 ;
  wire \u_EXU_LSU/n8 ;
  wire \u_EXU_LSU/n80 ;
  wire \u_EXU_LSU/n81 ;
  wire \u_EXU_LSU/n82 ;
  wire \u_EXU_LSU/n83 ;
  wire \u_EXU_LSU/n84 ;
  wire \u_EXU_LSU/n85 ;
  wire \u_EXU_LSU/n86 ;
  wire \u_EXU_LSU/n87 ;
  wire \u_EXU_LSU/n88 ;
  wire \u_EXU_LSU/n89 ;
  wire \u_EXU_LSU/n9 ;
  wire \u_EXU_LSU/n90 ;
  wire \u_EXU_LSU/n91 ;
  wire \u_EXU_LSU/n96 ;
  wire \u_EXU_LSU/n97 ;
  wire \u_EXU_LSU/n98 ;
  wire \u_EXU_LSU/n99 ;
  wire \u_EXU_LSU/sub0_2_co ;
  wire \u_EXU_LSU/sub0_2_co_neg ;
  wire \u_EXU_LSU/trans_finish ;  // ../RTL/core/exu_lsu.v(71)
  wire \u_EXU_LSU/u21_sel_is_2_o ;
  wire \u_EXU_LSU/u21_sel_is_2_o_neg ;
  wire \u_EXU_LSU/u22_sel_is_0_o ;
  wire \u_EXU_LSU/u29_sel_is_0_o ;
  wire \u_EXU_LSU/u336_sel_is_0_o ;
  wire \u_EXU_LSU/working ;  // ../RTL/core/exu_lsu.v(91)

  assign o_csridx[11] = i_csridx[11];
  assign o_csridx[10] = i_csridx[10];
  assign o_csridx[9] = i_csridx[9];
  assign o_csridx[8] = i_csridx[8];
  assign o_csridx[7] = i_csridx[7];
  assign o_csridx[6] = i_csridx[6];
  assign o_csridx[5] = i_csridx[5];
  assign o_csridx[4] = i_csridx[4];
  assign o_csridx[3] = i_csridx[3];
  assign o_csridx[2] = i_csridx[2];
  assign o_csridx[1] = i_csridx[1];
  assign o_csridx[0] = i_csridx[0];
  assign o_rdidx0[4] = i_rdidx[4];
  assign o_rdidx0[3] = i_rdidx[3];
  assign o_rdidx0[2] = i_rdidx[2];
  assign o_rdidx0[1] = i_rdidx[1];
  assign o_rdidx0[0] = i_rdidx[0];
  assign o_exu_rdwen0 = i_rdwen;
  assign o_exu_rdidx0[4] = i_rdidx[4];
  assign o_exu_rdidx0[3] = i_rdidx[3];
  assign o_exu_rdidx0[2] = i_rdidx[2];
  assign o_exu_rdidx0[1] = i_rdidx[1];
  assign o_exu_rdidx0[0] = i_rdidx[0];
  assign o_exu_rdidx2[4] = o_rdidx2[4];
  assign o_exu_rdidx2[3] = o_rdidx2[3];
  assign o_exu_rdidx2[2] = o_rdidx2[2];
  assign o_exu_rdidx2[1] = o_rdidx2[1];
  assign o_exu_rdidx2[0] = o_rdidx2[0];
  assign o_ribm_addr[1] = 1'b0;
  assign o_ribm_addr[0] = 1'b0;
  assign o_ribm_rdy = i_ribm_rsp;
  not \alu2lsu_result[1]_inv  (\alu2lsu_result[1]_neg , alu2lsu_result[1]);
  eq_w5 eq0 (
    .i0(o_rdidx0),
    .i1(o_exu_rdidx1),
    .o(n5));  // ../RTL/core/exu.v(172)
  eq_w5 eq1 (
    .i0(o_rdidx0),
    .i1(o_rdidx2),
    .o(n7));  // ../RTL/core/exu.v(209)
  not \i_decinfo[2]_inv  (\i_decinfo[2]_neg , i_decinfo[2]);
  not \i_decinfo[3]_inv  (\i_decinfo[3]_neg , i_decinfo[3]);
  not \i_decinfo[4]_inv  (\i_decinfo[4]_neg , i_decinfo[4]);
  not \i_exu_op2[4]_inv  (\i_exu_op2[4]_neg , i_exu_op2[4]);
  binary_mux_s1_w1 mux0_b0 (
    .i0(1'b0),
    .i1(i_csr_rdata[0]),
    .sel(i_decinfo_grp[4]),
    .o(n2[0]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b1 (
    .i0(1'b0),
    .i1(i_csr_rdata[1]),
    .sel(i_decinfo_grp[4]),
    .o(n2[1]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b10 (
    .i0(1'b0),
    .i1(i_csr_rdata[10]),
    .sel(i_decinfo_grp[4]),
    .o(n2[10]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b11 (
    .i0(1'b0),
    .i1(i_csr_rdata[11]),
    .sel(i_decinfo_grp[4]),
    .o(n2[11]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b12 (
    .i0(1'b0),
    .i1(i_csr_rdata[12]),
    .sel(i_decinfo_grp[4]),
    .o(n2[12]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b13 (
    .i0(1'b0),
    .i1(i_csr_rdata[13]),
    .sel(i_decinfo_grp[4]),
    .o(n2[13]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b14 (
    .i0(1'b0),
    .i1(i_csr_rdata[14]),
    .sel(i_decinfo_grp[4]),
    .o(n2[14]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b15 (
    .i0(1'b0),
    .i1(i_csr_rdata[15]),
    .sel(i_decinfo_grp[4]),
    .o(n2[15]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b16 (
    .i0(1'b0),
    .i1(i_csr_rdata[16]),
    .sel(i_decinfo_grp[4]),
    .o(n2[16]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b17 (
    .i0(1'b0),
    .i1(i_csr_rdata[17]),
    .sel(i_decinfo_grp[4]),
    .o(n2[17]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b18 (
    .i0(1'b0),
    .i1(i_csr_rdata[18]),
    .sel(i_decinfo_grp[4]),
    .o(n2[18]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b19 (
    .i0(1'b0),
    .i1(i_csr_rdata[19]),
    .sel(i_decinfo_grp[4]),
    .o(n2[19]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b2 (
    .i0(1'b0),
    .i1(i_csr_rdata[2]),
    .sel(i_decinfo_grp[4]),
    .o(n2[2]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b20 (
    .i0(1'b0),
    .i1(i_csr_rdata[20]),
    .sel(i_decinfo_grp[4]),
    .o(n2[20]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b21 (
    .i0(1'b0),
    .i1(i_csr_rdata[21]),
    .sel(i_decinfo_grp[4]),
    .o(n2[21]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b22 (
    .i0(1'b0),
    .i1(i_csr_rdata[22]),
    .sel(i_decinfo_grp[4]),
    .o(n2[22]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b23 (
    .i0(1'b0),
    .i1(i_csr_rdata[23]),
    .sel(i_decinfo_grp[4]),
    .o(n2[23]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b24 (
    .i0(1'b0),
    .i1(i_csr_rdata[24]),
    .sel(i_decinfo_grp[4]),
    .o(n2[24]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b25 (
    .i0(1'b0),
    .i1(i_csr_rdata[25]),
    .sel(i_decinfo_grp[4]),
    .o(n2[25]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b26 (
    .i0(1'b0),
    .i1(i_csr_rdata[26]),
    .sel(i_decinfo_grp[4]),
    .o(n2[26]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b27 (
    .i0(1'b0),
    .i1(i_csr_rdata[27]),
    .sel(i_decinfo_grp[4]),
    .o(n2[27]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b28 (
    .i0(1'b0),
    .i1(i_csr_rdata[28]),
    .sel(i_decinfo_grp[4]),
    .o(n2[28]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b29 (
    .i0(1'b0),
    .i1(i_csr_rdata[29]),
    .sel(i_decinfo_grp[4]),
    .o(n2[29]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b3 (
    .i0(1'b0),
    .i1(i_csr_rdata[3]),
    .sel(i_decinfo_grp[4]),
    .o(n2[3]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b30 (
    .i0(1'b0),
    .i1(i_csr_rdata[30]),
    .sel(i_decinfo_grp[4]),
    .o(n2[30]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b31 (
    .i0(1'b0),
    .i1(i_csr_rdata[31]),
    .sel(i_decinfo_grp[4]),
    .o(n2[31]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b4 (
    .i0(1'b0),
    .i1(i_csr_rdata[4]),
    .sel(i_decinfo_grp[4]),
    .o(n2[4]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b5 (
    .i0(1'b0),
    .i1(i_csr_rdata[5]),
    .sel(i_decinfo_grp[4]),
    .o(n2[5]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b6 (
    .i0(1'b0),
    .i1(i_csr_rdata[6]),
    .sel(i_decinfo_grp[4]),
    .o(n2[6]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b7 (
    .i0(1'b0),
    .i1(i_csr_rdata[7]),
    .sel(i_decinfo_grp[4]),
    .o(n2[7]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b8 (
    .i0(1'b0),
    .i1(i_csr_rdata[8]),
    .sel(i_decinfo_grp[4]),
    .o(n2[8]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux0_b9 (
    .i0(1'b0),
    .i1(i_csr_rdata[9]),
    .sel(i_decinfo_grp[4]),
    .o(n2[9]));  // ../RTL/core/exu.v(159)
  binary_mux_s1_w1 mux1_b0 (
    .i0(n2[0]),
    .i1(i_iaddr[0]),
    .sel(bju_rdwen),
    .o(n3[0]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b1 (
    .i0(n2[1]),
    .i1(i_iaddr[1]),
    .sel(bju_rdwen),
    .o(n3[1]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b10 (
    .i0(n2[10]),
    .i1(bju_rdwdata[10]),
    .sel(bju_rdwen),
    .o(n3[10]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b11 (
    .i0(n2[11]),
    .i1(bju_rdwdata[11]),
    .sel(bju_rdwen),
    .o(n3[11]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b12 (
    .i0(n2[12]),
    .i1(bju_rdwdata[12]),
    .sel(bju_rdwen),
    .o(n3[12]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b13 (
    .i0(n2[13]),
    .i1(bju_rdwdata[13]),
    .sel(bju_rdwen),
    .o(n3[13]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b14 (
    .i0(n2[14]),
    .i1(bju_rdwdata[14]),
    .sel(bju_rdwen),
    .o(n3[14]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b15 (
    .i0(n2[15]),
    .i1(bju_rdwdata[15]),
    .sel(bju_rdwen),
    .o(n3[15]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b16 (
    .i0(n2[16]),
    .i1(bju_rdwdata[16]),
    .sel(bju_rdwen),
    .o(n3[16]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b17 (
    .i0(n2[17]),
    .i1(bju_rdwdata[17]),
    .sel(bju_rdwen),
    .o(n3[17]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b18 (
    .i0(n2[18]),
    .i1(bju_rdwdata[18]),
    .sel(bju_rdwen),
    .o(n3[18]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b19 (
    .i0(n2[19]),
    .i1(bju_rdwdata[19]),
    .sel(bju_rdwen),
    .o(n3[19]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b2 (
    .i0(n2[2]),
    .i1(bju_rdwdata[2]),
    .sel(bju_rdwen),
    .o(n3[2]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b20 (
    .i0(n2[20]),
    .i1(bju_rdwdata[20]),
    .sel(bju_rdwen),
    .o(n3[20]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b21 (
    .i0(n2[21]),
    .i1(bju_rdwdata[21]),
    .sel(bju_rdwen),
    .o(n3[21]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b22 (
    .i0(n2[22]),
    .i1(bju_rdwdata[22]),
    .sel(bju_rdwen),
    .o(n3[22]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b23 (
    .i0(n2[23]),
    .i1(bju_rdwdata[23]),
    .sel(bju_rdwen),
    .o(n3[23]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b24 (
    .i0(n2[24]),
    .i1(bju_rdwdata[24]),
    .sel(bju_rdwen),
    .o(n3[24]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b25 (
    .i0(n2[25]),
    .i1(bju_rdwdata[25]),
    .sel(bju_rdwen),
    .o(n3[25]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b26 (
    .i0(n2[26]),
    .i1(bju_rdwdata[26]),
    .sel(bju_rdwen),
    .o(n3[26]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b27 (
    .i0(n2[27]),
    .i1(bju_rdwdata[27]),
    .sel(bju_rdwen),
    .o(n3[27]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b28 (
    .i0(n2[28]),
    .i1(bju_rdwdata[28]),
    .sel(bju_rdwen),
    .o(n3[28]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b29 (
    .i0(n2[29]),
    .i1(bju_rdwdata[29]),
    .sel(bju_rdwen),
    .o(n3[29]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b3 (
    .i0(n2[3]),
    .i1(bju_rdwdata[3]),
    .sel(bju_rdwen),
    .o(n3[3]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b30 (
    .i0(n2[30]),
    .i1(bju_rdwdata[30]),
    .sel(bju_rdwen),
    .o(n3[30]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b31 (
    .i0(n2[31]),
    .i1(bju_rdwdata[31]),
    .sel(bju_rdwen),
    .o(n3[31]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b4 (
    .i0(n2[4]),
    .i1(bju_rdwdata[4]),
    .sel(bju_rdwen),
    .o(n3[4]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b5 (
    .i0(n2[5]),
    .i1(bju_rdwdata[5]),
    .sel(bju_rdwen),
    .o(n3[5]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b6 (
    .i0(n2[6]),
    .i1(bju_rdwdata[6]),
    .sel(bju_rdwen),
    .o(n3[6]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b7 (
    .i0(n2[7]),
    .i1(bju_rdwdata[7]),
    .sel(bju_rdwen),
    .o(n3[7]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b8 (
    .i0(n2[8]),
    .i1(bju_rdwdata[8]),
    .sel(bju_rdwen),
    .o(n3[8]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux1_b9 (
    .i0(n2[9]),
    .i1(bju_rdwdata[9]),
    .sel(bju_rdwen),
    .o(n3[9]));  // ../RTL/core/exu.v(158)
  binary_mux_s1_w1 mux2_b0 (
    .i0(n3[0]),
    .i1(alu_rdwdata[0]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[0]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b1 (
    .i0(n3[1]),
    .i1(\u_EXU_ALU/n309 [1]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[1]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b10 (
    .i0(n3[10]),
    .i1(\u_EXU_ALU/n309 [10]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[10]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b11 (
    .i0(n3[11]),
    .i1(\u_EXU_ALU/n309 [11]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[11]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b12 (
    .i0(n3[12]),
    .i1(\u_EXU_ALU/n309 [12]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[12]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b13 (
    .i0(n3[13]),
    .i1(\u_EXU_ALU/n309 [13]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[13]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b14 (
    .i0(n3[14]),
    .i1(\u_EXU_ALU/n309 [14]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[14]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b15 (
    .i0(n3[15]),
    .i1(\u_EXU_ALU/n309 [15]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[15]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b16 (
    .i0(n3[16]),
    .i1(\u_EXU_ALU/n309 [16]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[16]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b17 (
    .i0(n3[17]),
    .i1(\u_EXU_ALU/n309 [17]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[17]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b18 (
    .i0(n3[18]),
    .i1(\u_EXU_ALU/n309 [18]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[18]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b19 (
    .i0(n3[19]),
    .i1(\u_EXU_ALU/n309 [19]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[19]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b2 (
    .i0(n3[2]),
    .i1(\u_EXU_ALU/n309 [2]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[2]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b20 (
    .i0(n3[20]),
    .i1(\u_EXU_ALU/n309 [20]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[20]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b21 (
    .i0(n3[21]),
    .i1(\u_EXU_ALU/n309 [21]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[21]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b22 (
    .i0(n3[22]),
    .i1(\u_EXU_ALU/n309 [22]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[22]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b23 (
    .i0(n3[23]),
    .i1(\u_EXU_ALU/n309 [23]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[23]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b24 (
    .i0(n3[24]),
    .i1(\u_EXU_ALU/n309 [24]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[24]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b25 (
    .i0(n3[25]),
    .i1(\u_EXU_ALU/n309 [25]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[25]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b26 (
    .i0(n3[26]),
    .i1(\u_EXU_ALU/n309 [26]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[26]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b27 (
    .i0(n3[27]),
    .i1(\u_EXU_ALU/n309 [27]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[27]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b28 (
    .i0(n3[28]),
    .i1(\u_EXU_ALU/n309 [28]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[28]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b29 (
    .i0(n3[29]),
    .i1(\u_EXU_ALU/n309 [29]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[29]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b3 (
    .i0(n3[3]),
    .i1(\u_EXU_ALU/n309 [3]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[3]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b30 (
    .i0(n3[30]),
    .i1(\u_EXU_ALU/n309 [30]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[30]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b31 (
    .i0(n3[31]),
    .i1(\u_EXU_ALU/n309 [31]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[31]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b4 (
    .i0(n3[4]),
    .i1(\u_EXU_ALU/n309 [4]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[4]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b5 (
    .i0(n3[5]),
    .i1(\u_EXU_ALU/n309 [5]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[5]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b6 (
    .i0(n3[6]),
    .i1(\u_EXU_ALU/n309 [6]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[6]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b7 (
    .i0(n3[7]),
    .i1(\u_EXU_ALU/n309 [7]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[7]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b8 (
    .i0(n3[8]),
    .i1(\u_EXU_ALU/n309 [8]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[8]));  // ../RTL/core/exu.v(157)
  binary_mux_s1_w1 mux2_b9 (
    .i0(n3[9]),
    .i1(\u_EXU_ALU/n309 [9]),
    .sel(i_decinfo_grp[0]),
    .o(o_rdwdata0[9]));  // ../RTL/core/exu.v(157)
  and u10 (n4, o_exu_rdwen0, o_exu_rdwen1);  // ../RTL/core/exu.v(172)
  AL_MUX u11 (
    .i0(1'b0),
    .i1(n5),
    .sel(n4),
    .o(mdu_flush));  // ../RTL/core/exu.v(172)
  and u13 (n6, o_exu_rdwen0, o_exu_rdwen2);  // ../RTL/core/exu.v(209)
  AL_MUX u14 (
    .i0(1'b0),
    .i1(n7),
    .sel(n6),
    .o(lsu_flush));  // ../RTL/core/exu.v(209)
  and u16 (n8, i_decinfo_grp[3], o_mdu_working);  // ../RTL/core/exu.v(249)
  and u17 (n9, i_decinfo_grp[1], o_lsu_working);  // ../RTL/core/exu.v(250)
  or u18 (o_exu_resource_match, n8, n9);  // ../RTL/core/exu.v(249)
  or u4 (n0, i_decinfo_grp[0], bju_rdwen);  // ../RTL/core/exu.v(155)
  or u5 (n1, n0, i_decinfo_grp[4]);  // ../RTL/core/exu.v(155)
  and u6 (o_rdwen0, n1, o_exu_rdwen0);  // ../RTL/core/exu.v(155)
  add_pu32_pu32_o32 \u_EXU_ALU/add0  (
    .i0(i_exu_op1),
    .i1(i_exu_op2),
    .o(\u_EXU_ALU/n0 ));  // ../RTL/core/exu_alu.v(39)
  lt_u32_u32 \u_EXU_ALU/lt0  (
    .ci(1'b0),
    .i0({i_exu_op2[31],i_exu_op1[30:0]}),
    .i1({i_exu_op1[31],i_exu_op2[30:0]}),
    .o(\u_EXU_ALU/n253 ));  // ../RTL/core/exu_alu.v(55)
  lt_u32_u32 \u_EXU_ALU/lt1  (
    .ci(1'b0),
    .i0(i_exu_op1),
    .i1(i_exu_op2),
    .o(\u_EXU_ALU/n261 ));  // ../RTL/core/exu_alu.v(57)
  not \u_EXU_ALU/n179_inv  (\u_EXU_ALU/n179_neg , \u_EXU_ALU/n179 );
  not \u_EXU_ALU/n281_inv  (\u_EXU_ALU/n281_neg , \u_EXU_ALU/n281 );
  add_pu32_mu32_o32 \u_EXU_ALU/sub0  (
    .i0(i_exu_op1),
    .i1(i_exu_op2),
    .o(\u_EXU_ALU/n33 ));  // ../RTL/core/exu_alu.v(41)
  or \u_EXU_ALU/u10  (alu_rdwdata[0], \u_EXU_ALU/n310 [0], \u_EXU_ALU/alu_sltu [0]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u100  (\u_EXU_ALU/n309 [11], \u_EXU_ALU/n308 [11], \u_EXU_ALU/alu_or [11]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u1000  (\u_EXU_ALU/n293 , i_exu_op2[18], \u_EXU_ALU/n461 );  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u1001  (\u_EXU_ALU/n292 , i_exu_op2[21], i_exu_op2[22]);  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u1002  (\u_EXU_ALU/n291 , i_exu_op2[23], i_exu_op2[24]);  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u1003  (\u_EXU_ALU/n290 , \u_EXU_ALU/n292 , \u_EXU_ALU/n291 );  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u1004  (\u_EXU_ALU/n289 , \u_EXU_ALU/n293 , \u_EXU_ALU/n290 );  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u1005  (\u_EXU_ALU/n288 , i_exu_op2[26], i_exu_op2[27]);  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u1006  (\u_EXU_ALU/n287 , i_exu_op2[25], \u_EXU_ALU/n288 );  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u1007  (\u_EXU_ALU/n286 , i_exu_op2[28], i_exu_op2[29]);  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u1008  (\u_EXU_ALU/n285 , i_exu_op2[30], i_exu_op2[31]);  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u1009  (\u_EXU_ALU/n284 , \u_EXU_ALU/n286 , \u_EXU_ALU/n285 );  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u101  (\u_EXU_ALU/n309 [12], \u_EXU_ALU/n308 [12], \u_EXU_ALU/alu_or [12]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u1010  (\u_EXU_ALU/n283 , \u_EXU_ALU/n287 , \u_EXU_ALU/n284 );  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u1011  (\u_EXU_ALU/n282 , \u_EXU_ALU/n289 , \u_EXU_ALU/n283 );  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u1012  (\u_EXU_ALU/n281 , \u_EXU_ALU/n460 , \u_EXU_ALU/n282 );  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1013  (
    .i0(\u_EXU_ALU/n43 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [0]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1014  (
    .i0(\u_EXU_ALU/n42 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [1]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1015  (
    .i0(\u_EXU_ALU/n41 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [2]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1016  (
    .i0(\u_EXU_ALU/n40 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [3]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1017  (
    .i0(\u_EXU_ALU/n39 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [4]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1018  (
    .i0(\u_EXU_ALU/n38 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [5]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1019  (
    .i0(\u_EXU_ALU/n37 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [6]));  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u102  (\u_EXU_ALU/n309 [13], \u_EXU_ALU/n308 [13], \u_EXU_ALU/alu_or [13]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1020  (
    .i0(\u_EXU_ALU/n36 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [7]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1021  (
    .i0(\u_EXU_ALU/n35 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [8]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1022  (
    .i0(\u_EXU_ALU/n34 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [9]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1023  (
    .i0(\u_EXU_ALU/n32 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [10]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1024  (
    .i0(\u_EXU_ALU/n31 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [11]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1025  (
    .i0(\u_EXU_ALU/n30 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [12]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1026  (
    .i0(\u_EXU_ALU/n29 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [13]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1027  (
    .i0(\u_EXU_ALU/n28 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [14]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1028  (
    .i0(\u_EXU_ALU/n27 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n99 [15]));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u1029  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n59 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [16]));
  and \u_EXU_ALU/u1029_sel_is_0  (\u_EXU_ALU/u1029_sel_is_0_o , \u_EXU_ALU/n281_neg , \i_exu_op2[4]_neg );
  or \u_EXU_ALU/u103  (\u_EXU_ALU/n309 [14], \u_EXU_ALU/n308 [14], \u_EXU_ALU/alu_or [14]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1030  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n58 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [17]));
  AL_MUX \u_EXU_ALU/u1031  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n57 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [18]));
  AL_MUX \u_EXU_ALU/u1032  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n56 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [19]));
  AL_MUX \u_EXU_ALU/u1033  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n55 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [20]));
  AL_MUX \u_EXU_ALU/u1034  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n54 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [21]));
  AL_MUX \u_EXU_ALU/u1035  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n53 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [22]));
  AL_MUX \u_EXU_ALU/u1036  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n52 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [23]));
  AL_MUX \u_EXU_ALU/u1037  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n51 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [24]));
  AL_MUX \u_EXU_ALU/u1038  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n50 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [25]));
  AL_MUX \u_EXU_ALU/u1039  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n49 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [26]));
  or \u_EXU_ALU/u104  (\u_EXU_ALU/n309 [15], \u_EXU_ALU/n308 [15], \u_EXU_ALU/alu_or [15]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1040  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n48 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [27]));
  AL_MUX \u_EXU_ALU/u1041  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n47 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [28]));
  AL_MUX \u_EXU_ALU/u1042  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n46 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [29]));
  AL_MUX \u_EXU_ALU/u1043  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n45 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [30]));
  AL_MUX \u_EXU_ALU/u1044  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n44 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n99 [31]));
  and \u_EXU_ALU/u1045  (\u_EXU_ALU/alu_sll [1], i_decinfo[2], \u_EXU_ALU/n66 [1]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1046  (\u_EXU_ALU/alu_sll [2], i_decinfo[2], \u_EXU_ALU/n66 [2]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1047  (\u_EXU_ALU/alu_sll [3], i_decinfo[2], \u_EXU_ALU/n66 [3]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1048  (\u_EXU_ALU/alu_sll [4], i_decinfo[2], \u_EXU_ALU/n66 [4]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1049  (\u_EXU_ALU/alu_sll [5], i_decinfo[2], \u_EXU_ALU/n66 [5]);  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u105  (\u_EXU_ALU/n309 [16], \u_EXU_ALU/n308 [16], \u_EXU_ALU/alu_or [16]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u1050  (\u_EXU_ALU/alu_sll [6], i_decinfo[2], \u_EXU_ALU/n66 [6]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1051  (\u_EXU_ALU/alu_sll [7], i_decinfo[2], \u_EXU_ALU/n66 [7]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1052  (\u_EXU_ALU/alu_sll [8], i_decinfo[2], \u_EXU_ALU/n66 [8]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1053  (\u_EXU_ALU/alu_sll [9], i_decinfo[2], \u_EXU_ALU/n66 [9]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1054  (\u_EXU_ALU/alu_sll [10], i_decinfo[2], \u_EXU_ALU/n66 [10]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1055  (\u_EXU_ALU/alu_sll [11], i_decinfo[2], \u_EXU_ALU/n66 [11]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1056  (\u_EXU_ALU/alu_sll [12], i_decinfo[2], \u_EXU_ALU/n66 [12]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1057  (\u_EXU_ALU/alu_sll [13], i_decinfo[2], \u_EXU_ALU/n66 [13]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1058  (\u_EXU_ALU/alu_sll [14], i_decinfo[2], \u_EXU_ALU/n66 [14]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1059  (\u_EXU_ALU/alu_sll [15], i_decinfo[2], \u_EXU_ALU/n66 [15]);  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u106  (\u_EXU_ALU/n309 [17], \u_EXU_ALU/n308 [17], \u_EXU_ALU/alu_or [17]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u1060  (\u_EXU_ALU/alu_sll [16], i_decinfo[2], \u_EXU_ALU/n66 [16]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1061  (\u_EXU_ALU/alu_sll [17], i_decinfo[2], \u_EXU_ALU/n66 [17]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1062  (\u_EXU_ALU/alu_sll [18], i_decinfo[2], \u_EXU_ALU/n66 [18]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1063  (\u_EXU_ALU/alu_sll [19], i_decinfo[2], \u_EXU_ALU/n66 [19]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1064  (\u_EXU_ALU/alu_sll [20], i_decinfo[2], \u_EXU_ALU/n66 [20]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1065  (\u_EXU_ALU/alu_sll [21], i_decinfo[2], \u_EXU_ALU/n66 [21]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1066  (\u_EXU_ALU/alu_sll [22], i_decinfo[2], \u_EXU_ALU/n66 [22]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1067  (\u_EXU_ALU/alu_sll [23], i_decinfo[2], \u_EXU_ALU/n66 [23]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1068  (\u_EXU_ALU/alu_sll [24], i_decinfo[2], \u_EXU_ALU/n66 [24]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1069  (\u_EXU_ALU/alu_sll [25], i_decinfo[2], \u_EXU_ALU/n66 [25]);  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u107  (\u_EXU_ALU/n309 [18], \u_EXU_ALU/n308 [18], \u_EXU_ALU/alu_or [18]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u1070  (\u_EXU_ALU/alu_sll [26], i_decinfo[2], \u_EXU_ALU/n66 [26]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1071  (\u_EXU_ALU/alu_sll [27], i_decinfo[2], \u_EXU_ALU/n66 [27]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1072  (\u_EXU_ALU/alu_sll [28], i_decinfo[2], \u_EXU_ALU/n66 [28]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1073  (\u_EXU_ALU/alu_sll [29], i_decinfo[2], \u_EXU_ALU/n66 [29]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1074  (\u_EXU_ALU/alu_sll [30], i_decinfo[2], \u_EXU_ALU/n66 [30]);  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u1075  (\u_EXU_ALU/alu_sll [31], i_decinfo[2], \u_EXU_ALU/n66 [31]);  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1076  (
    .i0(i_exu_op1[30]),
    .i1(i_exu_op1[29]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n279 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1077  (
    .i0(i_exu_op1[29]),
    .i1(i_exu_op1[28]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n278 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1078  (
    .i0(i_exu_op1[28]),
    .i1(i_exu_op1[27]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n277 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1079  (
    .i0(i_exu_op1[27]),
    .i1(i_exu_op1[26]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n276 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u108  (\u_EXU_ALU/n309 [19], \u_EXU_ALU/n308 [19], \u_EXU_ALU/alu_or [19]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1080  (
    .i0(i_exu_op1[26]),
    .i1(i_exu_op1[25]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n275 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1081  (
    .i0(i_exu_op1[25]),
    .i1(i_exu_op1[24]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n274 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1082  (
    .i0(i_exu_op1[24]),
    .i1(i_exu_op1[23]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n273 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1083  (
    .i0(i_exu_op1[23]),
    .i1(i_exu_op1[22]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n272 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1084  (
    .i0(i_exu_op1[22]),
    .i1(i_exu_op1[21]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n271 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1085  (
    .i0(i_exu_op1[21]),
    .i1(i_exu_op1[20]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n270 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1086  (
    .i0(i_exu_op1[20]),
    .i1(i_exu_op1[19]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n269 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1087  (
    .i0(i_exu_op1[19]),
    .i1(i_exu_op1[18]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n268 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1088  (
    .i0(i_exu_op1[18]),
    .i1(i_exu_op1[17]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n267 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1089  (
    .i0(i_exu_op1[17]),
    .i1(i_exu_op1[16]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n266 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u109  (\u_EXU_ALU/n309 [20], \u_EXU_ALU/n308 [20], \u_EXU_ALU/alu_or [20]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1090  (
    .i0(i_exu_op1[16]),
    .i1(i_exu_op1[15]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n265 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1091  (
    .i0(i_exu_op1[15]),
    .i1(i_exu_op1[14]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n342 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1092  (
    .i0(i_exu_op1[14]),
    .i1(i_exu_op1[13]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n341 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1093  (
    .i0(i_exu_op1[13]),
    .i1(i_exu_op1[12]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n340 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1094  (
    .i0(i_exu_op1[12]),
    .i1(i_exu_op1[11]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n339 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1095  (
    .i0(i_exu_op1[11]),
    .i1(i_exu_op1[10]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n338 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1096  (
    .i0(i_exu_op1[10]),
    .i1(i_exu_op1[9]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n337 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1097  (
    .i0(i_exu_op1[9]),
    .i1(i_exu_op1[8]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n336 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1098  (
    .i0(i_exu_op1[8]),
    .i1(i_exu_op1[7]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n335 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1099  (
    .i0(i_exu_op1[7]),
    .i1(i_exu_op1[6]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n334 ));  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u11  (\u_EXU_ALU/alu_sra [0], i_decinfo[4], \u_EXU_ALU/n99 [0]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u110  (\u_EXU_ALU/n309 [21], \u_EXU_ALU/n308 [21], \u_EXU_ALU/alu_or [21]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1100  (
    .i0(i_exu_op1[6]),
    .i1(i_exu_op1[5]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n333 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1101  (
    .i0(i_exu_op1[5]),
    .i1(i_exu_op1[4]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n332 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1102  (
    .i0(i_exu_op1[4]),
    .i1(i_exu_op1[3]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n331 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1103  (
    .i0(i_exu_op1[3]),
    .i1(i_exu_op1[2]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n330 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1104  (
    .i0(i_exu_op1[2]),
    .i1(i_exu_op1[1]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n329 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1105  (
    .i0(i_exu_op1[1]),
    .i1(i_exu_op1[0]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n328 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1106  (
    .i0(i_exu_op1[0]),
    .i1(1'b0),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n327 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1107  (
    .i0(\u_EXU_ALU/n280 ),
    .i1(\u_EXU_ALU/n278 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n326 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1108  (
    .i0(\u_EXU_ALU/n279 ),
    .i1(\u_EXU_ALU/n277 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n325 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1109  (
    .i0(\u_EXU_ALU/n278 ),
    .i1(\u_EXU_ALU/n276 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n324 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u111  (\u_EXU_ALU/n309 [22], \u_EXU_ALU/n308 [22], \u_EXU_ALU/alu_or [22]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1110  (
    .i0(\u_EXU_ALU/n277 ),
    .i1(\u_EXU_ALU/n275 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n323 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1111  (
    .i0(\u_EXU_ALU/n276 ),
    .i1(\u_EXU_ALU/n274 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n322 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1112  (
    .i0(\u_EXU_ALU/n275 ),
    .i1(\u_EXU_ALU/n273 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n321 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1113  (
    .i0(\u_EXU_ALU/n274 ),
    .i1(\u_EXU_ALU/n272 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n320 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1114  (
    .i0(\u_EXU_ALU/n273 ),
    .i1(\u_EXU_ALU/n271 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n319 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1115  (
    .i0(\u_EXU_ALU/n272 ),
    .i1(\u_EXU_ALU/n270 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n318 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1116  (
    .i0(\u_EXU_ALU/n271 ),
    .i1(\u_EXU_ALU/n269 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n317 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1117  (
    .i0(\u_EXU_ALU/n270 ),
    .i1(\u_EXU_ALU/n268 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n316 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1118  (
    .i0(\u_EXU_ALU/n269 ),
    .i1(\u_EXU_ALU/n267 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n315 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1119  (
    .i0(\u_EXU_ALU/n268 ),
    .i1(\u_EXU_ALU/n266 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n314 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u112  (\u_EXU_ALU/n309 [23], \u_EXU_ALU/n308 [23], \u_EXU_ALU/alu_or [23]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1120  (
    .i0(\u_EXU_ALU/n267 ),
    .i1(\u_EXU_ALU/n265 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n313 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1121  (
    .i0(\u_EXU_ALU/n266 ),
    .i1(\u_EXU_ALU/n342 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n312 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1122  (
    .i0(\u_EXU_ALU/n265 ),
    .i1(\u_EXU_ALU/n341 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n311 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1123  (
    .i0(\u_EXU_ALU/n342 ),
    .i1(\u_EXU_ALU/n340 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n302 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1124  (
    .i0(\u_EXU_ALU/n341 ),
    .i1(\u_EXU_ALU/n339 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n301 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1125  (
    .i0(\u_EXU_ALU/n340 ),
    .i1(\u_EXU_ALU/n338 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n300 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1126  (
    .i0(\u_EXU_ALU/n339 ),
    .i1(\u_EXU_ALU/n337 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n299 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1127  (
    .i0(\u_EXU_ALU/n338 ),
    .i1(\u_EXU_ALU/n336 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n298 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1128  (
    .i0(\u_EXU_ALU/n337 ),
    .i1(\u_EXU_ALU/n335 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n297 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1129  (
    .i0(\u_EXU_ALU/n336 ),
    .i1(\u_EXU_ALU/n334 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n343 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u113  (\u_EXU_ALU/n309 [24], \u_EXU_ALU/n308 [24], \u_EXU_ALU/alu_or [24]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1130  (
    .i0(\u_EXU_ALU/n335 ),
    .i1(\u_EXU_ALU/n333 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n344 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1131  (
    .i0(\u_EXU_ALU/n334 ),
    .i1(\u_EXU_ALU/n332 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n345 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1132  (
    .i0(\u_EXU_ALU/n333 ),
    .i1(\u_EXU_ALU/n331 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n346 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1133  (
    .i0(\u_EXU_ALU/n332 ),
    .i1(\u_EXU_ALU/n330 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n347 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1134  (
    .i0(\u_EXU_ALU/n331 ),
    .i1(\u_EXU_ALU/n329 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n348 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1135  (
    .i0(\u_EXU_ALU/n330 ),
    .i1(\u_EXU_ALU/n328 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n349 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1136  (
    .i0(\u_EXU_ALU/n329 ),
    .i1(\u_EXU_ALU/n327 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n350 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1137  (
    .i0(\u_EXU_ALU/n328 ),
    .i1(1'b0),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n351 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1138  (
    .i0(\u_EXU_ALU/n327 ),
    .i1(1'b0),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n352 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1139  (
    .i0(\u_EXU_ALU/n326 ),
    .i1(\u_EXU_ALU/n322 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n353 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u114  (\u_EXU_ALU/n309 [25], \u_EXU_ALU/n308 [25], \u_EXU_ALU/alu_or [25]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1140  (
    .i0(\u_EXU_ALU/n325 ),
    .i1(\u_EXU_ALU/n321 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n354 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1141  (
    .i0(\u_EXU_ALU/n324 ),
    .i1(\u_EXU_ALU/n320 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n355 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1142  (
    .i0(\u_EXU_ALU/n323 ),
    .i1(\u_EXU_ALU/n319 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n356 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1143  (
    .i0(\u_EXU_ALU/n322 ),
    .i1(\u_EXU_ALU/n318 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n357 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1144  (
    .i0(\u_EXU_ALU/n321 ),
    .i1(\u_EXU_ALU/n317 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n358 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1145  (
    .i0(\u_EXU_ALU/n320 ),
    .i1(\u_EXU_ALU/n316 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n359 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1146  (
    .i0(\u_EXU_ALU/n319 ),
    .i1(\u_EXU_ALU/n315 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n360 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1147  (
    .i0(\u_EXU_ALU/n318 ),
    .i1(\u_EXU_ALU/n314 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n361 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1148  (
    .i0(\u_EXU_ALU/n317 ),
    .i1(\u_EXU_ALU/n313 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n362 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1149  (
    .i0(\u_EXU_ALU/n316 ),
    .i1(\u_EXU_ALU/n312 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n363 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u115  (\u_EXU_ALU/n309 [26], \u_EXU_ALU/n308 [26], \u_EXU_ALU/alu_or [26]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1150  (
    .i0(\u_EXU_ALU/n315 ),
    .i1(\u_EXU_ALU/n311 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n364 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1151  (
    .i0(\u_EXU_ALU/n314 ),
    .i1(\u_EXU_ALU/n302 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n365 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1152  (
    .i0(\u_EXU_ALU/n313 ),
    .i1(\u_EXU_ALU/n301 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n366 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1153  (
    .i0(\u_EXU_ALU/n312 ),
    .i1(\u_EXU_ALU/n300 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n367 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1154  (
    .i0(\u_EXU_ALU/n311 ),
    .i1(\u_EXU_ALU/n299 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n368 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1155  (
    .i0(\u_EXU_ALU/n302 ),
    .i1(\u_EXU_ALU/n298 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n369 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1156  (
    .i0(\u_EXU_ALU/n301 ),
    .i1(\u_EXU_ALU/n297 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n370 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1157  (
    .i0(\u_EXU_ALU/n300 ),
    .i1(\u_EXU_ALU/n343 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n371 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1158  (
    .i0(\u_EXU_ALU/n299 ),
    .i1(\u_EXU_ALU/n344 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n372 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1159  (
    .i0(\u_EXU_ALU/n298 ),
    .i1(\u_EXU_ALU/n345 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n373 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u116  (\u_EXU_ALU/n309 [27], \u_EXU_ALU/n308 [27], \u_EXU_ALU/alu_or [27]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1160  (
    .i0(\u_EXU_ALU/n297 ),
    .i1(\u_EXU_ALU/n346 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n374 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1161  (
    .i0(\u_EXU_ALU/n343 ),
    .i1(\u_EXU_ALU/n347 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n375 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1162  (
    .i0(\u_EXU_ALU/n344 ),
    .i1(\u_EXU_ALU/n348 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n376 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1163  (
    .i0(\u_EXU_ALU/n345 ),
    .i1(\u_EXU_ALU/n349 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n377 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1164  (
    .i0(\u_EXU_ALU/n346 ),
    .i1(\u_EXU_ALU/n350 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n378 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1165  (
    .i0(\u_EXU_ALU/n347 ),
    .i1(\u_EXU_ALU/n351 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n379 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1166  (
    .i0(\u_EXU_ALU/n348 ),
    .i1(\u_EXU_ALU/n352 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n380 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1167  (
    .i0(\u_EXU_ALU/n349 ),
    .i1(1'b0),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n381 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1168  (
    .i0(\u_EXU_ALU/n350 ),
    .i1(1'b0),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n382 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1169  (
    .i0(\u_EXU_ALU/n351 ),
    .i1(1'b0),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n383 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u117  (\u_EXU_ALU/n309 [28], \u_EXU_ALU/n308 [28], \u_EXU_ALU/alu_or [28]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1170  (
    .i0(\u_EXU_ALU/n352 ),
    .i1(1'b0),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n384 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1171  (
    .i0(\u_EXU_ALU/n353 ),
    .i1(\u_EXU_ALU/n361 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n385 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1172  (
    .i0(\u_EXU_ALU/n354 ),
    .i1(\u_EXU_ALU/n362 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n386 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1173  (
    .i0(\u_EXU_ALU/n355 ),
    .i1(\u_EXU_ALU/n363 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n387 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1174  (
    .i0(\u_EXU_ALU/n356 ),
    .i1(\u_EXU_ALU/n364 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n388 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1175  (
    .i0(\u_EXU_ALU/n357 ),
    .i1(\u_EXU_ALU/n365 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n389 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1176  (
    .i0(\u_EXU_ALU/n358 ),
    .i1(\u_EXU_ALU/n366 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n390 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1177  (
    .i0(\u_EXU_ALU/n359 ),
    .i1(\u_EXU_ALU/n367 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n391 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1178  (
    .i0(\u_EXU_ALU/n360 ),
    .i1(\u_EXU_ALU/n368 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n392 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1179  (
    .i0(\u_EXU_ALU/n361 ),
    .i1(\u_EXU_ALU/n369 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n393 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u118  (\u_EXU_ALU/n309 [29], \u_EXU_ALU/n308 [29], \u_EXU_ALU/alu_or [29]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1180  (
    .i0(\u_EXU_ALU/n362 ),
    .i1(\u_EXU_ALU/n370 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n394 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1181  (
    .i0(\u_EXU_ALU/n363 ),
    .i1(\u_EXU_ALU/n371 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n395 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1182  (
    .i0(\u_EXU_ALU/n364 ),
    .i1(\u_EXU_ALU/n372 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n396 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1183  (
    .i0(\u_EXU_ALU/n365 ),
    .i1(\u_EXU_ALU/n373 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n397 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1184  (
    .i0(\u_EXU_ALU/n366 ),
    .i1(\u_EXU_ALU/n374 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n398 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1185  (
    .i0(\u_EXU_ALU/n367 ),
    .i1(\u_EXU_ALU/n375 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n399 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1186  (
    .i0(\u_EXU_ALU/n368 ),
    .i1(\u_EXU_ALU/n376 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n400 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1187  (
    .i0(\u_EXU_ALU/n369 ),
    .i1(\u_EXU_ALU/n377 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n401 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1188  (
    .i0(\u_EXU_ALU/n370 ),
    .i1(\u_EXU_ALU/n378 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n402 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1189  (
    .i0(\u_EXU_ALU/n371 ),
    .i1(\u_EXU_ALU/n379 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n403 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u119  (\u_EXU_ALU/n309 [30], \u_EXU_ALU/n308 [30], \u_EXU_ALU/alu_or [30]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1190  (
    .i0(\u_EXU_ALU/n372 ),
    .i1(\u_EXU_ALU/n380 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n404 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1191  (
    .i0(\u_EXU_ALU/n373 ),
    .i1(\u_EXU_ALU/n381 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n405 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1192  (
    .i0(\u_EXU_ALU/n374 ),
    .i1(\u_EXU_ALU/n382 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n406 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1193  (
    .i0(\u_EXU_ALU/n375 ),
    .i1(\u_EXU_ALU/n383 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n407 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1194  (
    .i0(\u_EXU_ALU/n376 ),
    .i1(\u_EXU_ALU/n384 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n408 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1195  (
    .i0(\u_EXU_ALU/n377 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n409 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1196  (
    .i0(\u_EXU_ALU/n378 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n410 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1197  (
    .i0(\u_EXU_ALU/n379 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n411 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1198  (
    .i0(\u_EXU_ALU/n380 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n412 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1199  (
    .i0(\u_EXU_ALU/n381 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n413 ));  // ../RTL/core/exu_alu.v(43)
  xor \u_EXU_ALU/u12  (\u_EXU_ALU/n168 [0], i_exu_op1[0], i_exu_op2[0]);  // ../RTL/core/exu_alu.v(49)
  or \u_EXU_ALU/u120  (\u_EXU_ALU/n309 [31], \u_EXU_ALU/n308 [31], \u_EXU_ALU/alu_or [31]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1200  (
    .i0(\u_EXU_ALU/n382 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n414 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1201  (
    .i0(\u_EXU_ALU/n383 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n415 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1202  (
    .i0(\u_EXU_ALU/n384 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n416 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1203  (
    .i0(\u_EXU_ALU/n385 ),
    .i1(\u_EXU_ALU/n401 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n417 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1204  (
    .i0(\u_EXU_ALU/n386 ),
    .i1(\u_EXU_ALU/n402 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n418 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1205  (
    .i0(\u_EXU_ALU/n387 ),
    .i1(\u_EXU_ALU/n403 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n419 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1206  (
    .i0(\u_EXU_ALU/n388 ),
    .i1(\u_EXU_ALU/n404 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n420 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1207  (
    .i0(\u_EXU_ALU/n389 ),
    .i1(\u_EXU_ALU/n405 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n421 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1208  (
    .i0(\u_EXU_ALU/n390 ),
    .i1(\u_EXU_ALU/n406 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n422 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1209  (
    .i0(\u_EXU_ALU/n391 ),
    .i1(\u_EXU_ALU/n407 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n423 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u121  (\u_EXU_ALU/n308 [1], \u_EXU_ALU/n307 [1], \u_EXU_ALU/alu_and [1]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1210  (
    .i0(\u_EXU_ALU/n392 ),
    .i1(\u_EXU_ALU/n408 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n424 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1211  (
    .i0(\u_EXU_ALU/n393 ),
    .i1(\u_EXU_ALU/n409 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n425 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1212  (
    .i0(\u_EXU_ALU/n394 ),
    .i1(\u_EXU_ALU/n410 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n426 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1213  (
    .i0(\u_EXU_ALU/n395 ),
    .i1(\u_EXU_ALU/n411 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n427 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1214  (
    .i0(\u_EXU_ALU/n396 ),
    .i1(\u_EXU_ALU/n412 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n428 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1215  (
    .i0(\u_EXU_ALU/n397 ),
    .i1(\u_EXU_ALU/n413 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n429 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1216  (
    .i0(\u_EXU_ALU/n398 ),
    .i1(\u_EXU_ALU/n414 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n430 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1217  (
    .i0(\u_EXU_ALU/n399 ),
    .i1(\u_EXU_ALU/n415 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n431 ));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1218  (
    .i0(\u_EXU_ALU/n400 ),
    .i1(\u_EXU_ALU/n416 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n432 ));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u122  (\u_EXU_ALU/n308 [2], \u_EXU_ALU/n307 [2], \u_EXU_ALU/alu_and [2]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u123  (\u_EXU_ALU/n308 [3], \u_EXU_ALU/n307 [3], \u_EXU_ALU/alu_and [3]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u1235  (\u_EXU_ALU/n449 , i_exu_op2[6], i_exu_op2[7]);  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u1236  (\u_EXU_ALU/n450 , i_exu_op2[5], \u_EXU_ALU/n449 );  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u1237  (\u_EXU_ALU/n451 , i_exu_op2[9], i_exu_op2[10]);  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u1238  (\u_EXU_ALU/n452 , i_exu_op2[8], \u_EXU_ALU/n451 );  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u1239  (\u_EXU_ALU/n453 , \u_EXU_ALU/n450 , \u_EXU_ALU/n452 );  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u124  (\u_EXU_ALU/n308 [4], \u_EXU_ALU/n307 [4], \u_EXU_ALU/alu_and [4]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u1240  (\u_EXU_ALU/n454 , i_exu_op2[12], i_exu_op2[13]);  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u1241  (\u_EXU_ALU/n455 , i_exu_op2[11], \u_EXU_ALU/n454 );  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u1242  (\u_EXU_ALU/n456 , i_exu_op2[14], i_exu_op2[15]);  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u1243  (\u_EXU_ALU/n457 , i_exu_op2[16], i_exu_op2[17]);  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u1244  (\u_EXU_ALU/n458 , \u_EXU_ALU/n456 , \u_EXU_ALU/n457 );  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u1245  (\u_EXU_ALU/n459 , \u_EXU_ALU/n455 , \u_EXU_ALU/n458 );  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u1246  (\u_EXU_ALU/n460 , \u_EXU_ALU/n453 , \u_EXU_ALU/n459 );  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u1247  (\u_EXU_ALU/n461 , i_exu_op2[19], i_exu_op2[20]);  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u125  (\u_EXU_ALU/n308 [5], \u_EXU_ALU/n307 [5], \u_EXU_ALU/alu_and [5]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u126  (\u_EXU_ALU/n308 [6], \u_EXU_ALU/n307 [6], \u_EXU_ALU/alu_and [6]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1261  (
    .i0(\u_EXU_ALU/n417 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [31]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1262  (
    .i0(\u_EXU_ALU/n418 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [30]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1263  (
    .i0(\u_EXU_ALU/n419 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [29]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1264  (
    .i0(\u_EXU_ALU/n420 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [28]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1265  (
    .i0(\u_EXU_ALU/n421 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [27]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1266  (
    .i0(\u_EXU_ALU/n422 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [26]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1267  (
    .i0(\u_EXU_ALU/n423 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [25]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1268  (
    .i0(\u_EXU_ALU/n424 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [24]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1269  (
    .i0(\u_EXU_ALU/n425 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [23]));  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u127  (\u_EXU_ALU/n308 [7], \u_EXU_ALU/n307 [7], \u_EXU_ALU/alu_and [7]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1270  (
    .i0(\u_EXU_ALU/n426 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [22]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1271  (
    .i0(\u_EXU_ALU/n427 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [21]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1272  (
    .i0(\u_EXU_ALU/n428 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [20]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1273  (
    .i0(\u_EXU_ALU/n429 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [19]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1274  (
    .i0(\u_EXU_ALU/n430 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [18]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1275  (
    .i0(\u_EXU_ALU/n431 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [17]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1276  (
    .i0(\u_EXU_ALU/n432 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n281 ),
    .o(\u_EXU_ALU/n66 [16]));  // ../RTL/core/exu_alu.v(43)
  AL_MUX \u_EXU_ALU/u1277  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n401 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [15]));
  AL_MUX \u_EXU_ALU/u1278  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n402 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [14]));
  AL_MUX \u_EXU_ALU/u1279  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n403 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [13]));
  or \u_EXU_ALU/u128  (\u_EXU_ALU/n308 [8], \u_EXU_ALU/n307 [8], \u_EXU_ALU/alu_and [8]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1280  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n404 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [12]));
  AL_MUX \u_EXU_ALU/u1281  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n405 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [11]));
  AL_MUX \u_EXU_ALU/u1282  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n406 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [10]));
  AL_MUX \u_EXU_ALU/u1283  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n407 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [9]));
  AL_MUX \u_EXU_ALU/u1284  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n408 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [8]));
  AL_MUX \u_EXU_ALU/u1285  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n409 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [7]));
  AL_MUX \u_EXU_ALU/u1286  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n410 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [6]));
  AL_MUX \u_EXU_ALU/u1287  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n411 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [5]));
  AL_MUX \u_EXU_ALU/u1288  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n412 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [4]));
  AL_MUX \u_EXU_ALU/u1289  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n413 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [3]));
  or \u_EXU_ALU/u129  (\u_EXU_ALU/n308 [9], \u_EXU_ALU/n307 [9], \u_EXU_ALU/alu_and [9]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u1290  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n414 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [2]));
  AL_MUX \u_EXU_ALU/u1291  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n415 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [1]));
  AL_MUX \u_EXU_ALU/u1292  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n416 ),
    .sel(\u_EXU_ALU/u1029_sel_is_0_o ),
    .o(\u_EXU_ALU/n66 [0]));
  and \u_EXU_ALU/u1293  (\u_EXU_ALU/alu_sub [1], i_decinfo[1], \u_EXU_ALU/n33 [1]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1294  (\u_EXU_ALU/alu_sub [2], i_decinfo[1], \u_EXU_ALU/n33 [2]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1295  (\u_EXU_ALU/alu_sub [3], i_decinfo[1], \u_EXU_ALU/n33 [3]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1296  (\u_EXU_ALU/alu_sub [4], i_decinfo[1], \u_EXU_ALU/n33 [4]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1297  (\u_EXU_ALU/alu_sub [5], i_decinfo[1], \u_EXU_ALU/n33 [5]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1298  (\u_EXU_ALU/alu_sub [6], i_decinfo[1], \u_EXU_ALU/n33 [6]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1299  (\u_EXU_ALU/alu_sub [7], i_decinfo[1], \u_EXU_ALU/n33 [7]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u13  (\u_EXU_ALU/alu_xor [0], i_decinfo[5], \u_EXU_ALU/n168 [0]);  // ../RTL/core/exu_alu.v(49)
  or \u_EXU_ALU/u130  (\u_EXU_ALU/n308 [10], \u_EXU_ALU/n307 [10], \u_EXU_ALU/alu_and [10]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u1300  (\u_EXU_ALU/alu_sub [8], i_decinfo[1], \u_EXU_ALU/n33 [8]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1301  (\u_EXU_ALU/alu_sub [9], i_decinfo[1], \u_EXU_ALU/n33 [9]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1302  (\u_EXU_ALU/alu_sub [10], i_decinfo[1], \u_EXU_ALU/n33 [10]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1303  (\u_EXU_ALU/alu_sub [11], i_decinfo[1], \u_EXU_ALU/n33 [11]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1304  (\u_EXU_ALU/alu_sub [12], i_decinfo[1], \u_EXU_ALU/n33 [12]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1305  (\u_EXU_ALU/alu_sub [13], i_decinfo[1], \u_EXU_ALU/n33 [13]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1306  (\u_EXU_ALU/alu_sub [14], i_decinfo[1], \u_EXU_ALU/n33 [14]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1307  (\u_EXU_ALU/alu_sub [15], i_decinfo[1], \u_EXU_ALU/n33 [15]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1308  (\u_EXU_ALU/alu_sub [16], i_decinfo[1], \u_EXU_ALU/n33 [16]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1309  (\u_EXU_ALU/alu_sub [17], i_decinfo[1], \u_EXU_ALU/n33 [17]);  // ../RTL/core/exu_alu.v(41)
  or \u_EXU_ALU/u131  (\u_EXU_ALU/n308 [11], \u_EXU_ALU/n307 [11], \u_EXU_ALU/alu_and [11]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u1310  (\u_EXU_ALU/alu_sub [18], i_decinfo[1], \u_EXU_ALU/n33 [18]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1311  (\u_EXU_ALU/alu_sub [19], i_decinfo[1], \u_EXU_ALU/n33 [19]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1312  (\u_EXU_ALU/alu_sub [20], i_decinfo[1], \u_EXU_ALU/n33 [20]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1313  (\u_EXU_ALU/alu_sub [21], i_decinfo[1], \u_EXU_ALU/n33 [21]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1314  (\u_EXU_ALU/alu_sub [22], i_decinfo[1], \u_EXU_ALU/n33 [22]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1315  (\u_EXU_ALU/alu_sub [23], i_decinfo[1], \u_EXU_ALU/n33 [23]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1316  (\u_EXU_ALU/alu_sub [24], i_decinfo[1], \u_EXU_ALU/n33 [24]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1317  (\u_EXU_ALU/alu_sub [25], i_decinfo[1], \u_EXU_ALU/n33 [25]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1318  (\u_EXU_ALU/alu_sub [26], i_decinfo[1], \u_EXU_ALU/n33 [26]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1319  (\u_EXU_ALU/alu_sub [27], i_decinfo[1], \u_EXU_ALU/n33 [27]);  // ../RTL/core/exu_alu.v(41)
  or \u_EXU_ALU/u132  (\u_EXU_ALU/n308 [12], \u_EXU_ALU/n307 [12], \u_EXU_ALU/alu_and [12]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u1320  (\u_EXU_ALU/alu_sub [28], i_decinfo[1], \u_EXU_ALU/n33 [28]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1321  (\u_EXU_ALU/alu_sub [29], i_decinfo[1], \u_EXU_ALU/n33 [29]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1322  (\u_EXU_ALU/alu_sub [30], i_decinfo[1], \u_EXU_ALU/n33 [30]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1323  (\u_EXU_ALU/alu_sub [31], i_decinfo[1], \u_EXU_ALU/n33 [31]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u1324  (alu2lsu_result[1], i_decinfo_grp[5], \u_EXU_ALU/n0 [1]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1325  (alu2lsu_result[2], i_decinfo_grp[5], \u_EXU_ALU/n0 [2]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1326  (alu2lsu_result[3], i_decinfo_grp[5], \u_EXU_ALU/n0 [3]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1327  (alu2lsu_result[4], i_decinfo_grp[5], \u_EXU_ALU/n0 [4]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1328  (alu2lsu_result[5], i_decinfo_grp[5], \u_EXU_ALU/n0 [5]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1329  (alu2lsu_result[6], i_decinfo_grp[5], \u_EXU_ALU/n0 [6]);  // ../RTL/core/exu_alu.v(39)
  or \u_EXU_ALU/u133  (\u_EXU_ALU/n308 [13], \u_EXU_ALU/n307 [13], \u_EXU_ALU/alu_and [13]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u1330  (alu2lsu_result[7], i_decinfo_grp[5], \u_EXU_ALU/n0 [7]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1331  (alu2lsu_result[8], i_decinfo_grp[5], \u_EXU_ALU/n0 [8]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1332  (alu2lsu_result[9], i_decinfo_grp[5], \u_EXU_ALU/n0 [9]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1333  (alu2lsu_result[10], i_decinfo_grp[5], \u_EXU_ALU/n0 [10]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1334  (alu2lsu_result[11], i_decinfo_grp[5], \u_EXU_ALU/n0 [11]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1335  (alu2lsu_result[12], i_decinfo_grp[5], \u_EXU_ALU/n0 [12]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1336  (alu2lsu_result[13], i_decinfo_grp[5], \u_EXU_ALU/n0 [13]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1337  (alu2lsu_result[14], i_decinfo_grp[5], \u_EXU_ALU/n0 [14]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1338  (alu2lsu_result[15], i_decinfo_grp[5], \u_EXU_ALU/n0 [15]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1339  (alu2lsu_result[16], i_decinfo_grp[5], \u_EXU_ALU/n0 [16]);  // ../RTL/core/exu_alu.v(39)
  or \u_EXU_ALU/u134  (\u_EXU_ALU/n308 [14], \u_EXU_ALU/n307 [14], \u_EXU_ALU/alu_and [14]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u1340  (alu2lsu_result[17], i_decinfo_grp[5], \u_EXU_ALU/n0 [17]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1341  (alu2lsu_result[18], i_decinfo_grp[5], \u_EXU_ALU/n0 [18]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1342  (alu2lsu_result[19], i_decinfo_grp[5], \u_EXU_ALU/n0 [19]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1343  (alu2lsu_result[20], i_decinfo_grp[5], \u_EXU_ALU/n0 [20]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1344  (alu2lsu_result[21], i_decinfo_grp[5], \u_EXU_ALU/n0 [21]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1345  (alu2lsu_result[22], i_decinfo_grp[5], \u_EXU_ALU/n0 [22]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1346  (alu2lsu_result[23], i_decinfo_grp[5], \u_EXU_ALU/n0 [23]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1347  (alu2lsu_result[24], i_decinfo_grp[5], \u_EXU_ALU/n0 [24]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1348  (alu2lsu_result[25], i_decinfo_grp[5], \u_EXU_ALU/n0 [25]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1349  (alu2lsu_result[26], i_decinfo_grp[5], \u_EXU_ALU/n0 [26]);  // ../RTL/core/exu_alu.v(39)
  or \u_EXU_ALU/u135  (\u_EXU_ALU/n308 [15], \u_EXU_ALU/n307 [15], \u_EXU_ALU/alu_and [15]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u1350  (alu2lsu_result[27], i_decinfo_grp[5], \u_EXU_ALU/n0 [27]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1351  (alu2lsu_result[28], i_decinfo_grp[5], \u_EXU_ALU/n0 [28]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1352  (alu2lsu_result[29], i_decinfo_grp[5], \u_EXU_ALU/n0 [29]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1353  (alu2lsu_result[30], i_decinfo_grp[5], \u_EXU_ALU/n0 [30]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u1354  (alu2lsu_result[31], i_decinfo_grp[5], \u_EXU_ALU/n0 [31]);  // ../RTL/core/exu_alu.v(39)
  or \u_EXU_ALU/u136  (\u_EXU_ALU/n308 [16], \u_EXU_ALU/n307 [16], \u_EXU_ALU/alu_and [16]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u137  (\u_EXU_ALU/n308 [17], \u_EXU_ALU/n307 [17], \u_EXU_ALU/alu_and [17]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u138  (\u_EXU_ALU/n308 [18], \u_EXU_ALU/n307 [18], \u_EXU_ALU/alu_and [18]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u139  (\u_EXU_ALU/n308 [19], \u_EXU_ALU/n307 [19], \u_EXU_ALU/alu_and [19]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u14  (\u_EXU_ALU/n201 [0], i_exu_op1[0], i_exu_op2[0]);  // ../RTL/core/exu_alu.v(51)
  or \u_EXU_ALU/u140  (\u_EXU_ALU/n308 [20], \u_EXU_ALU/n307 [20], \u_EXU_ALU/alu_and [20]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u141  (\u_EXU_ALU/n308 [21], \u_EXU_ALU/n307 [21], \u_EXU_ALU/alu_and [21]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u142  (\u_EXU_ALU/n308 [22], \u_EXU_ALU/n307 [22], \u_EXU_ALU/alu_and [22]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u143  (\u_EXU_ALU/n308 [23], \u_EXU_ALU/n307 [23], \u_EXU_ALU/alu_and [23]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u144  (\u_EXU_ALU/n308 [24], \u_EXU_ALU/n307 [24], \u_EXU_ALU/alu_and [24]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u145  (\u_EXU_ALU/n308 [25], \u_EXU_ALU/n307 [25], \u_EXU_ALU/alu_and [25]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u146  (\u_EXU_ALU/n308 [26], \u_EXU_ALU/n307 [26], \u_EXU_ALU/alu_and [26]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u147  (\u_EXU_ALU/n308 [27], \u_EXU_ALU/n307 [27], \u_EXU_ALU/alu_and [27]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u148  (\u_EXU_ALU/n308 [28], \u_EXU_ALU/n307 [28], \u_EXU_ALU/alu_and [28]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u149  (\u_EXU_ALU/n308 [29], \u_EXU_ALU/n307 [29], \u_EXU_ALU/alu_and [29]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u15  (\u_EXU_ALU/alu_and [0], i_decinfo[6], \u_EXU_ALU/n201 [0]);  // ../RTL/core/exu_alu.v(51)
  or \u_EXU_ALU/u150  (\u_EXU_ALU/n308 [30], \u_EXU_ALU/n307 [30], \u_EXU_ALU/alu_and [30]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u151  (\u_EXU_ALU/n308 [31], \u_EXU_ALU/n307 [31], \u_EXU_ALU/alu_and [31]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u152  (\u_EXU_ALU/n307 [1], \u_EXU_ALU/n306 [1], \u_EXU_ALU/alu_xor [1]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u153  (\u_EXU_ALU/n307 [2], \u_EXU_ALU/n306 [2], \u_EXU_ALU/alu_xor [2]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u154  (\u_EXU_ALU/n307 [3], \u_EXU_ALU/n306 [3], \u_EXU_ALU/alu_xor [3]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u155  (\u_EXU_ALU/n307 [4], \u_EXU_ALU/n306 [4], \u_EXU_ALU/alu_xor [4]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u156  (\u_EXU_ALU/n307 [5], \u_EXU_ALU/n306 [5], \u_EXU_ALU/alu_xor [5]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u157  (\u_EXU_ALU/n307 [6], \u_EXU_ALU/n306 [6], \u_EXU_ALU/alu_xor [6]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u158  (\u_EXU_ALU/n307 [7], \u_EXU_ALU/n306 [7], \u_EXU_ALU/alu_xor [7]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u159  (\u_EXU_ALU/n307 [8], \u_EXU_ALU/n306 [8], \u_EXU_ALU/alu_xor [8]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u16  (\u_EXU_ALU/n233 [0], i_exu_op1[0], i_exu_op2[0]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u160  (\u_EXU_ALU/n307 [9], \u_EXU_ALU/n306 [9], \u_EXU_ALU/alu_xor [9]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u161  (\u_EXU_ALU/n307 [10], \u_EXU_ALU/n306 [10], \u_EXU_ALU/alu_xor [10]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u162  (\u_EXU_ALU/n307 [11], \u_EXU_ALU/n306 [11], \u_EXU_ALU/alu_xor [11]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u163  (\u_EXU_ALU/n307 [12], \u_EXU_ALU/n306 [12], \u_EXU_ALU/alu_xor [12]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u164  (\u_EXU_ALU/n307 [13], \u_EXU_ALU/n306 [13], \u_EXU_ALU/alu_xor [13]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u165  (\u_EXU_ALU/n307 [14], \u_EXU_ALU/n306 [14], \u_EXU_ALU/alu_xor [14]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u166  (\u_EXU_ALU/n307 [15], \u_EXU_ALU/n306 [15], \u_EXU_ALU/alu_xor [15]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u167  (\u_EXU_ALU/n307 [16], \u_EXU_ALU/n306 [16], \u_EXU_ALU/alu_xor [16]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u168  (\u_EXU_ALU/n307 [17], \u_EXU_ALU/n306 [17], \u_EXU_ALU/alu_xor [17]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u169  (\u_EXU_ALU/n307 [18], \u_EXU_ALU/n306 [18], \u_EXU_ALU/alu_xor [18]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u17  (\u_EXU_ALU/alu_or [0], i_decinfo[7], \u_EXU_ALU/n233 [0]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u170  (\u_EXU_ALU/n307 [19], \u_EXU_ALU/n306 [19], \u_EXU_ALU/alu_xor [19]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u171  (\u_EXU_ALU/n307 [20], \u_EXU_ALU/n306 [20], \u_EXU_ALU/alu_xor [20]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u172  (\u_EXU_ALU/n307 [21], \u_EXU_ALU/n306 [21], \u_EXU_ALU/alu_xor [21]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u173  (\u_EXU_ALU/n307 [22], \u_EXU_ALU/n306 [22], \u_EXU_ALU/alu_xor [22]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u174  (\u_EXU_ALU/n307 [23], \u_EXU_ALU/n306 [23], \u_EXU_ALU/alu_xor [23]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u175  (\u_EXU_ALU/n307 [24], \u_EXU_ALU/n306 [24], \u_EXU_ALU/alu_xor [24]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u176  (\u_EXU_ALU/n307 [25], \u_EXU_ALU/n306 [25], \u_EXU_ALU/alu_xor [25]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u177  (\u_EXU_ALU/n307 [26], \u_EXU_ALU/n306 [26], \u_EXU_ALU/alu_xor [26]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u178  (\u_EXU_ALU/n307 [27], \u_EXU_ALU/n306 [27], \u_EXU_ALU/alu_xor [27]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u179  (\u_EXU_ALU/n307 [28], \u_EXU_ALU/n306 [28], \u_EXU_ALU/alu_xor [28]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u18  (\u_EXU_ALU/alu_slt [0], i_decinfo[8], \u_EXU_ALU/n253 );  // ../RTL/core/exu_alu.v(55)
  or \u_EXU_ALU/u180  (\u_EXU_ALU/n307 [29], \u_EXU_ALU/n306 [29], \u_EXU_ALU/alu_xor [29]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u181  (\u_EXU_ALU/n307 [30], \u_EXU_ALU/n306 [30], \u_EXU_ALU/alu_xor [30]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u182  (\u_EXU_ALU/n307 [31], \u_EXU_ALU/n306 [31], \u_EXU_ALU/alu_xor [31]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u183  (\u_EXU_ALU/n306 [1], \u_EXU_ALU/n305 [1], \u_EXU_ALU/alu_sra [1]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u184  (\u_EXU_ALU/n306 [2], \u_EXU_ALU/n305 [2], \u_EXU_ALU/alu_sra [2]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u185  (\u_EXU_ALU/n306 [3], \u_EXU_ALU/n305 [3], \u_EXU_ALU/alu_sra [3]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u186  (\u_EXU_ALU/n306 [4], \u_EXU_ALU/n305 [4], \u_EXU_ALU/alu_sra [4]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u187  (\u_EXU_ALU/n306 [5], \u_EXU_ALU/n305 [5], \u_EXU_ALU/alu_sra [5]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u188  (\u_EXU_ALU/n306 [6], \u_EXU_ALU/n305 [6], \u_EXU_ALU/alu_sra [6]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u189  (\u_EXU_ALU/n306 [7], \u_EXU_ALU/n305 [7], \u_EXU_ALU/alu_sra [7]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u19  (\u_EXU_ALU/alu_sltu [0], i_decinfo[9], \u_EXU_ALU/n261 );  // ../RTL/core/exu_alu.v(57)
  or \u_EXU_ALU/u190  (\u_EXU_ALU/n306 [8], \u_EXU_ALU/n305 [8], \u_EXU_ALU/alu_sra [8]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u191  (\u_EXU_ALU/n306 [9], \u_EXU_ALU/n305 [9], \u_EXU_ALU/alu_sra [9]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u192  (\u_EXU_ALU/n306 [10], \u_EXU_ALU/n305 [10], \u_EXU_ALU/alu_sra [10]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u193  (\u_EXU_ALU/n306 [11], \u_EXU_ALU/n305 [11], \u_EXU_ALU/alu_sra [11]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u194  (\u_EXU_ALU/n306 [12], \u_EXU_ALU/n305 [12], \u_EXU_ALU/alu_sra [12]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u195  (\u_EXU_ALU/n306 [13], \u_EXU_ALU/n305 [13], \u_EXU_ALU/alu_sra [13]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u196  (\u_EXU_ALU/n306 [14], \u_EXU_ALU/n305 [14], \u_EXU_ALU/alu_sra [14]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u197  (\u_EXU_ALU/n306 [15], \u_EXU_ALU/n305 [15], \u_EXU_ALU/alu_sra [15]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u198  (\u_EXU_ALU/n306 [16], \u_EXU_ALU/n305 [16], \u_EXU_ALU/alu_sra [16]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u199  (\u_EXU_ALU/n306 [17], \u_EXU_ALU/n305 [17], \u_EXU_ALU/alu_sra [17]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u200  (\u_EXU_ALU/n306 [18], \u_EXU_ALU/n305 [18], \u_EXU_ALU/alu_sra [18]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u201  (\u_EXU_ALU/n306 [19], \u_EXU_ALU/n305 [19], \u_EXU_ALU/alu_sra [19]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u202  (\u_EXU_ALU/n306 [20], \u_EXU_ALU/n305 [20], \u_EXU_ALU/alu_sra [20]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u203  (\u_EXU_ALU/n306 [21], \u_EXU_ALU/n305 [21], \u_EXU_ALU/alu_sra [21]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u204  (\u_EXU_ALU/n306 [22], \u_EXU_ALU/n305 [22], \u_EXU_ALU/alu_sra [22]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u205  (\u_EXU_ALU/n306 [23], \u_EXU_ALU/n305 [23], \u_EXU_ALU/alu_sra [23]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u206  (\u_EXU_ALU/n306 [24], \u_EXU_ALU/n305 [24], \u_EXU_ALU/alu_sra [24]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u207  (\u_EXU_ALU/n306 [25], \u_EXU_ALU/n305 [25], \u_EXU_ALU/alu_sra [25]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u208  (\u_EXU_ALU/n306 [26], \u_EXU_ALU/n305 [26], \u_EXU_ALU/alu_sra [26]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u209  (\u_EXU_ALU/n306 [27], \u_EXU_ALU/n305 [27], \u_EXU_ALU/alu_sra [27]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u210  (\u_EXU_ALU/n306 [28], \u_EXU_ALU/n305 [28], \u_EXU_ALU/alu_sra [28]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u211  (\u_EXU_ALU/n306 [29], \u_EXU_ALU/n305 [29], \u_EXU_ALU/alu_sra [29]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u212  (\u_EXU_ALU/n306 [30], \u_EXU_ALU/n305 [30], \u_EXU_ALU/alu_sra [30]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u213  (\u_EXU_ALU/n306 [31], \u_EXU_ALU/n305 [31], \u_EXU_ALU/alu_sra [31]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u214  (\u_EXU_ALU/n305 [1], \u_EXU_ALU/n304 [1], \u_EXU_ALU/alu_srl [1]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u215  (\u_EXU_ALU/n305 [2], \u_EXU_ALU/n304 [2], \u_EXU_ALU/alu_srl [2]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u216  (\u_EXU_ALU/n305 [3], \u_EXU_ALU/n304 [3], \u_EXU_ALU/alu_srl [3]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u217  (\u_EXU_ALU/n305 [4], \u_EXU_ALU/n304 [4], \u_EXU_ALU/alu_srl [4]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u218  (\u_EXU_ALU/n305 [5], \u_EXU_ALU/n304 [5], \u_EXU_ALU/alu_srl [5]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u219  (\u_EXU_ALU/n305 [6], \u_EXU_ALU/n304 [6], \u_EXU_ALU/alu_srl [6]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u220  (\u_EXU_ALU/n305 [7], \u_EXU_ALU/n304 [7], \u_EXU_ALU/alu_srl [7]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u221  (\u_EXU_ALU/n305 [8], \u_EXU_ALU/n304 [8], \u_EXU_ALU/alu_srl [8]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u222  (\u_EXU_ALU/n305 [9], \u_EXU_ALU/n304 [9], \u_EXU_ALU/alu_srl [9]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u223  (\u_EXU_ALU/n305 [10], \u_EXU_ALU/n304 [10], \u_EXU_ALU/alu_srl [10]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u224  (\u_EXU_ALU/n305 [11], \u_EXU_ALU/n304 [11], \u_EXU_ALU/alu_srl [11]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u225  (\u_EXU_ALU/n305 [12], \u_EXU_ALU/n304 [12], \u_EXU_ALU/alu_srl [12]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u226  (\u_EXU_ALU/n305 [13], \u_EXU_ALU/n304 [13], \u_EXU_ALU/alu_srl [13]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u227  (\u_EXU_ALU/n305 [14], \u_EXU_ALU/n304 [14], \u_EXU_ALU/alu_srl [14]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u228  (\u_EXU_ALU/n305 [15], \u_EXU_ALU/n304 [15], \u_EXU_ALU/alu_srl [15]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u229  (\u_EXU_ALU/n305 [16], \u_EXU_ALU/n304 [16], \u_EXU_ALU/alu_srl [16]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u23  (\u_EXU_ALU/n303 [0], alu2lsu_result[0], \u_EXU_ALU/alu_sub [0]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u230  (\u_EXU_ALU/n305 [17], \u_EXU_ALU/n304 [17], \u_EXU_ALU/alu_srl [17]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u231  (\u_EXU_ALU/n305 [18], \u_EXU_ALU/n304 [18], \u_EXU_ALU/alu_srl [18]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u232  (\u_EXU_ALU/n305 [19], \u_EXU_ALU/n304 [19], \u_EXU_ALU/alu_srl [19]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u233  (\u_EXU_ALU/n305 [20], \u_EXU_ALU/n304 [20], \u_EXU_ALU/alu_srl [20]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u234  (\u_EXU_ALU/n305 [21], \u_EXU_ALU/n304 [21], \u_EXU_ALU/alu_srl [21]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u235  (\u_EXU_ALU/n305 [22], \u_EXU_ALU/n304 [22], \u_EXU_ALU/alu_srl [22]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u236  (\u_EXU_ALU/n305 [23], \u_EXU_ALU/n304 [23], \u_EXU_ALU/alu_srl [23]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u237  (\u_EXU_ALU/n305 [24], \u_EXU_ALU/n304 [24], \u_EXU_ALU/alu_srl [24]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u238  (\u_EXU_ALU/n305 [25], \u_EXU_ALU/n304 [25], \u_EXU_ALU/alu_srl [25]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u239  (\u_EXU_ALU/n305 [26], \u_EXU_ALU/n304 [26], \u_EXU_ALU/alu_srl [26]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u24  (\u_EXU_ALU/n304 [0], \u_EXU_ALU/n303 [0], \u_EXU_ALU/alu_sll [0]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u240  (\u_EXU_ALU/n305 [27], \u_EXU_ALU/n304 [27], \u_EXU_ALU/alu_srl [27]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u241  (\u_EXU_ALU/n305 [28], \u_EXU_ALU/n304 [28], \u_EXU_ALU/alu_srl [28]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u242  (\u_EXU_ALU/n305 [29], \u_EXU_ALU/n304 [29], \u_EXU_ALU/alu_srl [29]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u243  (\u_EXU_ALU/n305 [30], \u_EXU_ALU/n304 [30], \u_EXU_ALU/alu_srl [30]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u244  (\u_EXU_ALU/n305 [31], \u_EXU_ALU/n304 [31], \u_EXU_ALU/alu_srl [31]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u245  (\u_EXU_ALU/n304 [1], \u_EXU_ALU/n303 [1], \u_EXU_ALU/alu_sll [1]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u246  (\u_EXU_ALU/n304 [2], \u_EXU_ALU/n303 [2], \u_EXU_ALU/alu_sll [2]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u247  (\u_EXU_ALU/n304 [3], \u_EXU_ALU/n303 [3], \u_EXU_ALU/alu_sll [3]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u248  (\u_EXU_ALU/n304 [4], \u_EXU_ALU/n303 [4], \u_EXU_ALU/alu_sll [4]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u249  (\u_EXU_ALU/n304 [5], \u_EXU_ALU/n303 [5], \u_EXU_ALU/alu_sll [5]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u25  (\u_EXU_ALU/n305 [0], \u_EXU_ALU/n304 [0], \u_EXU_ALU/alu_srl [0]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u250  (\u_EXU_ALU/n304 [6], \u_EXU_ALU/n303 [6], \u_EXU_ALU/alu_sll [6]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u251  (\u_EXU_ALU/n304 [7], \u_EXU_ALU/n303 [7], \u_EXU_ALU/alu_sll [7]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u252  (\u_EXU_ALU/n304 [8], \u_EXU_ALU/n303 [8], \u_EXU_ALU/alu_sll [8]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u253  (\u_EXU_ALU/n304 [9], \u_EXU_ALU/n303 [9], \u_EXU_ALU/alu_sll [9]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u254  (\u_EXU_ALU/n304 [10], \u_EXU_ALU/n303 [10], \u_EXU_ALU/alu_sll [10]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u255  (\u_EXU_ALU/n304 [11], \u_EXU_ALU/n303 [11], \u_EXU_ALU/alu_sll [11]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u256  (\u_EXU_ALU/n304 [12], \u_EXU_ALU/n303 [12], \u_EXU_ALU/alu_sll [12]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u257  (\u_EXU_ALU/n304 [13], \u_EXU_ALU/n303 [13], \u_EXU_ALU/alu_sll [13]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u258  (\u_EXU_ALU/n304 [14], \u_EXU_ALU/n303 [14], \u_EXU_ALU/alu_sll [14]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u259  (\u_EXU_ALU/n304 [15], \u_EXU_ALU/n303 [15], \u_EXU_ALU/alu_sll [15]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u26  (\u_EXU_ALU/n306 [0], \u_EXU_ALU/n305 [0], \u_EXU_ALU/alu_sra [0]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u260  (\u_EXU_ALU/n304 [16], \u_EXU_ALU/n303 [16], \u_EXU_ALU/alu_sll [16]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u261  (\u_EXU_ALU/n304 [17], \u_EXU_ALU/n303 [17], \u_EXU_ALU/alu_sll [17]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u262  (\u_EXU_ALU/n304 [18], \u_EXU_ALU/n303 [18], \u_EXU_ALU/alu_sll [18]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u263  (\u_EXU_ALU/n304 [19], \u_EXU_ALU/n303 [19], \u_EXU_ALU/alu_sll [19]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u264  (\u_EXU_ALU/n304 [20], \u_EXU_ALU/n303 [20], \u_EXU_ALU/alu_sll [20]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u265  (\u_EXU_ALU/n304 [21], \u_EXU_ALU/n303 [21], \u_EXU_ALU/alu_sll [21]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u266  (\u_EXU_ALU/n304 [22], \u_EXU_ALU/n303 [22], \u_EXU_ALU/alu_sll [22]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u267  (\u_EXU_ALU/n304 [23], \u_EXU_ALU/n303 [23], \u_EXU_ALU/alu_sll [23]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u268  (\u_EXU_ALU/n304 [24], \u_EXU_ALU/n303 [24], \u_EXU_ALU/alu_sll [24]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u269  (\u_EXU_ALU/n304 [25], \u_EXU_ALU/n303 [25], \u_EXU_ALU/alu_sll [25]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u27  (\u_EXU_ALU/n307 [0], \u_EXU_ALU/n306 [0], \u_EXU_ALU/alu_xor [0]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u270  (\u_EXU_ALU/n304 [26], \u_EXU_ALU/n303 [26], \u_EXU_ALU/alu_sll [26]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u271  (\u_EXU_ALU/n304 [27], \u_EXU_ALU/n303 [27], \u_EXU_ALU/alu_sll [27]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u272  (\u_EXU_ALU/n304 [28], \u_EXU_ALU/n303 [28], \u_EXU_ALU/alu_sll [28]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u273  (\u_EXU_ALU/n304 [29], \u_EXU_ALU/n303 [29], \u_EXU_ALU/alu_sll [29]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u274  (\u_EXU_ALU/n304 [30], \u_EXU_ALU/n303 [30], \u_EXU_ALU/alu_sll [30]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u275  (\u_EXU_ALU/n304 [31], \u_EXU_ALU/n303 [31], \u_EXU_ALU/alu_sll [31]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u276  (\u_EXU_ALU/n303 [1], alu2lsu_result[1], \u_EXU_ALU/alu_sub [1]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u277  (\u_EXU_ALU/n303 [2], alu2lsu_result[2], \u_EXU_ALU/alu_sub [2]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u278  (\u_EXU_ALU/n303 [3], alu2lsu_result[3], \u_EXU_ALU/alu_sub [3]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u279  (\u_EXU_ALU/n303 [4], alu2lsu_result[4], \u_EXU_ALU/alu_sub [4]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u28  (\u_EXU_ALU/n308 [0], \u_EXU_ALU/n307 [0], \u_EXU_ALU/alu_and [0]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u280  (\u_EXU_ALU/n303 [5], alu2lsu_result[5], \u_EXU_ALU/alu_sub [5]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u281  (\u_EXU_ALU/n303 [6], alu2lsu_result[6], \u_EXU_ALU/alu_sub [6]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u282  (\u_EXU_ALU/n303 [7], alu2lsu_result[7], \u_EXU_ALU/alu_sub [7]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u283  (\u_EXU_ALU/n303 [8], alu2lsu_result[8], \u_EXU_ALU/alu_sub [8]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u284  (\u_EXU_ALU/n303 [9], alu2lsu_result[9], \u_EXU_ALU/alu_sub [9]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u285  (\u_EXU_ALU/n303 [10], alu2lsu_result[10], \u_EXU_ALU/alu_sub [10]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u286  (\u_EXU_ALU/n303 [11], alu2lsu_result[11], \u_EXU_ALU/alu_sub [11]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u287  (\u_EXU_ALU/n303 [12], alu2lsu_result[12], \u_EXU_ALU/alu_sub [12]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u288  (\u_EXU_ALU/n303 [13], alu2lsu_result[13], \u_EXU_ALU/alu_sub [13]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u289  (\u_EXU_ALU/n303 [14], alu2lsu_result[14], \u_EXU_ALU/alu_sub [14]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u29  (\u_EXU_ALU/n309 [0], \u_EXU_ALU/n308 [0], \u_EXU_ALU/alu_or [0]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u290  (\u_EXU_ALU/n303 [15], alu2lsu_result[15], \u_EXU_ALU/alu_sub [15]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u291  (\u_EXU_ALU/n303 [16], alu2lsu_result[16], \u_EXU_ALU/alu_sub [16]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u292  (\u_EXU_ALU/n303 [17], alu2lsu_result[17], \u_EXU_ALU/alu_sub [17]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u293  (\u_EXU_ALU/n303 [18], alu2lsu_result[18], \u_EXU_ALU/alu_sub [18]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u294  (\u_EXU_ALU/n303 [19], alu2lsu_result[19], \u_EXU_ALU/alu_sub [19]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u295  (\u_EXU_ALU/n303 [20], alu2lsu_result[20], \u_EXU_ALU/alu_sub [20]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u296  (\u_EXU_ALU/n303 [21], alu2lsu_result[21], \u_EXU_ALU/alu_sub [21]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u297  (\u_EXU_ALU/n303 [22], alu2lsu_result[22], \u_EXU_ALU/alu_sub [22]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u298  (\u_EXU_ALU/n303 [23], alu2lsu_result[23], \u_EXU_ALU/alu_sub [23]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u299  (\u_EXU_ALU/n303 [24], alu2lsu_result[24], \u_EXU_ALU/alu_sub [24]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u30  (\u_EXU_ALU/n310 [0], \u_EXU_ALU/n309 [0], \u_EXU_ALU/alu_slt [0]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u300  (\u_EXU_ALU/n303 [25], alu2lsu_result[25], \u_EXU_ALU/alu_sub [25]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u301  (\u_EXU_ALU/n303 [26], alu2lsu_result[26], \u_EXU_ALU/alu_sub [26]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u302  (\u_EXU_ALU/n303 [27], alu2lsu_result[27], \u_EXU_ALU/alu_sub [27]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u303  (\u_EXU_ALU/n303 [28], alu2lsu_result[28], \u_EXU_ALU/alu_sub [28]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u304  (\u_EXU_ALU/n303 [29], alu2lsu_result[29], \u_EXU_ALU/alu_sub [29]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u305  (\u_EXU_ALU/n303 [30], alu2lsu_result[30], \u_EXU_ALU/alu_sub [30]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u306  (\u_EXU_ALU/n303 [31], alu2lsu_result[31], \u_EXU_ALU/alu_sub [31]);  // ../RTL/core/exu_alu.v(66)
  and \u_EXU_ALU/u4  (alu2lsu_result[0], i_decinfo_grp[5], \u_EXU_ALU/n0 [0]);  // ../RTL/core/exu_alu.v(39)
  and \u_EXU_ALU/u404  (\u_EXU_ALU/alu_or [1], i_decinfo[7], \u_EXU_ALU/n233 [1]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u405  (\u_EXU_ALU/alu_or [2], i_decinfo[7], \u_EXU_ALU/n233 [2]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u406  (\u_EXU_ALU/alu_or [3], i_decinfo[7], \u_EXU_ALU/n233 [3]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u407  (\u_EXU_ALU/alu_or [4], i_decinfo[7], \u_EXU_ALU/n233 [4]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u408  (\u_EXU_ALU/alu_or [5], i_decinfo[7], \u_EXU_ALU/n233 [5]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u409  (\u_EXU_ALU/alu_or [6], i_decinfo[7], \u_EXU_ALU/n233 [6]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u410  (\u_EXU_ALU/alu_or [7], i_decinfo[7], \u_EXU_ALU/n233 [7]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u411  (\u_EXU_ALU/alu_or [8], i_decinfo[7], \u_EXU_ALU/n233 [8]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u412  (\u_EXU_ALU/alu_or [9], i_decinfo[7], \u_EXU_ALU/n233 [9]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u413  (\u_EXU_ALU/alu_or [10], i_decinfo[7], \u_EXU_ALU/n233 [10]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u414  (\u_EXU_ALU/alu_or [11], i_decinfo[7], \u_EXU_ALU/n233 [11]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u415  (\u_EXU_ALU/alu_or [12], i_decinfo[7], \u_EXU_ALU/n233 [12]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u416  (\u_EXU_ALU/alu_or [13], i_decinfo[7], \u_EXU_ALU/n233 [13]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u417  (\u_EXU_ALU/alu_or [14], i_decinfo[7], \u_EXU_ALU/n233 [14]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u418  (\u_EXU_ALU/alu_or [15], i_decinfo[7], \u_EXU_ALU/n233 [15]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u419  (\u_EXU_ALU/alu_or [16], i_decinfo[7], \u_EXU_ALU/n233 [16]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u420  (\u_EXU_ALU/alu_or [17], i_decinfo[7], \u_EXU_ALU/n233 [17]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u421  (\u_EXU_ALU/alu_or [18], i_decinfo[7], \u_EXU_ALU/n233 [18]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u422  (\u_EXU_ALU/alu_or [19], i_decinfo[7], \u_EXU_ALU/n233 [19]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u423  (\u_EXU_ALU/alu_or [20], i_decinfo[7], \u_EXU_ALU/n233 [20]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u424  (\u_EXU_ALU/alu_or [21], i_decinfo[7], \u_EXU_ALU/n233 [21]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u425  (\u_EXU_ALU/alu_or [22], i_decinfo[7], \u_EXU_ALU/n233 [22]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u426  (\u_EXU_ALU/alu_or [23], i_decinfo[7], \u_EXU_ALU/n233 [23]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u427  (\u_EXU_ALU/alu_or [24], i_decinfo[7], \u_EXU_ALU/n233 [24]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u428  (\u_EXU_ALU/alu_or [25], i_decinfo[7], \u_EXU_ALU/n233 [25]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u429  (\u_EXU_ALU/alu_or [26], i_decinfo[7], \u_EXU_ALU/n233 [26]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u430  (\u_EXU_ALU/alu_or [27], i_decinfo[7], \u_EXU_ALU/n233 [27]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u431  (\u_EXU_ALU/alu_or [28], i_decinfo[7], \u_EXU_ALU/n233 [28]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u432  (\u_EXU_ALU/alu_or [29], i_decinfo[7], \u_EXU_ALU/n233 [29]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u433  (\u_EXU_ALU/alu_or [30], i_decinfo[7], \u_EXU_ALU/n233 [30]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u434  (\u_EXU_ALU/alu_or [31], i_decinfo[7], \u_EXU_ALU/n233 [31]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u435  (\u_EXU_ALU/n233 [1], i_exu_op1[1], i_exu_op2[1]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u436  (\u_EXU_ALU/n233 [2], i_exu_op1[2], i_exu_op2[2]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u437  (\u_EXU_ALU/n233 [3], i_exu_op1[3], i_exu_op2[3]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u438  (\u_EXU_ALU/n233 [4], i_exu_op1[4], i_exu_op2[4]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u439  (\u_EXU_ALU/n233 [5], i_exu_op1[5], i_exu_op2[5]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u440  (\u_EXU_ALU/n233 [6], i_exu_op1[6], i_exu_op2[6]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u441  (\u_EXU_ALU/n233 [7], i_exu_op1[7], i_exu_op2[7]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u442  (\u_EXU_ALU/n233 [8], i_exu_op1[8], i_exu_op2[8]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u443  (\u_EXU_ALU/n233 [9], i_exu_op1[9], i_exu_op2[9]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u444  (\u_EXU_ALU/n233 [10], i_exu_op1[10], i_exu_op2[10]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u445  (\u_EXU_ALU/n233 [11], i_exu_op1[11], i_exu_op2[11]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u446  (\u_EXU_ALU/n233 [12], i_exu_op1[12], i_exu_op2[12]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u447  (\u_EXU_ALU/n233 [13], i_exu_op1[13], i_exu_op2[13]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u448  (\u_EXU_ALU/n233 [14], i_exu_op1[14], i_exu_op2[14]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u449  (\u_EXU_ALU/n233 [15], i_exu_op1[15], i_exu_op2[15]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u450  (\u_EXU_ALU/n233 [16], i_exu_op1[16], i_exu_op2[16]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u451  (\u_EXU_ALU/n233 [17], i_exu_op1[17], i_exu_op2[17]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u452  (\u_EXU_ALU/n233 [18], i_exu_op1[18], i_exu_op2[18]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u453  (\u_EXU_ALU/n233 [19], i_exu_op1[19], i_exu_op2[19]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u454  (\u_EXU_ALU/n233 [20], i_exu_op1[20], i_exu_op2[20]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u455  (\u_EXU_ALU/n233 [21], i_exu_op1[21], i_exu_op2[21]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u456  (\u_EXU_ALU/n233 [22], i_exu_op1[22], i_exu_op2[22]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u457  (\u_EXU_ALU/n233 [23], i_exu_op1[23], i_exu_op2[23]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u458  (\u_EXU_ALU/n233 [24], i_exu_op1[24], i_exu_op2[24]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u459  (\u_EXU_ALU/n233 [25], i_exu_op1[25], i_exu_op2[25]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u460  (\u_EXU_ALU/n233 [26], i_exu_op1[26], i_exu_op2[26]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u461  (\u_EXU_ALU/n233 [27], i_exu_op1[27], i_exu_op2[27]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u462  (\u_EXU_ALU/n233 [28], i_exu_op1[28], i_exu_op2[28]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u463  (\u_EXU_ALU/n233 [29], i_exu_op1[29], i_exu_op2[29]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u464  (\u_EXU_ALU/n233 [30], i_exu_op1[30], i_exu_op2[30]);  // ../RTL/core/exu_alu.v(53)
  or \u_EXU_ALU/u465  (\u_EXU_ALU/n233 [31], i_exu_op1[31], i_exu_op2[31]);  // ../RTL/core/exu_alu.v(53)
  and \u_EXU_ALU/u466  (\u_EXU_ALU/alu_and [1], i_decinfo[6], \u_EXU_ALU/n201 [1]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u467  (\u_EXU_ALU/alu_and [2], i_decinfo[6], \u_EXU_ALU/n201 [2]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u468  (\u_EXU_ALU/alu_and [3], i_decinfo[6], \u_EXU_ALU/n201 [3]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u469  (\u_EXU_ALU/alu_and [4], i_decinfo[6], \u_EXU_ALU/n201 [4]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u470  (\u_EXU_ALU/alu_and [5], i_decinfo[6], \u_EXU_ALU/n201 [5]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u471  (\u_EXU_ALU/alu_and [6], i_decinfo[6], \u_EXU_ALU/n201 [6]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u472  (\u_EXU_ALU/alu_and [7], i_decinfo[6], \u_EXU_ALU/n201 [7]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u473  (\u_EXU_ALU/alu_and [8], i_decinfo[6], \u_EXU_ALU/n201 [8]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u474  (\u_EXU_ALU/alu_and [9], i_decinfo[6], \u_EXU_ALU/n201 [9]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u475  (\u_EXU_ALU/alu_and [10], i_decinfo[6], \u_EXU_ALU/n201 [10]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u476  (\u_EXU_ALU/alu_and [11], i_decinfo[6], \u_EXU_ALU/n201 [11]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u477  (\u_EXU_ALU/alu_and [12], i_decinfo[6], \u_EXU_ALU/n201 [12]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u478  (\u_EXU_ALU/alu_and [13], i_decinfo[6], \u_EXU_ALU/n201 [13]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u479  (\u_EXU_ALU/alu_and [14], i_decinfo[6], \u_EXU_ALU/n201 [14]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u480  (\u_EXU_ALU/alu_and [15], i_decinfo[6], \u_EXU_ALU/n201 [15]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u481  (\u_EXU_ALU/alu_and [16], i_decinfo[6], \u_EXU_ALU/n201 [16]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u482  (\u_EXU_ALU/alu_and [17], i_decinfo[6], \u_EXU_ALU/n201 [17]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u483  (\u_EXU_ALU/alu_and [18], i_decinfo[6], \u_EXU_ALU/n201 [18]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u484  (\u_EXU_ALU/alu_and [19], i_decinfo[6], \u_EXU_ALU/n201 [19]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u485  (\u_EXU_ALU/alu_and [20], i_decinfo[6], \u_EXU_ALU/n201 [20]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u486  (\u_EXU_ALU/alu_and [21], i_decinfo[6], \u_EXU_ALU/n201 [21]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u487  (\u_EXU_ALU/alu_and [22], i_decinfo[6], \u_EXU_ALU/n201 [22]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u488  (\u_EXU_ALU/alu_and [23], i_decinfo[6], \u_EXU_ALU/n201 [23]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u489  (\u_EXU_ALU/alu_and [24], i_decinfo[6], \u_EXU_ALU/n201 [24]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u490  (\u_EXU_ALU/alu_and [25], i_decinfo[6], \u_EXU_ALU/n201 [25]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u491  (\u_EXU_ALU/alu_and [26], i_decinfo[6], \u_EXU_ALU/n201 [26]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u492  (\u_EXU_ALU/alu_and [27], i_decinfo[6], \u_EXU_ALU/n201 [27]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u493  (\u_EXU_ALU/alu_and [28], i_decinfo[6], \u_EXU_ALU/n201 [28]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u494  (\u_EXU_ALU/alu_and [29], i_decinfo[6], \u_EXU_ALU/n201 [29]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u495  (\u_EXU_ALU/alu_and [30], i_decinfo[6], \u_EXU_ALU/n201 [30]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u496  (\u_EXU_ALU/alu_and [31], i_decinfo[6], \u_EXU_ALU/n201 [31]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u497  (\u_EXU_ALU/n201 [1], i_exu_op1[1], i_exu_op2[1]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u498  (\u_EXU_ALU/n201 [2], i_exu_op1[2], i_exu_op2[2]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u499  (\u_EXU_ALU/n201 [3], i_exu_op1[3], i_exu_op2[3]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u5  (\u_EXU_ALU/alu_sub [0], i_decinfo[1], \u_EXU_ALU/n33 [0]);  // ../RTL/core/exu_alu.v(41)
  and \u_EXU_ALU/u500  (\u_EXU_ALU/n201 [4], i_exu_op1[4], i_exu_op2[4]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u501  (\u_EXU_ALU/n201 [5], i_exu_op1[5], i_exu_op2[5]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u502  (\u_EXU_ALU/n201 [6], i_exu_op1[6], i_exu_op2[6]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u503  (\u_EXU_ALU/n201 [7], i_exu_op1[7], i_exu_op2[7]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u504  (\u_EXU_ALU/n201 [8], i_exu_op1[8], i_exu_op2[8]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u505  (\u_EXU_ALU/n201 [9], i_exu_op1[9], i_exu_op2[9]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u506  (\u_EXU_ALU/n201 [10], i_exu_op1[10], i_exu_op2[10]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u507  (\u_EXU_ALU/n201 [11], i_exu_op1[11], i_exu_op2[11]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u508  (\u_EXU_ALU/n201 [12], i_exu_op1[12], i_exu_op2[12]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u509  (\u_EXU_ALU/n201 [13], i_exu_op1[13], i_exu_op2[13]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u510  (\u_EXU_ALU/n201 [14], i_exu_op1[14], i_exu_op2[14]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u511  (\u_EXU_ALU/n201 [15], i_exu_op1[15], i_exu_op2[15]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u512  (\u_EXU_ALU/n201 [16], i_exu_op1[16], i_exu_op2[16]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u513  (\u_EXU_ALU/n201 [17], i_exu_op1[17], i_exu_op2[17]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u514  (\u_EXU_ALU/n201 [18], i_exu_op1[18], i_exu_op2[18]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u515  (\u_EXU_ALU/n201 [19], i_exu_op1[19], i_exu_op2[19]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u516  (\u_EXU_ALU/n201 [20], i_exu_op1[20], i_exu_op2[20]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u517  (\u_EXU_ALU/n201 [21], i_exu_op1[21], i_exu_op2[21]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u518  (\u_EXU_ALU/n201 [22], i_exu_op1[22], i_exu_op2[22]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u519  (\u_EXU_ALU/n201 [23], i_exu_op1[23], i_exu_op2[23]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u520  (\u_EXU_ALU/n201 [24], i_exu_op1[24], i_exu_op2[24]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u521  (\u_EXU_ALU/n201 [25], i_exu_op1[25], i_exu_op2[25]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u522  (\u_EXU_ALU/n201 [26], i_exu_op1[26], i_exu_op2[26]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u523  (\u_EXU_ALU/n201 [27], i_exu_op1[27], i_exu_op2[27]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u524  (\u_EXU_ALU/n201 [28], i_exu_op1[28], i_exu_op2[28]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u525  (\u_EXU_ALU/n201 [29], i_exu_op1[29], i_exu_op2[29]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u526  (\u_EXU_ALU/n201 [30], i_exu_op1[30], i_exu_op2[30]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u527  (\u_EXU_ALU/n201 [31], i_exu_op1[31], i_exu_op2[31]);  // ../RTL/core/exu_alu.v(51)
  and \u_EXU_ALU/u528  (\u_EXU_ALU/alu_xor [1], i_decinfo[5], \u_EXU_ALU/n168 [1]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u529  (\u_EXU_ALU/alu_xor [2], i_decinfo[5], \u_EXU_ALU/n168 [2]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u530  (\u_EXU_ALU/alu_xor [3], i_decinfo[5], \u_EXU_ALU/n168 [3]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u531  (\u_EXU_ALU/alu_xor [4], i_decinfo[5], \u_EXU_ALU/n168 [4]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u532  (\u_EXU_ALU/alu_xor [5], i_decinfo[5], \u_EXU_ALU/n168 [5]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u533  (\u_EXU_ALU/alu_xor [6], i_decinfo[5], \u_EXU_ALU/n168 [6]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u534  (\u_EXU_ALU/alu_xor [7], i_decinfo[5], \u_EXU_ALU/n168 [7]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u535  (\u_EXU_ALU/alu_xor [8], i_decinfo[5], \u_EXU_ALU/n168 [8]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u536  (\u_EXU_ALU/alu_xor [9], i_decinfo[5], \u_EXU_ALU/n168 [9]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u537  (\u_EXU_ALU/alu_xor [10], i_decinfo[5], \u_EXU_ALU/n168 [10]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u538  (\u_EXU_ALU/alu_xor [11], i_decinfo[5], \u_EXU_ALU/n168 [11]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u539  (\u_EXU_ALU/alu_xor [12], i_decinfo[5], \u_EXU_ALU/n168 [12]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u540  (\u_EXU_ALU/alu_xor [13], i_decinfo[5], \u_EXU_ALU/n168 [13]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u541  (\u_EXU_ALU/alu_xor [14], i_decinfo[5], \u_EXU_ALU/n168 [14]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u542  (\u_EXU_ALU/alu_xor [15], i_decinfo[5], \u_EXU_ALU/n168 [15]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u543  (\u_EXU_ALU/alu_xor [16], i_decinfo[5], \u_EXU_ALU/n168 [16]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u544  (\u_EXU_ALU/alu_xor [17], i_decinfo[5], \u_EXU_ALU/n168 [17]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u545  (\u_EXU_ALU/alu_xor [18], i_decinfo[5], \u_EXU_ALU/n168 [18]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u546  (\u_EXU_ALU/alu_xor [19], i_decinfo[5], \u_EXU_ALU/n168 [19]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u547  (\u_EXU_ALU/alu_xor [20], i_decinfo[5], \u_EXU_ALU/n168 [20]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u548  (\u_EXU_ALU/alu_xor [21], i_decinfo[5], \u_EXU_ALU/n168 [21]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u549  (\u_EXU_ALU/alu_xor [22], i_decinfo[5], \u_EXU_ALU/n168 [22]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u550  (\u_EXU_ALU/alu_xor [23], i_decinfo[5], \u_EXU_ALU/n168 [23]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u551  (\u_EXU_ALU/alu_xor [24], i_decinfo[5], \u_EXU_ALU/n168 [24]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u552  (\u_EXU_ALU/alu_xor [25], i_decinfo[5], \u_EXU_ALU/n168 [25]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u553  (\u_EXU_ALU/alu_xor [26], i_decinfo[5], \u_EXU_ALU/n168 [26]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u554  (\u_EXU_ALU/alu_xor [27], i_decinfo[5], \u_EXU_ALU/n168 [27]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u555  (\u_EXU_ALU/alu_xor [28], i_decinfo[5], \u_EXU_ALU/n168 [28]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u556  (\u_EXU_ALU/alu_xor [29], i_decinfo[5], \u_EXU_ALU/n168 [29]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u557  (\u_EXU_ALU/alu_xor [30], i_decinfo[5], \u_EXU_ALU/n168 [30]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u558  (\u_EXU_ALU/alu_xor [31], i_decinfo[5], \u_EXU_ALU/n168 [31]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u559  (\u_EXU_ALU/n168 [1], i_exu_op1[1], i_exu_op2[1]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u560  (\u_EXU_ALU/n168 [2], i_exu_op1[2], i_exu_op2[2]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u561  (\u_EXU_ALU/n168 [3], i_exu_op1[3], i_exu_op2[3]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u562  (\u_EXU_ALU/n168 [4], i_exu_op1[4], i_exu_op2[4]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u563  (\u_EXU_ALU/n168 [5], i_exu_op1[5], i_exu_op2[5]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u564  (\u_EXU_ALU/n168 [6], i_exu_op1[6], i_exu_op2[6]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u565  (\u_EXU_ALU/n168 [7], i_exu_op1[7], i_exu_op2[7]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u566  (\u_EXU_ALU/n168 [8], i_exu_op1[8], i_exu_op2[8]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u567  (\u_EXU_ALU/n168 [9], i_exu_op1[9], i_exu_op2[9]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u568  (\u_EXU_ALU/n168 [10], i_exu_op1[10], i_exu_op2[10]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u569  (\u_EXU_ALU/n168 [11], i_exu_op1[11], i_exu_op2[11]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u570  (\u_EXU_ALU/n168 [12], i_exu_op1[12], i_exu_op2[12]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u571  (\u_EXU_ALU/n168 [13], i_exu_op1[13], i_exu_op2[13]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u572  (\u_EXU_ALU/n168 [14], i_exu_op1[14], i_exu_op2[14]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u573  (\u_EXU_ALU/n168 [15], i_exu_op1[15], i_exu_op2[15]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u574  (\u_EXU_ALU/n168 [16], i_exu_op1[16], i_exu_op2[16]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u575  (\u_EXU_ALU/n168 [17], i_exu_op1[17], i_exu_op2[17]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u576  (\u_EXU_ALU/n168 [18], i_exu_op1[18], i_exu_op2[18]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u577  (\u_EXU_ALU/n168 [19], i_exu_op1[19], i_exu_op2[19]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u578  (\u_EXU_ALU/n168 [20], i_exu_op1[20], i_exu_op2[20]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u579  (\u_EXU_ALU/n168 [21], i_exu_op1[21], i_exu_op2[21]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u580  (\u_EXU_ALU/n168 [22], i_exu_op1[22], i_exu_op2[22]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u581  (\u_EXU_ALU/n168 [23], i_exu_op1[23], i_exu_op2[23]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u582  (\u_EXU_ALU/n168 [24], i_exu_op1[24], i_exu_op2[24]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u583  (\u_EXU_ALU/n168 [25], i_exu_op1[25], i_exu_op2[25]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u584  (\u_EXU_ALU/n168 [26], i_exu_op1[26], i_exu_op2[26]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u585  (\u_EXU_ALU/n168 [27], i_exu_op1[27], i_exu_op2[27]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u586  (\u_EXU_ALU/n168 [28], i_exu_op1[28], i_exu_op2[28]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u587  (\u_EXU_ALU/n168 [29], i_exu_op1[29], i_exu_op2[29]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u588  (\u_EXU_ALU/n168 [30], i_exu_op1[30], i_exu_op2[30]);  // ../RTL/core/exu_alu.v(49)
  xor \u_EXU_ALU/u589  (\u_EXU_ALU/n168 [31], i_exu_op1[31], i_exu_op2[31]);  // ../RTL/core/exu_alu.v(49)
  and \u_EXU_ALU/u590  (\u_EXU_ALU/alu_sra [1], i_decinfo[4], \u_EXU_ALU/n135 [1]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u591  (\u_EXU_ALU/alu_sra [2], i_decinfo[4], \u_EXU_ALU/n135 [2]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u592  (\u_EXU_ALU/alu_sra [3], i_decinfo[4], \u_EXU_ALU/n135 [3]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u593  (\u_EXU_ALU/alu_sra [4], i_decinfo[4], \u_EXU_ALU/n135 [4]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u594  (\u_EXU_ALU/alu_sra [5], i_decinfo[4], \u_EXU_ALU/n135 [5]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u595  (\u_EXU_ALU/alu_sra [6], i_decinfo[4], \u_EXU_ALU/n135 [6]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u596  (\u_EXU_ALU/alu_sra [7], i_decinfo[4], \u_EXU_ALU/n135 [7]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u597  (\u_EXU_ALU/alu_sra [8], i_decinfo[4], \u_EXU_ALU/n135 [8]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u598  (\u_EXU_ALU/alu_sra [9], i_decinfo[4], \u_EXU_ALU/n135 [9]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u599  (\u_EXU_ALU/alu_sra [10], i_decinfo[4], \u_EXU_ALU/n135 [10]);  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u6  (
    .i0(i_exu_op1[31]),
    .i1(i_exu_op1[30]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n280 ));  // ../RTL/core/exu_alu.v(43)
  and \u_EXU_ALU/u600  (\u_EXU_ALU/alu_sra [11], i_decinfo[4], \u_EXU_ALU/n135 [11]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u601  (\u_EXU_ALU/alu_sra [12], i_decinfo[4], \u_EXU_ALU/n135 [12]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u602  (\u_EXU_ALU/alu_sra [13], i_decinfo[4], \u_EXU_ALU/n135 [13]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u603  (\u_EXU_ALU/alu_sra [14], i_decinfo[4], \u_EXU_ALU/n135 [14]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u604  (\u_EXU_ALU/alu_sra [15], i_decinfo[4], \u_EXU_ALU/n135 [15]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u605  (\u_EXU_ALU/alu_sra [16], i_decinfo[4], \u_EXU_ALU/n135 [16]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u606  (\u_EXU_ALU/alu_sra [17], i_decinfo[4], \u_EXU_ALU/n135 [17]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u607  (\u_EXU_ALU/alu_sra [18], i_decinfo[4], \u_EXU_ALU/n135 [18]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u608  (\u_EXU_ALU/alu_sra [19], i_decinfo[4], \u_EXU_ALU/n135 [19]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u609  (\u_EXU_ALU/alu_sra [20], i_decinfo[4], \u_EXU_ALU/n135 [20]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u610  (\u_EXU_ALU/alu_sra [21], i_decinfo[4], \u_EXU_ALU/n135 [21]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u611  (\u_EXU_ALU/alu_sra [22], i_decinfo[4], \u_EXU_ALU/n135 [22]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u612  (\u_EXU_ALU/alu_sra [23], i_decinfo[4], \u_EXU_ALU/n135 [23]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u613  (\u_EXU_ALU/alu_sra [24], i_decinfo[4], \u_EXU_ALU/n135 [24]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u614  (\u_EXU_ALU/alu_sra [25], i_decinfo[4], \u_EXU_ALU/n135 [25]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u615  (\u_EXU_ALU/alu_sra [26], i_decinfo[4], \u_EXU_ALU/n135 [26]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u616  (\u_EXU_ALU/alu_sra [27], i_decinfo[4], \u_EXU_ALU/n135 [27]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u617  (\u_EXU_ALU/alu_sra [28], i_decinfo[4], \u_EXU_ALU/n135 [28]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u618  (\u_EXU_ALU/alu_sra [29], i_decinfo[4], \u_EXU_ALU/n135 [29]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u619  (\u_EXU_ALU/alu_sra [30], i_decinfo[4], \u_EXU_ALU/n135 [30]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u620  (\u_EXU_ALU/alu_sra [31], i_decinfo[4], \u_EXU_ALU/n135 [31]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u621  (\u_EXU_ALU/n135 [1], \u_EXU_ALU/n133 [1], \u_EXU_ALU/n99 [1]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u622  (\u_EXU_ALU/n135 [2], \u_EXU_ALU/n133 [2], \u_EXU_ALU/n99 [2]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u623  (\u_EXU_ALU/n135 [3], \u_EXU_ALU/n133 [3], \u_EXU_ALU/n99 [3]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u624  (\u_EXU_ALU/n135 [4], \u_EXU_ALU/n133 [4], \u_EXU_ALU/n99 [4]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u625  (\u_EXU_ALU/n135 [5], \u_EXU_ALU/n133 [5], \u_EXU_ALU/n99 [5]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u626  (\u_EXU_ALU/n135 [6], \u_EXU_ALU/n133 [6], \u_EXU_ALU/n99 [6]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u627  (\u_EXU_ALU/n135 [7], \u_EXU_ALU/n133 [7], \u_EXU_ALU/n99 [7]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u628  (\u_EXU_ALU/n135 [8], \u_EXU_ALU/n133 [8], \u_EXU_ALU/n99 [8]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u629  (\u_EXU_ALU/n135 [9], \u_EXU_ALU/n133 [9], \u_EXU_ALU/n99 [9]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u630  (\u_EXU_ALU/n135 [10], \u_EXU_ALU/n133 [10], \u_EXU_ALU/n99 [10]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u631  (\u_EXU_ALU/n135 [11], \u_EXU_ALU/n133 [11], \u_EXU_ALU/n99 [11]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u632  (\u_EXU_ALU/n135 [12], \u_EXU_ALU/n133 [12], \u_EXU_ALU/n99 [12]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u633  (\u_EXU_ALU/n135 [13], \u_EXU_ALU/n133 [13], \u_EXU_ALU/n99 [13]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u634  (\u_EXU_ALU/n135 [14], \u_EXU_ALU/n133 [14], \u_EXU_ALU/n99 [14]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u635  (\u_EXU_ALU/n135 [15], \u_EXU_ALU/n133 [15], \u_EXU_ALU/n99 [15]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u636  (\u_EXU_ALU/n135 [16], \u_EXU_ALU/n133 [16], \u_EXU_ALU/n99 [16]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u637  (\u_EXU_ALU/n135 [17], \u_EXU_ALU/n133 [17], \u_EXU_ALU/n99 [17]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u638  (\u_EXU_ALU/n135 [18], \u_EXU_ALU/n133 [18], \u_EXU_ALU/n99 [18]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u639  (\u_EXU_ALU/n135 [19], \u_EXU_ALU/n133 [19], \u_EXU_ALU/n99 [19]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u640  (\u_EXU_ALU/n135 [20], \u_EXU_ALU/n133 [20], \u_EXU_ALU/n99 [20]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u641  (\u_EXU_ALU/n135 [21], \u_EXU_ALU/n133 [21], \u_EXU_ALU/n99 [21]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u642  (\u_EXU_ALU/n135 [22], \u_EXU_ALU/n133 [22], \u_EXU_ALU/n99 [22]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u643  (\u_EXU_ALU/n135 [23], \u_EXU_ALU/n133 [23], \u_EXU_ALU/n99 [23]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u644  (\u_EXU_ALU/n135 [24], \u_EXU_ALU/n133 [24], \u_EXU_ALU/n99 [24]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u645  (\u_EXU_ALU/n135 [25], \u_EXU_ALU/n133 [25], \u_EXU_ALU/n99 [25]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u646  (\u_EXU_ALU/n135 [26], \u_EXU_ALU/n133 [26], \u_EXU_ALU/n99 [26]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u647  (\u_EXU_ALU/n135 [27], \u_EXU_ALU/n133 [27], \u_EXU_ALU/n99 [27]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u648  (\u_EXU_ALU/n135 [28], \u_EXU_ALU/n133 [28], \u_EXU_ALU/n99 [28]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u649  (\u_EXU_ALU/n135 [29], \u_EXU_ALU/n133 [29], \u_EXU_ALU/n99 [29]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u650  (\u_EXU_ALU/n135 [30], \u_EXU_ALU/n133 [30], \u_EXU_ALU/n99 [30]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u651  (\u_EXU_ALU/n135 [31], \u_EXU_ALU/n133 [31], \u_EXU_ALU/n99 [31]);  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u652  (
    .i0(1'b0),
    .i1(i_exu_op1[31]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n134 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u653  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n134 ),
    .sel(\u_EXU_ALU/n132 [1]),
    .o(\u_EXU_ALU/n264 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u654  (
    .i0(i_exu_op1[31]),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [1]),
    .o(\u_EXU_ALU/n263 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u655  (
    .i0(\u_EXU_ALU/n134 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [1]),
    .o(\u_EXU_ALU/n262 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u656  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n264 ),
    .sel(\u_EXU_ALU/n132 [2]),
    .o(\u_EXU_ALU/n260 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u657  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n263 ),
    .sel(\u_EXU_ALU/n132 [2]),
    .o(\u_EXU_ALU/n259 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u658  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n262 ),
    .sel(\u_EXU_ALU/n132 [2]),
    .o(\u_EXU_ALU/n258 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u659  (
    .i0(i_exu_op1[31]),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [2]),
    .o(\u_EXU_ALU/n257 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u660  (
    .i0(\u_EXU_ALU/n264 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [2]),
    .o(\u_EXU_ALU/n256 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u661  (
    .i0(\u_EXU_ALU/n263 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [2]),
    .o(\u_EXU_ALU/n255 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u662  (
    .i0(\u_EXU_ALU/n262 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [2]),
    .o(\u_EXU_ALU/n254 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u663  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n260 ),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n252 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u664  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n259 ),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n251 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u665  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n258 ),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n250 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u666  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n257 ),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n249 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u667  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n256 ),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n248 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u668  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n255 ),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n247 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u669  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n254 ),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n246 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u670  (
    .i0(i_exu_op1[31]),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n245 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u671  (
    .i0(\u_EXU_ALU/n260 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n244 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u672  (
    .i0(\u_EXU_ALU/n259 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n243 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u673  (
    .i0(\u_EXU_ALU/n258 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n242 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u674  (
    .i0(\u_EXU_ALU/n257 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n241 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u675  (
    .i0(\u_EXU_ALU/n256 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n240 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u676  (
    .i0(\u_EXU_ALU/n255 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n239 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u677  (
    .i0(\u_EXU_ALU/n254 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n132 [3]),
    .o(\u_EXU_ALU/n238 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u678  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n252 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n237 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u679  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n251 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n236 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u680  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n250 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n235 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u681  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n249 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n234 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u682  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n248 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n232 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u683  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n247 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n231 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u684  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n246 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n230 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u685  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n245 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n229 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u686  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n244 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n228 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u687  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n243 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n227 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u688  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n242 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n226 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u689  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n241 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n225 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u690  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n240 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n224 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u691  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n239 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n223 ));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u692  (
    .i0(i_exu_op1[31]),
    .i1(\u_EXU_ALU/n238 ),
    .sel(\i_exu_op2[4]_neg ),
    .o(\u_EXU_ALU/n222 ));  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u7  (\u_EXU_ALU/alu_sll [0], i_decinfo[2], \u_EXU_ALU/n66 [0]);  // ../RTL/core/exu_alu.v(43)
  or \u_EXU_ALU/u709  (\u_EXU_ALU/n205 , \u_EXU_ALU/n132 [6], \u_EXU_ALU/n132 [7]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u710  (\u_EXU_ALU/n204 , \u_EXU_ALU/n132 [5], \u_EXU_ALU/n205 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u711  (\u_EXU_ALU/n203 , \u_EXU_ALU/n132 [9], \u_EXU_ALU/n132 [10]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u712  (\u_EXU_ALU/n202 , \u_EXU_ALU/n132 [8], \u_EXU_ALU/n203 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u713  (\u_EXU_ALU/n200 , \u_EXU_ALU/n204 , \u_EXU_ALU/n202 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u714  (\u_EXU_ALU/n199 , \u_EXU_ALU/n132 [12], \u_EXU_ALU/n132 [13]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u715  (\u_EXU_ALU/n198 , \u_EXU_ALU/n132 [11], \u_EXU_ALU/n199 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u716  (\u_EXU_ALU/n197 , \u_EXU_ALU/n132 [14], \u_EXU_ALU/n132 [15]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u717  (\u_EXU_ALU/n196 , \u_EXU_ALU/n132 [16], \u_EXU_ALU/n132 [17]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u718  (\u_EXU_ALU/n195 , \u_EXU_ALU/n197 , \u_EXU_ALU/n196 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u719  (\u_EXU_ALU/n194 , \u_EXU_ALU/n198 , \u_EXU_ALU/n195 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u720  (\u_EXU_ALU/n193 , \u_EXU_ALU/n200 , \u_EXU_ALU/n194 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u721  (\u_EXU_ALU/n192 , \u_EXU_ALU/n132 [19], \u_EXU_ALU/n132 [20]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u722  (\u_EXU_ALU/n191 , \u_EXU_ALU/n132 [18], \u_EXU_ALU/n192 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u723  (\u_EXU_ALU/n190 , \u_EXU_ALU/n132 [21], \u_EXU_ALU/n132 [22]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u724  (\u_EXU_ALU/n189 , \u_EXU_ALU/n132 [23], \u_EXU_ALU/n132 [24]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u725  (\u_EXU_ALU/n188 , \u_EXU_ALU/n190 , \u_EXU_ALU/n189 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u726  (\u_EXU_ALU/n187 , \u_EXU_ALU/n191 , \u_EXU_ALU/n188 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u727  (\u_EXU_ALU/n186 , \u_EXU_ALU/n132 [26], \u_EXU_ALU/n132 [27]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u728  (\u_EXU_ALU/n185 , \u_EXU_ALU/n132 [25], \u_EXU_ALU/n186 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u729  (\u_EXU_ALU/n184 , \u_EXU_ALU/n132 [28], \u_EXU_ALU/n132 [29]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u730  (\u_EXU_ALU/n183 , \u_EXU_ALU/n132 [30], \u_EXU_ALU/n132 [31]);  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u731  (\u_EXU_ALU/n182 , \u_EXU_ALU/n184 , \u_EXU_ALU/n183 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u732  (\u_EXU_ALU/n181 , \u_EXU_ALU/n185 , \u_EXU_ALU/n182 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u733  (\u_EXU_ALU/n180 , \u_EXU_ALU/n187 , \u_EXU_ALU/n181 );  // ../RTL/core/exu_alu.v(47)
  or \u_EXU_ALU/u734  (\u_EXU_ALU/n179 , \u_EXU_ALU/n193 , \u_EXU_ALU/n180 );  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u735  (
    .i0(\u_EXU_ALU/n237 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [31]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u736  (
    .i0(\u_EXU_ALU/n236 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [30]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u737  (
    .i0(\u_EXU_ALU/n235 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [29]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u738  (
    .i0(\u_EXU_ALU/n234 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [28]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u739  (
    .i0(\u_EXU_ALU/n232 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [27]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u740  (
    .i0(\u_EXU_ALU/n231 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [26]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u741  (
    .i0(\u_EXU_ALU/n230 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [25]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u742  (
    .i0(\u_EXU_ALU/n229 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [24]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u743  (
    .i0(\u_EXU_ALU/n228 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [23]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u744  (
    .i0(\u_EXU_ALU/n227 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [22]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u745  (
    .i0(\u_EXU_ALU/n226 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [21]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u746  (
    .i0(\u_EXU_ALU/n225 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [20]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u747  (
    .i0(\u_EXU_ALU/n224 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [19]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u748  (
    .i0(\u_EXU_ALU/n223 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [18]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u749  (
    .i0(\u_EXU_ALU/n222 ),
    .i1(1'b0),
    .sel(\u_EXU_ALU/n179 ),
    .o(\u_EXU_ALU/n133 [17]));  // ../RTL/core/exu_alu.v(47)
  AL_MUX \u_EXU_ALU/u750  (
    .i0(1'b0),
    .i1(i_exu_op1[31]),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [16]));
  and \u_EXU_ALU/u750_sel_is_0  (\u_EXU_ALU/u750_sel_is_0_o , \u_EXU_ALU/n179_neg , i_exu_op2[4]);
  AL_MUX \u_EXU_ALU/u751  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n252 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [15]));
  AL_MUX \u_EXU_ALU/u752  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n251 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [14]));
  AL_MUX \u_EXU_ALU/u753  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n250 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [13]));
  AL_MUX \u_EXU_ALU/u754  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n249 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [12]));
  AL_MUX \u_EXU_ALU/u755  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n248 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [11]));
  AL_MUX \u_EXU_ALU/u756  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n247 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [10]));
  AL_MUX \u_EXU_ALU/u757  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n246 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [9]));
  AL_MUX \u_EXU_ALU/u758  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n245 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [8]));
  AL_MUX \u_EXU_ALU/u759  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n244 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [7]));
  AL_MUX \u_EXU_ALU/u760  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n243 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [6]));
  AL_MUX \u_EXU_ALU/u761  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n242 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [5]));
  AL_MUX \u_EXU_ALU/u762  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n241 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [4]));
  AL_MUX \u_EXU_ALU/u763  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n240 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [3]));
  AL_MUX \u_EXU_ALU/u764  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n239 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [2]));
  AL_MUX \u_EXU_ALU/u765  (
    .i0(1'b0),
    .i1(\u_EXU_ALU/n238 ),
    .sel(\u_EXU_ALU/u750_sel_is_0_o ),
    .o(\u_EXU_ALU/n133 [1]));
  not \u_EXU_ALU/u766  (\u_EXU_ALU/n132 [1], i_exu_op2[1]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u767  (\u_EXU_ALU/n132 [2], i_exu_op2[2]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u768  (\u_EXU_ALU/n132 [3], i_exu_op2[3]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u770  (\u_EXU_ALU/n132 [5], i_exu_op2[5]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u771  (\u_EXU_ALU/n132 [6], i_exu_op2[6]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u772  (\u_EXU_ALU/n132 [7], i_exu_op2[7]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u773  (\u_EXU_ALU/n132 [8], i_exu_op2[8]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u774  (\u_EXU_ALU/n132 [9], i_exu_op2[9]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u775  (\u_EXU_ALU/n132 [10], i_exu_op2[10]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u776  (\u_EXU_ALU/n132 [11], i_exu_op2[11]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u777  (\u_EXU_ALU/n132 [12], i_exu_op2[12]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u778  (\u_EXU_ALU/n132 [13], i_exu_op2[13]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u779  (\u_EXU_ALU/n132 [14], i_exu_op2[14]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u780  (\u_EXU_ALU/n132 [15], i_exu_op2[15]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u781  (\u_EXU_ALU/n132 [16], i_exu_op2[16]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u782  (\u_EXU_ALU/n132 [17], i_exu_op2[17]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u783  (\u_EXU_ALU/n132 [18], i_exu_op2[18]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u784  (\u_EXU_ALU/n132 [19], i_exu_op2[19]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u785  (\u_EXU_ALU/n132 [20], i_exu_op2[20]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u786  (\u_EXU_ALU/n132 [21], i_exu_op2[21]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u787  (\u_EXU_ALU/n132 [22], i_exu_op2[22]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u788  (\u_EXU_ALU/n132 [23], i_exu_op2[23]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u789  (\u_EXU_ALU/n132 [24], i_exu_op2[24]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u790  (\u_EXU_ALU/n132 [25], i_exu_op2[25]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u791  (\u_EXU_ALU/n132 [26], i_exu_op2[26]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u792  (\u_EXU_ALU/n132 [27], i_exu_op2[27]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u793  (\u_EXU_ALU/n132 [28], i_exu_op2[28]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u794  (\u_EXU_ALU/n132 [29], i_exu_op2[29]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u795  (\u_EXU_ALU/n132 [30], i_exu_op2[30]);  // ../RTL/core/exu_alu.v(47)
  not \u_EXU_ALU/u796  (\u_EXU_ALU/n132 [31], i_exu_op2[31]);  // ../RTL/core/exu_alu.v(47)
  and \u_EXU_ALU/u797  (\u_EXU_ALU/alu_srl [1], i_decinfo[3], \u_EXU_ALU/n99 [1]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u798  (\u_EXU_ALU/alu_srl [2], i_decinfo[3], \u_EXU_ALU/n99 [2]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u799  (\u_EXU_ALU/alu_srl [3], i_decinfo[3], \u_EXU_ALU/n99 [3]);  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u8  (
    .i0(i_exu_op1[0]),
    .i1(i_exu_op1[1]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n178 ));  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u800  (\u_EXU_ALU/alu_srl [4], i_decinfo[3], \u_EXU_ALU/n99 [4]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u801  (\u_EXU_ALU/alu_srl [5], i_decinfo[3], \u_EXU_ALU/n99 [5]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u802  (\u_EXU_ALU/alu_srl [6], i_decinfo[3], \u_EXU_ALU/n99 [6]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u803  (\u_EXU_ALU/alu_srl [7], i_decinfo[3], \u_EXU_ALU/n99 [7]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u804  (\u_EXU_ALU/alu_srl [8], i_decinfo[3], \u_EXU_ALU/n99 [8]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u805  (\u_EXU_ALU/alu_srl [9], i_decinfo[3], \u_EXU_ALU/n99 [9]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u806  (\u_EXU_ALU/alu_srl [10], i_decinfo[3], \u_EXU_ALU/n99 [10]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u807  (\u_EXU_ALU/alu_srl [11], i_decinfo[3], \u_EXU_ALU/n99 [11]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u808  (\u_EXU_ALU/alu_srl [12], i_decinfo[3], \u_EXU_ALU/n99 [12]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u809  (\u_EXU_ALU/alu_srl [13], i_decinfo[3], \u_EXU_ALU/n99 [13]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u810  (\u_EXU_ALU/alu_srl [14], i_decinfo[3], \u_EXU_ALU/n99 [14]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u811  (\u_EXU_ALU/alu_srl [15], i_decinfo[3], \u_EXU_ALU/n99 [15]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u812  (\u_EXU_ALU/alu_srl [16], i_decinfo[3], \u_EXU_ALU/n99 [16]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u813  (\u_EXU_ALU/alu_srl [17], i_decinfo[3], \u_EXU_ALU/n99 [17]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u814  (\u_EXU_ALU/alu_srl [18], i_decinfo[3], \u_EXU_ALU/n99 [18]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u815  (\u_EXU_ALU/alu_srl [19], i_decinfo[3], \u_EXU_ALU/n99 [19]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u816  (\u_EXU_ALU/alu_srl [20], i_decinfo[3], \u_EXU_ALU/n99 [20]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u817  (\u_EXU_ALU/alu_srl [21], i_decinfo[3], \u_EXU_ALU/n99 [21]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u818  (\u_EXU_ALU/alu_srl [22], i_decinfo[3], \u_EXU_ALU/n99 [22]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u819  (\u_EXU_ALU/alu_srl [23], i_decinfo[3], \u_EXU_ALU/n99 [23]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u820  (\u_EXU_ALU/alu_srl [24], i_decinfo[3], \u_EXU_ALU/n99 [24]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u821  (\u_EXU_ALU/alu_srl [25], i_decinfo[3], \u_EXU_ALU/n99 [25]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u822  (\u_EXU_ALU/alu_srl [26], i_decinfo[3], \u_EXU_ALU/n99 [26]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u823  (\u_EXU_ALU/alu_srl [27], i_decinfo[3], \u_EXU_ALU/n99 [27]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u824  (\u_EXU_ALU/alu_srl [28], i_decinfo[3], \u_EXU_ALU/n99 [28]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u825  (\u_EXU_ALU/alu_srl [29], i_decinfo[3], \u_EXU_ALU/n99 [29]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u826  (\u_EXU_ALU/alu_srl [30], i_decinfo[3], \u_EXU_ALU/n99 [30]);  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u827  (\u_EXU_ALU/alu_srl [31], i_decinfo[3], \u_EXU_ALU/n99 [31]);  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u828  (
    .i0(i_exu_op1[1]),
    .i1(i_exu_op1[2]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n177 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u829  (
    .i0(i_exu_op1[2]),
    .i1(i_exu_op1[3]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n176 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u830  (
    .i0(i_exu_op1[3]),
    .i1(i_exu_op1[4]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n175 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u831  (
    .i0(i_exu_op1[4]),
    .i1(i_exu_op1[5]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n174 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u832  (
    .i0(i_exu_op1[5]),
    .i1(i_exu_op1[6]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n173 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u833  (
    .i0(i_exu_op1[6]),
    .i1(i_exu_op1[7]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n172 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u834  (
    .i0(i_exu_op1[7]),
    .i1(i_exu_op1[8]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n171 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u835  (
    .i0(i_exu_op1[8]),
    .i1(i_exu_op1[9]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n170 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u836  (
    .i0(i_exu_op1[9]),
    .i1(i_exu_op1[10]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n169 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u837  (
    .i0(i_exu_op1[10]),
    .i1(i_exu_op1[11]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n167 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u838  (
    .i0(i_exu_op1[11]),
    .i1(i_exu_op1[12]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n166 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u839  (
    .i0(i_exu_op1[12]),
    .i1(i_exu_op1[13]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n165 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u840  (
    .i0(i_exu_op1[13]),
    .i1(i_exu_op1[14]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n164 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u841  (
    .i0(i_exu_op1[14]),
    .i1(i_exu_op1[15]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n163 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u842  (
    .i0(i_exu_op1[15]),
    .i1(i_exu_op1[16]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n162 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u843  (
    .i0(i_exu_op1[16]),
    .i1(i_exu_op1[17]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n161 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u844  (
    .i0(i_exu_op1[17]),
    .i1(i_exu_op1[18]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n160 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u845  (
    .i0(i_exu_op1[18]),
    .i1(i_exu_op1[19]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n159 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u846  (
    .i0(i_exu_op1[19]),
    .i1(i_exu_op1[20]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n158 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u847  (
    .i0(i_exu_op1[20]),
    .i1(i_exu_op1[21]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n157 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u848  (
    .i0(i_exu_op1[21]),
    .i1(i_exu_op1[22]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n156 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u849  (
    .i0(i_exu_op1[22]),
    .i1(i_exu_op1[23]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n155 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u850  (
    .i0(i_exu_op1[23]),
    .i1(i_exu_op1[24]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n154 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u851  (
    .i0(i_exu_op1[24]),
    .i1(i_exu_op1[25]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n153 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u852  (
    .i0(i_exu_op1[25]),
    .i1(i_exu_op1[26]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n152 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u853  (
    .i0(i_exu_op1[26]),
    .i1(i_exu_op1[27]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n151 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u854  (
    .i0(i_exu_op1[27]),
    .i1(i_exu_op1[28]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n150 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u855  (
    .i0(i_exu_op1[28]),
    .i1(i_exu_op1[29]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n149 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u856  (
    .i0(i_exu_op1[29]),
    .i1(i_exu_op1[30]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n148 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u857  (
    .i0(i_exu_op1[30]),
    .i1(i_exu_op1[31]),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n147 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u858  (
    .i0(i_exu_op1[31]),
    .i1(1'b0),
    .sel(i_exu_op2[0]),
    .o(\u_EXU_ALU/n146 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u859  (
    .i0(\u_EXU_ALU/n178 ),
    .i1(\u_EXU_ALU/n176 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n145 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u860  (
    .i0(\u_EXU_ALU/n177 ),
    .i1(\u_EXU_ALU/n175 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n144 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u861  (
    .i0(\u_EXU_ALU/n176 ),
    .i1(\u_EXU_ALU/n174 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n143 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u862  (
    .i0(\u_EXU_ALU/n175 ),
    .i1(\u_EXU_ALU/n173 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n142 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u863  (
    .i0(\u_EXU_ALU/n174 ),
    .i1(\u_EXU_ALU/n172 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n141 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u864  (
    .i0(\u_EXU_ALU/n173 ),
    .i1(\u_EXU_ALU/n171 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n140 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u865  (
    .i0(\u_EXU_ALU/n172 ),
    .i1(\u_EXU_ALU/n170 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n139 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u866  (
    .i0(\u_EXU_ALU/n171 ),
    .i1(\u_EXU_ALU/n169 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n138 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u867  (
    .i0(\u_EXU_ALU/n170 ),
    .i1(\u_EXU_ALU/n167 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n137 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u868  (
    .i0(\u_EXU_ALU/n169 ),
    .i1(\u_EXU_ALU/n166 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n136 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u869  (
    .i0(\u_EXU_ALU/n167 ),
    .i1(\u_EXU_ALU/n165 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n131 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u870  (
    .i0(\u_EXU_ALU/n166 ),
    .i1(\u_EXU_ALU/n164 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n130 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u871  (
    .i0(\u_EXU_ALU/n165 ),
    .i1(\u_EXU_ALU/n163 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n129 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u872  (
    .i0(\u_EXU_ALU/n164 ),
    .i1(\u_EXU_ALU/n162 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n128 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u873  (
    .i0(\u_EXU_ALU/n163 ),
    .i1(\u_EXU_ALU/n161 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n127 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u874  (
    .i0(\u_EXU_ALU/n162 ),
    .i1(\u_EXU_ALU/n160 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n126 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u875  (
    .i0(\u_EXU_ALU/n161 ),
    .i1(\u_EXU_ALU/n159 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n125 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u876  (
    .i0(\u_EXU_ALU/n160 ),
    .i1(\u_EXU_ALU/n158 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n124 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u877  (
    .i0(\u_EXU_ALU/n159 ),
    .i1(\u_EXU_ALU/n157 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n123 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u878  (
    .i0(\u_EXU_ALU/n158 ),
    .i1(\u_EXU_ALU/n156 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n122 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u879  (
    .i0(\u_EXU_ALU/n157 ),
    .i1(\u_EXU_ALU/n155 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n121 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u880  (
    .i0(\u_EXU_ALU/n156 ),
    .i1(\u_EXU_ALU/n154 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n120 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u881  (
    .i0(\u_EXU_ALU/n155 ),
    .i1(\u_EXU_ALU/n153 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n119 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u882  (
    .i0(\u_EXU_ALU/n154 ),
    .i1(\u_EXU_ALU/n152 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n118 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u883  (
    .i0(\u_EXU_ALU/n153 ),
    .i1(\u_EXU_ALU/n151 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n117 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u884  (
    .i0(\u_EXU_ALU/n152 ),
    .i1(\u_EXU_ALU/n150 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n116 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u885  (
    .i0(\u_EXU_ALU/n151 ),
    .i1(\u_EXU_ALU/n149 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n115 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u886  (
    .i0(\u_EXU_ALU/n150 ),
    .i1(\u_EXU_ALU/n148 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n114 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u887  (
    .i0(\u_EXU_ALU/n149 ),
    .i1(\u_EXU_ALU/n147 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n113 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u888  (
    .i0(\u_EXU_ALU/n148 ),
    .i1(\u_EXU_ALU/n146 ),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n112 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u889  (
    .i0(\u_EXU_ALU/n147 ),
    .i1(1'b0),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n111 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u890  (
    .i0(\u_EXU_ALU/n146 ),
    .i1(1'b0),
    .sel(i_exu_op2[1]),
    .o(\u_EXU_ALU/n110 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u891  (
    .i0(\u_EXU_ALU/n145 ),
    .i1(\u_EXU_ALU/n141 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n109 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u892  (
    .i0(\u_EXU_ALU/n144 ),
    .i1(\u_EXU_ALU/n140 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n108 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u893  (
    .i0(\u_EXU_ALU/n143 ),
    .i1(\u_EXU_ALU/n139 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n107 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u894  (
    .i0(\u_EXU_ALU/n142 ),
    .i1(\u_EXU_ALU/n138 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n106 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u895  (
    .i0(\u_EXU_ALU/n141 ),
    .i1(\u_EXU_ALU/n137 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n105 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u896  (
    .i0(\u_EXU_ALU/n140 ),
    .i1(\u_EXU_ALU/n136 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n104 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u897  (
    .i0(\u_EXU_ALU/n139 ),
    .i1(\u_EXU_ALU/n131 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n103 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u898  (
    .i0(\u_EXU_ALU/n138 ),
    .i1(\u_EXU_ALU/n130 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n102 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u899  (
    .i0(\u_EXU_ALU/n137 ),
    .i1(\u_EXU_ALU/n129 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n101 ));  // ../RTL/core/exu_alu.v(45)
  and \u_EXU_ALU/u9  (\u_EXU_ALU/alu_srl [0], i_decinfo[3], \u_EXU_ALU/n99 [0]);  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u90  (\u_EXU_ALU/n309 [1], \u_EXU_ALU/n308 [1], \u_EXU_ALU/alu_or [1]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u900  (
    .i0(\u_EXU_ALU/n136 ),
    .i1(\u_EXU_ALU/n128 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n100 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u901  (
    .i0(\u_EXU_ALU/n131 ),
    .i1(\u_EXU_ALU/n127 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n98 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u902  (
    .i0(\u_EXU_ALU/n130 ),
    .i1(\u_EXU_ALU/n126 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n97 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u903  (
    .i0(\u_EXU_ALU/n129 ),
    .i1(\u_EXU_ALU/n125 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n96 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u904  (
    .i0(\u_EXU_ALU/n128 ),
    .i1(\u_EXU_ALU/n124 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n95 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u905  (
    .i0(\u_EXU_ALU/n127 ),
    .i1(\u_EXU_ALU/n123 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n94 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u906  (
    .i0(\u_EXU_ALU/n126 ),
    .i1(\u_EXU_ALU/n122 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n93 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u907  (
    .i0(\u_EXU_ALU/n125 ),
    .i1(\u_EXU_ALU/n121 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n92 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u908  (
    .i0(\u_EXU_ALU/n124 ),
    .i1(\u_EXU_ALU/n120 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n91 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u909  (
    .i0(\u_EXU_ALU/n123 ),
    .i1(\u_EXU_ALU/n119 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n90 ));  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u91  (\u_EXU_ALU/n309 [2], \u_EXU_ALU/n308 [2], \u_EXU_ALU/alu_or [2]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u910  (
    .i0(\u_EXU_ALU/n122 ),
    .i1(\u_EXU_ALU/n118 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n89 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u911  (
    .i0(\u_EXU_ALU/n121 ),
    .i1(\u_EXU_ALU/n117 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n88 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u912  (
    .i0(\u_EXU_ALU/n120 ),
    .i1(\u_EXU_ALU/n116 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n87 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u913  (
    .i0(\u_EXU_ALU/n119 ),
    .i1(\u_EXU_ALU/n115 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n86 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u914  (
    .i0(\u_EXU_ALU/n118 ),
    .i1(\u_EXU_ALU/n114 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n85 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u915  (
    .i0(\u_EXU_ALU/n117 ),
    .i1(\u_EXU_ALU/n113 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n84 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u916  (
    .i0(\u_EXU_ALU/n116 ),
    .i1(\u_EXU_ALU/n112 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n83 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u917  (
    .i0(\u_EXU_ALU/n115 ),
    .i1(\u_EXU_ALU/n111 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n82 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u918  (
    .i0(\u_EXU_ALU/n114 ),
    .i1(\u_EXU_ALU/n110 ),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n81 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u919  (
    .i0(\u_EXU_ALU/n113 ),
    .i1(1'b0),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n80 ));  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u92  (\u_EXU_ALU/n309 [3], \u_EXU_ALU/n308 [3], \u_EXU_ALU/alu_or [3]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u920  (
    .i0(\u_EXU_ALU/n112 ),
    .i1(1'b0),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n79 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u921  (
    .i0(\u_EXU_ALU/n111 ),
    .i1(1'b0),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n78 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u922  (
    .i0(\u_EXU_ALU/n110 ),
    .i1(1'b0),
    .sel(i_exu_op2[2]),
    .o(\u_EXU_ALU/n77 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u923  (
    .i0(\u_EXU_ALU/n109 ),
    .i1(\u_EXU_ALU/n101 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n76 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u924  (
    .i0(\u_EXU_ALU/n108 ),
    .i1(\u_EXU_ALU/n100 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n75 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u925  (
    .i0(\u_EXU_ALU/n107 ),
    .i1(\u_EXU_ALU/n98 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n74 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u926  (
    .i0(\u_EXU_ALU/n106 ),
    .i1(\u_EXU_ALU/n97 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n73 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u927  (
    .i0(\u_EXU_ALU/n105 ),
    .i1(\u_EXU_ALU/n96 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n72 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u928  (
    .i0(\u_EXU_ALU/n104 ),
    .i1(\u_EXU_ALU/n95 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n71 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u929  (
    .i0(\u_EXU_ALU/n103 ),
    .i1(\u_EXU_ALU/n94 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n70 ));  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u93  (\u_EXU_ALU/n309 [4], \u_EXU_ALU/n308 [4], \u_EXU_ALU/alu_or [4]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u930  (
    .i0(\u_EXU_ALU/n102 ),
    .i1(\u_EXU_ALU/n93 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n69 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u931  (
    .i0(\u_EXU_ALU/n101 ),
    .i1(\u_EXU_ALU/n92 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n68 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u932  (
    .i0(\u_EXU_ALU/n100 ),
    .i1(\u_EXU_ALU/n91 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n67 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u933  (
    .i0(\u_EXU_ALU/n98 ),
    .i1(\u_EXU_ALU/n90 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n65 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u934  (
    .i0(\u_EXU_ALU/n97 ),
    .i1(\u_EXU_ALU/n89 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n64 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u935  (
    .i0(\u_EXU_ALU/n96 ),
    .i1(\u_EXU_ALU/n88 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n63 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u936  (
    .i0(\u_EXU_ALU/n95 ),
    .i1(\u_EXU_ALU/n87 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n62 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u937  (
    .i0(\u_EXU_ALU/n94 ),
    .i1(\u_EXU_ALU/n86 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n61 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u938  (
    .i0(\u_EXU_ALU/n93 ),
    .i1(\u_EXU_ALU/n85 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n60 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u939  (
    .i0(\u_EXU_ALU/n92 ),
    .i1(\u_EXU_ALU/n84 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n59 ));  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u94  (\u_EXU_ALU/n309 [5], \u_EXU_ALU/n308 [5], \u_EXU_ALU/alu_or [5]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u940  (
    .i0(\u_EXU_ALU/n91 ),
    .i1(\u_EXU_ALU/n83 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n58 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u941  (
    .i0(\u_EXU_ALU/n90 ),
    .i1(\u_EXU_ALU/n82 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n57 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u942  (
    .i0(\u_EXU_ALU/n89 ),
    .i1(\u_EXU_ALU/n81 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n56 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u943  (
    .i0(\u_EXU_ALU/n88 ),
    .i1(\u_EXU_ALU/n80 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n55 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u944  (
    .i0(\u_EXU_ALU/n87 ),
    .i1(\u_EXU_ALU/n79 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n54 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u945  (
    .i0(\u_EXU_ALU/n86 ),
    .i1(\u_EXU_ALU/n78 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n53 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u946  (
    .i0(\u_EXU_ALU/n85 ),
    .i1(\u_EXU_ALU/n77 ),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n52 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u947  (
    .i0(\u_EXU_ALU/n84 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n51 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u948  (
    .i0(\u_EXU_ALU/n83 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n50 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u949  (
    .i0(\u_EXU_ALU/n82 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n49 ));  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u95  (\u_EXU_ALU/n309 [6], \u_EXU_ALU/n308 [6], \u_EXU_ALU/alu_or [6]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u950  (
    .i0(\u_EXU_ALU/n81 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n48 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u951  (
    .i0(\u_EXU_ALU/n80 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n47 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u952  (
    .i0(\u_EXU_ALU/n79 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n46 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u953  (
    .i0(\u_EXU_ALU/n78 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n45 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u954  (
    .i0(\u_EXU_ALU/n77 ),
    .i1(1'b0),
    .sel(i_exu_op2[3]),
    .o(\u_EXU_ALU/n44 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u955  (
    .i0(\u_EXU_ALU/n76 ),
    .i1(\u_EXU_ALU/n59 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n43 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u956  (
    .i0(\u_EXU_ALU/n75 ),
    .i1(\u_EXU_ALU/n58 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n42 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u957  (
    .i0(\u_EXU_ALU/n74 ),
    .i1(\u_EXU_ALU/n57 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n41 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u958  (
    .i0(\u_EXU_ALU/n73 ),
    .i1(\u_EXU_ALU/n56 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n40 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u959  (
    .i0(\u_EXU_ALU/n72 ),
    .i1(\u_EXU_ALU/n55 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n39 ));  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u96  (\u_EXU_ALU/n309 [7], \u_EXU_ALU/n308 [7], \u_EXU_ALU/alu_or [7]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u960  (
    .i0(\u_EXU_ALU/n71 ),
    .i1(\u_EXU_ALU/n54 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n38 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u961  (
    .i0(\u_EXU_ALU/n70 ),
    .i1(\u_EXU_ALU/n53 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n37 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u962  (
    .i0(\u_EXU_ALU/n69 ),
    .i1(\u_EXU_ALU/n52 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n36 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u963  (
    .i0(\u_EXU_ALU/n68 ),
    .i1(\u_EXU_ALU/n51 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n35 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u964  (
    .i0(\u_EXU_ALU/n67 ),
    .i1(\u_EXU_ALU/n50 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n34 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u965  (
    .i0(\u_EXU_ALU/n65 ),
    .i1(\u_EXU_ALU/n49 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n32 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u966  (
    .i0(\u_EXU_ALU/n64 ),
    .i1(\u_EXU_ALU/n48 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n31 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u967  (
    .i0(\u_EXU_ALU/n63 ),
    .i1(\u_EXU_ALU/n47 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n30 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u968  (
    .i0(\u_EXU_ALU/n62 ),
    .i1(\u_EXU_ALU/n46 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n29 ));  // ../RTL/core/exu_alu.v(45)
  AL_MUX \u_EXU_ALU/u969  (
    .i0(\u_EXU_ALU/n61 ),
    .i1(\u_EXU_ALU/n45 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n28 ));  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u97  (\u_EXU_ALU/n309 [8], \u_EXU_ALU/n308 [8], \u_EXU_ALU/alu_or [8]);  // ../RTL/core/exu_alu.v(66)
  AL_MUX \u_EXU_ALU/u970  (
    .i0(\u_EXU_ALU/n60 ),
    .i1(\u_EXU_ALU/n44 ),
    .sel(i_exu_op2[4]),
    .o(\u_EXU_ALU/n27 ));  // ../RTL/core/exu_alu.v(45)
  or \u_EXU_ALU/u98  (\u_EXU_ALU/n309 [9], \u_EXU_ALU/n308 [9], \u_EXU_ALU/alu_or [9]);  // ../RTL/core/exu_alu.v(66)
  or \u_EXU_ALU/u99  (\u_EXU_ALU/n309 [10], \u_EXU_ALU/n308 [10], \u_EXU_ALU/alu_or [10]);  // ../RTL/core/exu_alu.v(66)
  add_pu32_pu32_o32 \u_EXU_BJU/add0  (
    .i0(i_iaddr),
    .i1(i_imm),
    .o(\u_EXU_BJU/bxx_nxtpc ));  // ../RTL/core/exu_bju.v(57)
  add_pu30_pu30_o30 \u_EXU_BJU/add1  (
    .i0(i_iaddr[31:2]),
    .i1(30'b000000000000000000000000000001),
    .o(bju_rdwdata[31:2]));  // ../RTL/core/exu_bju.v(62)
  eq_w32 \u_EXU_BJU/eq0  (
    .i0(i_exu_op1),
    .i1(i_exu_op2),
    .o(\u_EXU_BJU/n0 ));  // ../RTL/core/exu_bju.v(42)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b0  (
    .i0(\u_EXU_BJU/bxx_nxtpc [0]),
    .i1(i_iaddr[0]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[0]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b1  (
    .i0(\u_EXU_BJU/bxx_nxtpc [1]),
    .i1(i_iaddr[1]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[1]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b10  (
    .i0(\u_EXU_BJU/bxx_nxtpc [10]),
    .i1(bju_rdwdata[10]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[10]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b11  (
    .i0(\u_EXU_BJU/bxx_nxtpc [11]),
    .i1(bju_rdwdata[11]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[11]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b12  (
    .i0(\u_EXU_BJU/bxx_nxtpc [12]),
    .i1(bju_rdwdata[12]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[12]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b13  (
    .i0(\u_EXU_BJU/bxx_nxtpc [13]),
    .i1(bju_rdwdata[13]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[13]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b14  (
    .i0(\u_EXU_BJU/bxx_nxtpc [14]),
    .i1(bju_rdwdata[14]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[14]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b15  (
    .i0(\u_EXU_BJU/bxx_nxtpc [15]),
    .i1(bju_rdwdata[15]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[15]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b16  (
    .i0(\u_EXU_BJU/bxx_nxtpc [16]),
    .i1(bju_rdwdata[16]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[16]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b17  (
    .i0(\u_EXU_BJU/bxx_nxtpc [17]),
    .i1(bju_rdwdata[17]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[17]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b18  (
    .i0(\u_EXU_BJU/bxx_nxtpc [18]),
    .i1(bju_rdwdata[18]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[18]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b19  (
    .i0(\u_EXU_BJU/bxx_nxtpc [19]),
    .i1(bju_rdwdata[19]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[19]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b2  (
    .i0(\u_EXU_BJU/bxx_nxtpc [2]),
    .i1(bju_rdwdata[2]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[2]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b20  (
    .i0(\u_EXU_BJU/bxx_nxtpc [20]),
    .i1(bju_rdwdata[20]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[20]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b21  (
    .i0(\u_EXU_BJU/bxx_nxtpc [21]),
    .i1(bju_rdwdata[21]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[21]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b22  (
    .i0(\u_EXU_BJU/bxx_nxtpc [22]),
    .i1(bju_rdwdata[22]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[22]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b23  (
    .i0(\u_EXU_BJU/bxx_nxtpc [23]),
    .i1(bju_rdwdata[23]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[23]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b24  (
    .i0(\u_EXU_BJU/bxx_nxtpc [24]),
    .i1(bju_rdwdata[24]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[24]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b25  (
    .i0(\u_EXU_BJU/bxx_nxtpc [25]),
    .i1(bju_rdwdata[25]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[25]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b26  (
    .i0(\u_EXU_BJU/bxx_nxtpc [26]),
    .i1(bju_rdwdata[26]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[26]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b27  (
    .i0(\u_EXU_BJU/bxx_nxtpc [27]),
    .i1(bju_rdwdata[27]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[27]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b28  (
    .i0(\u_EXU_BJU/bxx_nxtpc [28]),
    .i1(bju_rdwdata[28]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[28]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b29  (
    .i0(\u_EXU_BJU/bxx_nxtpc [29]),
    .i1(bju_rdwdata[29]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[29]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b3  (
    .i0(\u_EXU_BJU/bxx_nxtpc [3]),
    .i1(bju_rdwdata[3]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[3]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b30  (
    .i0(\u_EXU_BJU/bxx_nxtpc [30]),
    .i1(bju_rdwdata[30]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[30]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b31  (
    .i0(\u_EXU_BJU/bxx_nxtpc [31]),
    .i1(bju_rdwdata[31]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[31]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b4  (
    .i0(\u_EXU_BJU/bxx_nxtpc [4]),
    .i1(bju_rdwdata[4]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[4]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b5  (
    .i0(\u_EXU_BJU/bxx_nxtpc [5]),
    .i1(bju_rdwdata[5]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[5]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b6  (
    .i0(\u_EXU_BJU/bxx_nxtpc [6]),
    .i1(bju_rdwdata[6]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[6]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b7  (
    .i0(\u_EXU_BJU/bxx_nxtpc [7]),
    .i1(bju_rdwdata[7]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[7]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b8  (
    .i0(\u_EXU_BJU/bxx_nxtpc [8]),
    .i1(bju_rdwdata[8]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[8]));  // ../RTL/core/exu_bju.v(69)
  binary_mux_s1_w1 \u_EXU_BJU/mux0_b9  (
    .i0(\u_EXU_BJU/bxx_nxtpc [9]),
    .i1(bju_rdwdata[9]),
    .sel(i_decinfo[8]),
    .o(o_exu_jaddr[9]));  // ../RTL/core/exu_bju.v(69)
  ne_w32 \u_EXU_BJU/neq0  (
    .i0(i_exu_op1),
    .i1(i_exu_op2),
    .o(\u_EXU_BJU/n1 ));  // ../RTL/core/exu_bju.v(43)
  not \u_EXU_BJU/u10  (\u_EXU_BJU/n5 , \u_EXU_ALU/n261 );  // ../RTL/core/exu_bju.v(47)
  and \u_EXU_BJU/u11  (\u_EXU_BJU/bxx_bgeu , i_decinfo[7], \u_EXU_BJU/n5 );  // ../RTL/core/exu_bju.v(47)
  or \u_EXU_BJU/u12  (\u_EXU_BJU/n6 , \u_EXU_BJU/bxx_beq , \u_EXU_BJU/bxx_bne );  // ../RTL/core/exu_bju.v(49)
  or \u_EXU_BJU/u13  (\u_EXU_BJU/n7 , \u_EXU_BJU/n6 , \u_EXU_BJU/bxx_blt );  // ../RTL/core/exu_bju.v(49)
  or \u_EXU_BJU/u14  (\u_EXU_BJU/n8 , \u_EXU_BJU/n7 , \u_EXU_BJU/bxx_bge );  // ../RTL/core/exu_bju.v(49)
  or \u_EXU_BJU/u15  (\u_EXU_BJU/n9 , \u_EXU_BJU/n8 , \u_EXU_BJU/bxx_bltu );  // ../RTL/core/exu_bju.v(49)
  or \u_EXU_BJU/u16  (\u_EXU_BJU/judgeflag , \u_EXU_BJU/n9 , \u_EXU_BJU/bxx_bgeu );  // ../RTL/core/exu_bju.v(49)
  and \u_EXU_BJU/u17  (bju_rdwen, i_decinfo_grp[2], i_decinfo[1]);  // ../RTL/core/exu_bju.v(60)
  xor \u_EXU_BJU/u20  (\u_EXU_BJU/n10 , i_decinfo[8], \u_EXU_BJU/judgeflag );  // ../RTL/core/exu_bju.v(68)
  and \u_EXU_BJU/u21  (o_exu_taken, i_decinfo_grp[2], \u_EXU_BJU/n10 );  // ../RTL/core/exu_bju.v(68)
  and \u_EXU_BJU/u4  (\u_EXU_BJU/bxx_beq , i_decinfo[2], \u_EXU_BJU/n0 );  // ../RTL/core/exu_bju.v(42)
  and \u_EXU_BJU/u5  (\u_EXU_BJU/bxx_bne , i_decinfo[3], \u_EXU_BJU/n1 );  // ../RTL/core/exu_bju.v(43)
  and \u_EXU_BJU/u6  (\u_EXU_BJU/bxx_blt , i_decinfo[4], \u_EXU_ALU/n253 );  // ../RTL/core/exu_bju.v(44)
  not \u_EXU_BJU/u7  (\u_EXU_BJU/n3 , \u_EXU_ALU/n253 );  // ../RTL/core/exu_bju.v(45)
  and \u_EXU_BJU/u8  (\u_EXU_BJU/bxx_bge , i_decinfo[5], \u_EXU_BJU/n3 );  // ../RTL/core/exu_bju.v(45)
  and \u_EXU_BJU/u9  (\u_EXU_BJU/bxx_bltu , i_decinfo[6], \u_EXU_ALU/n261 );  // ../RTL/core/exu_bju.v(46)
  AL_DFF_X \u_EXU_LSU/access2_once_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n30 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/access2_once ));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/access2_vld_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n26 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/access2_vld ));  // ../RTL/core/exu_lsu.v(105)
  add_pu30_pu30_o30 \u_EXU_LSU/add0  (
    .i0(o_ribm_addr[31:2]),
    .i1(30'b000000000000000000000000000001),
    .o(\u_EXU_LSU/n59 ));  // ../RTL/core/exu_lsu.v(185)
  eq_w2 \u_EXU_LSU/eq0  (
    .i0(alu2lsu_result[1:0]),
    .i1(2'b11),
    .o(\u_EXU_LSU/n10 ));  // ../RTL/core/exu_lsu.v(121)
  AL_DFF_X \u_EXU_LSU/handshake_once_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n80 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/handshake_once ));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/handshake_rdy_last_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/handshake_rdy ),
    .en(\u_EXU_LSU/n1 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/handshake_rdy_last ));  // ../RTL/core/exu_lsu.v(73)
  not \u_EXU_LSU/lsu_finish_inv  (\u_EXU_LSU/lsu_finish_neg , \u_EXU_LSU/lsu_finish );
  not \u_EXU_LSU/lsu_vld_inv  (\u_EXU_LSU/lsu_vld_neg , \u_EXU_LSU/lsu_vld );
  not \u_EXU_LSU/lsuinfo[2]_inv  (\u_EXU_LSU/lsuinfo[2]_neg , \u_EXU_LSU/lsuinfo [2]);
  not \u_EXU_LSU/lsuinfo[3]_inv  (\u_EXU_LSU/lsuinfo[3]_neg , \u_EXU_LSU/lsuinfo [3]);
  not \u_EXU_LSU/lsuinfo[4]_inv  (\u_EXU_LSU/lsuinfo[4]_neg , \u_EXU_LSU/lsuinfo [4]);
  not \u_EXU_LSU/lsuinfo[5]_inv  (\u_EXU_LSU/lsuinfo[5]_neg , \u_EXU_LSU/lsuinfo [5]);
  and \u_EXU_LSU/mux10_b2_sel_is_2  (\u_EXU_LSU/mux10_b2_sel_is_2_o , i_rstn, \u_EXU_LSU/lsu_vld );
  and \u_EXU_LSU/mux11_b0_sel_is_2  (\u_EXU_LSU/mux11_b0_sel_is_2_o , i_rstn, \u_EXU_LSU/mux6_b0_sel_is_2_o );
  AL_MUX \u_EXU_LSU/mux12_b1  (
    .i0(1'b0),
    .i1(alu2lsu_result[0]),
    .sel(\u_EXU_LSU/mux12_b1_sel_is_1_o ),
    .o(\u_EXU_LSU/n52 [1]));
  and \u_EXU_LSU/mux12_b1_sel_is_1  (\u_EXU_LSU/mux12_b1_sel_is_1_o , i_decinfo[2], \alu2lsu_result[1]_neg );
  AL_MUX \u_EXU_LSU/mux12_b2  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n284 ),
    .sel(\u_EXU_LSU/mux12_b2_sel_is_3_o ),
    .o(\u_EXU_LSU/n52 [2]));
  and \u_EXU_LSU/mux12_b2_sel_is_3  (\u_EXU_LSU/mux12_b2_sel_is_3_o , i_decinfo[2], alu2lsu_result[1]);
  AL_MUX \u_EXU_LSU/mux12_b3  (
    .i0(1'b0),
    .i1(alu2lsu_result[0]),
    .sel(\u_EXU_LSU/mux12_b2_sel_is_3_o ),
    .o(\u_EXU_LSU/n52 [3]));
  and \u_EXU_LSU/mux13_b0_sel_is_0  (\u_EXU_LSU/mux13_b0_sel_is_0_o , \i_decinfo[3]_neg , \i_decinfo[2]_neg );
  binary_mux_s1_w1 \u_EXU_LSU/mux13_b2  (
    .i0(\u_EXU_LSU/n52 [2]),
    .i1(\u_EXU_LSU/n50 [2]),
    .sel(i_decinfo[3]),
    .o(\u_EXU_LSU/n53 [2]));  // ../RTL/core/exu_lsu.v(170)
  binary_mux_s1_w1 \u_EXU_LSU/mux13_b3  (
    .i0(\u_EXU_LSU/n52 [3]),
    .i1(alu2lsu_result[1]),
    .sel(i_decinfo[3]),
    .o(\u_EXU_LSU/n53 [3]));  // ../RTL/core/exu_lsu.v(170)
  AL_MUX \u_EXU_LSU/mux14_b0  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n284 ),
    .sel(\u_EXU_LSU/mux14_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n54 [0]));
  and \u_EXU_LSU/mux14_b0_sel_is_0  (\u_EXU_LSU/mux14_b0_sel_is_0_o , \u_EXU_LSU/mux14_b0_sel_is_2_o_neg , \alu2lsu_result[1]_neg );
  and \u_EXU_LSU/mux14_b0_sel_is_2  (\u_EXU_LSU/mux14_b0_sel_is_2_o , \i_decinfo[4]_neg , \u_EXU_LSU/mux13_b0_sel_is_0_o );
  not \u_EXU_LSU/mux14_b0_sel_is_2_o_inv  (\u_EXU_LSU/mux14_b0_sel_is_2_o_neg , \u_EXU_LSU/mux14_b0_sel_is_2_o );
  AL_MUX \u_EXU_LSU/mux14_b1  (
    .i0(\alu2lsu_result[1]_neg ),
    .i1(\u_EXU_LSU/n52 [1]),
    .sel(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .o(\u_EXU_LSU/n54 [1]));
  and \u_EXU_LSU/mux14_b1_sel_is_0  (\u_EXU_LSU/mux14_b1_sel_is_0_o , \i_decinfo[4]_neg , \i_decinfo[3]_neg );
  binary_mux_s1_w1 \u_EXU_LSU/mux14_b2  (
    .i0(\u_EXU_LSU/n53 [2]),
    .i1(\u_EXU_LSU/n49 [2]),
    .sel(i_decinfo[4]),
    .o(\u_EXU_LSU/n54 [2]));  // ../RTL/core/exu_lsu.v(169)
  binary_mux_s1_w1 \u_EXU_LSU/mux14_b3  (
    .i0(\u_EXU_LSU/n53 [3]),
    .i1(1'b1),
    .sel(i_decinfo[4]),
    .o(\u_EXU_LSU/n54 [3]));  // ../RTL/core/exu_lsu.v(169)
  binary_mux_s1_w1 \u_EXU_LSU/mux15_b2  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n63 [2]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n64 [2]));  // ../RTL/core/exu_lsu.v(191)
  AL_MUX \u_EXU_LSU/mux16_b0  (
    .i0(\u_EXU_LSU/n61 [0]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n65 [0]));
  and \u_EXU_LSU/mux16_b0_sel_is_0  (\u_EXU_LSU/mux16_b0_sel_is_0_o , \u_EXU_LSU/lsuinfo[4]_neg , \u_EXU_LSU/lsuinfo[3]_neg );
  AL_MUX \u_EXU_LSU/mux16_b1  (
    .i0(\u_EXU_LSU/align_mode_reg [1]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n65 [1]));
  binary_mux_s1_w1 \u_EXU_LSU/mux16_b2  (
    .i0(\u_EXU_LSU/n64 [2]),
    .i1(\u_EXU_LSU/n61 [2]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n65 [2]));  // ../RTL/core/exu_lsu.v(190)
  AL_MUX \u_EXU_LSU/mux16_b3  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n63 [3]),
    .sel(\u_EXU_LSU/mux16_b3_sel_is_2_o ),
    .o(\u_EXU_LSU/n65 [3]));
  and \u_EXU_LSU/mux16_b3_sel_is_2  (\u_EXU_LSU/mux16_b3_sel_is_2_o , \u_EXU_LSU/lsuinfo[4]_neg , \u_EXU_LSU/lsuinfo [3]);
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b10  (
    .i0(o_ribm_addr[10]),
    .i1(\u_EXU_LSU/n59 [8]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [10]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b11  (
    .i0(o_ribm_addr[11]),
    .i1(\u_EXU_LSU/n59 [9]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [11]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b12  (
    .i0(o_ribm_addr[12]),
    .i1(\u_EXU_LSU/n59 [10]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [12]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b13  (
    .i0(o_ribm_addr[13]),
    .i1(\u_EXU_LSU/n59 [11]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [13]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b14  (
    .i0(o_ribm_addr[14]),
    .i1(\u_EXU_LSU/n59 [12]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [14]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b15  (
    .i0(o_ribm_addr[15]),
    .i1(\u_EXU_LSU/n59 [13]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [15]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b16  (
    .i0(o_ribm_addr[16]),
    .i1(\u_EXU_LSU/n59 [14]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [16]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b17  (
    .i0(o_ribm_addr[17]),
    .i1(\u_EXU_LSU/n59 [15]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [17]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b18  (
    .i0(o_ribm_addr[18]),
    .i1(\u_EXU_LSU/n59 [16]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [18]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b19  (
    .i0(o_ribm_addr[19]),
    .i1(\u_EXU_LSU/n59 [17]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [19]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b2  (
    .i0(o_ribm_addr[2]),
    .i1(\u_EXU_LSU/n59 [0]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [2]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b20  (
    .i0(o_ribm_addr[20]),
    .i1(\u_EXU_LSU/n59 [18]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [20]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b21  (
    .i0(o_ribm_addr[21]),
    .i1(\u_EXU_LSU/n59 [19]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [21]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b22  (
    .i0(o_ribm_addr[22]),
    .i1(\u_EXU_LSU/n59 [20]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [22]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b23  (
    .i0(o_ribm_addr[23]),
    .i1(\u_EXU_LSU/n59 [21]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [23]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b24  (
    .i0(o_ribm_addr[24]),
    .i1(\u_EXU_LSU/n59 [22]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [24]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b25  (
    .i0(o_ribm_addr[25]),
    .i1(\u_EXU_LSU/n59 [23]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [25]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b26  (
    .i0(o_ribm_addr[26]),
    .i1(\u_EXU_LSU/n59 [24]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [26]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b27  (
    .i0(o_ribm_addr[27]),
    .i1(\u_EXU_LSU/n59 [25]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [27]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b28  (
    .i0(o_ribm_addr[28]),
    .i1(\u_EXU_LSU/n59 [26]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [28]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b29  (
    .i0(o_ribm_addr[29]),
    .i1(\u_EXU_LSU/n59 [27]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [29]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b3  (
    .i0(o_ribm_addr[3]),
    .i1(\u_EXU_LSU/n59 [1]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [3]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b30  (
    .i0(o_ribm_addr[30]),
    .i1(\u_EXU_LSU/n59 [28]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [30]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b31  (
    .i0(o_ribm_addr[31]),
    .i1(\u_EXU_LSU/n59 [29]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [31]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b4  (
    .i0(o_ribm_addr[4]),
    .i1(\u_EXU_LSU/n59 [2]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [4]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b5  (
    .i0(o_ribm_addr[5]),
    .i1(\u_EXU_LSU/n59 [3]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [5]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b6  (
    .i0(o_ribm_addr[6]),
    .i1(\u_EXU_LSU/n59 [4]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [6]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b7  (
    .i0(o_ribm_addr[7]),
    .i1(\u_EXU_LSU/n59 [5]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [7]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b8  (
    .i0(o_ribm_addr[8]),
    .i1(\u_EXU_LSU/n59 [6]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [8]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux17_b9  (
    .i0(o_ribm_addr[9]),
    .i1(\u_EXU_LSU/n59 [7]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n72 [9]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux18_b0  (
    .i0(o_ribm_mask[0]),
    .i1(\u_EXU_LSU/n65 [0]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n73 [0]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux18_b1  (
    .i0(o_ribm_mask[1]),
    .i1(\u_EXU_LSU/n65 [1]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n73 [1]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux18_b2  (
    .i0(o_ribm_mask[2]),
    .i1(\u_EXU_LSU/n65 [2]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n73 [2]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux18_b3  (
    .i0(o_ribm_mask[3]),
    .i1(\u_EXU_LSU/n65 [3]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n73 [3]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b0  (
    .i0(o_ribm_wdata[0]),
    .i1(\u_EXU_LSU/n67 [0]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [0]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b1  (
    .i0(o_ribm_wdata[1]),
    .i1(\u_EXU_LSU/n67 [1]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [1]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b10  (
    .i0(o_ribm_wdata[10]),
    .i1(\u_EXU_LSU/n67 [10]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [10]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b11  (
    .i0(o_ribm_wdata[11]),
    .i1(\u_EXU_LSU/n67 [11]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [11]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b12  (
    .i0(o_ribm_wdata[12]),
    .i1(\u_EXU_LSU/n67 [12]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [12]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b13  (
    .i0(o_ribm_wdata[13]),
    .i1(\u_EXU_LSU/n67 [13]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [13]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b14  (
    .i0(o_ribm_wdata[14]),
    .i1(\u_EXU_LSU/n67 [14]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [14]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b15  (
    .i0(o_ribm_wdata[15]),
    .i1(\u_EXU_LSU/n67 [15]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [15]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b16  (
    .i0(o_ribm_wdata[16]),
    .i1(\u_EXU_LSU/n67 [16]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [16]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b17  (
    .i0(o_ribm_wdata[17]),
    .i1(\u_EXU_LSU/n67 [17]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [17]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b18  (
    .i0(o_ribm_wdata[18]),
    .i1(\u_EXU_LSU/n67 [18]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [18]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b19  (
    .i0(o_ribm_wdata[19]),
    .i1(\u_EXU_LSU/n67 [19]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [19]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b2  (
    .i0(o_ribm_wdata[2]),
    .i1(\u_EXU_LSU/n67 [2]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [2]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b20  (
    .i0(o_ribm_wdata[20]),
    .i1(\u_EXU_LSU/n67 [20]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [20]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b21  (
    .i0(o_ribm_wdata[21]),
    .i1(\u_EXU_LSU/n67 [21]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [21]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b22  (
    .i0(o_ribm_wdata[22]),
    .i1(\u_EXU_LSU/n67 [22]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [22]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b23  (
    .i0(o_ribm_wdata[23]),
    .i1(\u_EXU_LSU/n67 [23]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [23]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b24  (
    .i0(o_ribm_wdata[24]),
    .i1(\u_EXU_LSU/n67 [24]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [24]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b25  (
    .i0(o_ribm_wdata[25]),
    .i1(\u_EXU_LSU/n67 [25]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [25]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b26  (
    .i0(o_ribm_wdata[26]),
    .i1(\u_EXU_LSU/n67 [26]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [26]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b27  (
    .i0(o_ribm_wdata[27]),
    .i1(\u_EXU_LSU/n67 [27]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [27]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b28  (
    .i0(o_ribm_wdata[28]),
    .i1(\u_EXU_LSU/n67 [28]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [28]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b29  (
    .i0(o_ribm_wdata[29]),
    .i1(\u_EXU_LSU/n67 [29]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [29]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b3  (
    .i0(o_ribm_wdata[3]),
    .i1(\u_EXU_LSU/n67 [3]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [3]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b30  (
    .i0(o_ribm_wdata[30]),
    .i1(\u_EXU_LSU/n67 [30]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [30]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b31  (
    .i0(o_ribm_wdata[31]),
    .i1(\u_EXU_LSU/n67 [31]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [31]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b4  (
    .i0(o_ribm_wdata[4]),
    .i1(\u_EXU_LSU/n67 [4]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [4]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b5  (
    .i0(o_ribm_wdata[5]),
    .i1(\u_EXU_LSU/n67 [5]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [5]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b6  (
    .i0(o_ribm_wdata[6]),
    .i1(\u_EXU_LSU/n67 [6]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [6]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b7  (
    .i0(o_ribm_wdata[7]),
    .i1(\u_EXU_LSU/n67 [7]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [7]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b8  (
    .i0(o_ribm_wdata[8]),
    .i1(\u_EXU_LSU/n67 [8]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [8]));  // ../RTL/core/exu_lsu.v(179)
  binary_mux_s1_w1 \u_EXU_LSU/mux19_b9  (
    .i0(o_ribm_wdata[9]),
    .i1(\u_EXU_LSU/n67 [9]),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n74 [9]));  // ../RTL/core/exu_lsu.v(179)
  and \u_EXU_LSU/mux1_b0_sel_is_2  (\u_EXU_LSU/mux1_b0_sel_is_2_o , \u_EXU_LSU/lsu_finish_neg , \u_EXU_LSU/n13 );
  and \u_EXU_LSU/mux20_b0_sel_is_0  (\u_EXU_LSU/mux20_b0_sel_is_0_o , \u_EXU_LSU/lsu_vld_neg , \u_EXU_LSU/n58_neg );
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b10  (
    .i0(\u_EXU_LSU/n72 [10]),
    .i1(alu2lsu_result[10]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [10]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b11  (
    .i0(\u_EXU_LSU/n72 [11]),
    .i1(alu2lsu_result[11]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [11]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b12  (
    .i0(\u_EXU_LSU/n72 [12]),
    .i1(alu2lsu_result[12]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [12]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b13  (
    .i0(\u_EXU_LSU/n72 [13]),
    .i1(alu2lsu_result[13]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [13]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b14  (
    .i0(\u_EXU_LSU/n72 [14]),
    .i1(alu2lsu_result[14]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [14]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b15  (
    .i0(\u_EXU_LSU/n72 [15]),
    .i1(alu2lsu_result[15]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [15]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b16  (
    .i0(\u_EXU_LSU/n72 [16]),
    .i1(alu2lsu_result[16]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [16]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b17  (
    .i0(\u_EXU_LSU/n72 [17]),
    .i1(alu2lsu_result[17]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [17]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b18  (
    .i0(\u_EXU_LSU/n72 [18]),
    .i1(alu2lsu_result[18]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [18]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b19  (
    .i0(\u_EXU_LSU/n72 [19]),
    .i1(alu2lsu_result[19]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [19]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b2  (
    .i0(\u_EXU_LSU/n72 [2]),
    .i1(alu2lsu_result[2]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [2]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b20  (
    .i0(\u_EXU_LSU/n72 [20]),
    .i1(alu2lsu_result[20]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [20]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b21  (
    .i0(\u_EXU_LSU/n72 [21]),
    .i1(alu2lsu_result[21]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [21]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b22  (
    .i0(\u_EXU_LSU/n72 [22]),
    .i1(alu2lsu_result[22]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [22]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b23  (
    .i0(\u_EXU_LSU/n72 [23]),
    .i1(alu2lsu_result[23]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [23]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b24  (
    .i0(\u_EXU_LSU/n72 [24]),
    .i1(alu2lsu_result[24]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [24]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b25  (
    .i0(\u_EXU_LSU/n72 [25]),
    .i1(alu2lsu_result[25]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [25]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b26  (
    .i0(\u_EXU_LSU/n72 [26]),
    .i1(alu2lsu_result[26]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [26]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b27  (
    .i0(\u_EXU_LSU/n72 [27]),
    .i1(alu2lsu_result[27]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [27]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b28  (
    .i0(\u_EXU_LSU/n72 [28]),
    .i1(alu2lsu_result[28]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [28]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b29  (
    .i0(\u_EXU_LSU/n72 [29]),
    .i1(alu2lsu_result[29]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [29]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b3  (
    .i0(\u_EXU_LSU/n72 [3]),
    .i1(alu2lsu_result[3]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [3]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b30  (
    .i0(\u_EXU_LSU/n72 [30]),
    .i1(alu2lsu_result[30]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [30]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b31  (
    .i0(\u_EXU_LSU/n72 [31]),
    .i1(alu2lsu_result[31]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [31]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b4  (
    .i0(\u_EXU_LSU/n72 [4]),
    .i1(alu2lsu_result[4]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [4]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b5  (
    .i0(\u_EXU_LSU/n72 [5]),
    .i1(alu2lsu_result[5]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [5]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b6  (
    .i0(\u_EXU_LSU/n72 [6]),
    .i1(alu2lsu_result[6]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [6]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b7  (
    .i0(\u_EXU_LSU/n72 [7]),
    .i1(alu2lsu_result[7]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [7]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b8  (
    .i0(\u_EXU_LSU/n72 [8]),
    .i1(alu2lsu_result[8]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [8]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux20_b9  (
    .i0(\u_EXU_LSU/n72 [9]),
    .i1(alu2lsu_result[9]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n76 [9]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux21_b0  (
    .i0(\u_EXU_LSU/n73 [0]),
    .i1(\u_EXU_LSU/n54 [0]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n78 [0]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux21_b1  (
    .i0(\u_EXU_LSU/n73 [1]),
    .i1(\u_EXU_LSU/n54 [1]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n78 [1]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux21_b2  (
    .i0(\u_EXU_LSU/n73 [2]),
    .i1(\u_EXU_LSU/n54 [2]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n78 [2]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux21_b3  (
    .i0(\u_EXU_LSU/n73 [3]),
    .i1(\u_EXU_LSU/n54 [3]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n78 [3]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b0  (
    .i0(\u_EXU_LSU/n74 [0]),
    .i1(\u_EXU_LSU/n55 [0]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [0]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b1  (
    .i0(\u_EXU_LSU/n74 [1]),
    .i1(\u_EXU_LSU/n55 [1]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [1]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b10  (
    .i0(\u_EXU_LSU/n74 [10]),
    .i1(\u_EXU_LSU/n55 [10]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [10]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b11  (
    .i0(\u_EXU_LSU/n74 [11]),
    .i1(\u_EXU_LSU/n55 [11]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [11]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b12  (
    .i0(\u_EXU_LSU/n74 [12]),
    .i1(\u_EXU_LSU/n55 [12]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [12]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b13  (
    .i0(\u_EXU_LSU/n74 [13]),
    .i1(\u_EXU_LSU/n55 [13]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [13]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b14  (
    .i0(\u_EXU_LSU/n74 [14]),
    .i1(\u_EXU_LSU/n55 [14]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [14]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b15  (
    .i0(\u_EXU_LSU/n74 [15]),
    .i1(\u_EXU_LSU/n55 [15]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [15]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b16  (
    .i0(\u_EXU_LSU/n74 [16]),
    .i1(\u_EXU_LSU/n55 [16]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [16]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b17  (
    .i0(\u_EXU_LSU/n74 [17]),
    .i1(\u_EXU_LSU/n55 [17]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [17]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b18  (
    .i0(\u_EXU_LSU/n74 [18]),
    .i1(\u_EXU_LSU/n55 [18]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [18]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b19  (
    .i0(\u_EXU_LSU/n74 [19]),
    .i1(\u_EXU_LSU/n55 [19]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [19]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b2  (
    .i0(\u_EXU_LSU/n74 [2]),
    .i1(\u_EXU_LSU/n55 [2]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [2]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b20  (
    .i0(\u_EXU_LSU/n74 [20]),
    .i1(\u_EXU_LSU/n55 [20]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [20]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b21  (
    .i0(\u_EXU_LSU/n74 [21]),
    .i1(\u_EXU_LSU/n55 [21]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [21]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b22  (
    .i0(\u_EXU_LSU/n74 [22]),
    .i1(\u_EXU_LSU/n55 [22]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [22]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b23  (
    .i0(\u_EXU_LSU/n74 [23]),
    .i1(\u_EXU_LSU/n55 [23]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [23]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b24  (
    .i0(\u_EXU_LSU/n74 [24]),
    .i1(\u_EXU_LSU/n55 [24]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [24]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b25  (
    .i0(\u_EXU_LSU/n74 [25]),
    .i1(\u_EXU_LSU/n55 [25]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [25]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b26  (
    .i0(\u_EXU_LSU/n74 [26]),
    .i1(\u_EXU_LSU/n55 [26]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [26]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b27  (
    .i0(\u_EXU_LSU/n74 [27]),
    .i1(\u_EXU_LSU/n55 [27]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [27]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b28  (
    .i0(\u_EXU_LSU/n74 [28]),
    .i1(\u_EXU_LSU/n55 [28]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [28]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b29  (
    .i0(\u_EXU_LSU/n74 [29]),
    .i1(\u_EXU_LSU/n55 [29]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [29]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b3  (
    .i0(\u_EXU_LSU/n74 [3]),
    .i1(\u_EXU_LSU/n55 [3]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [3]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b30  (
    .i0(\u_EXU_LSU/n74 [30]),
    .i1(\u_EXU_LSU/n55 [30]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [30]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b31  (
    .i0(\u_EXU_LSU/n74 [31]),
    .i1(\u_EXU_LSU/n55 [31]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [31]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b4  (
    .i0(\u_EXU_LSU/n74 [4]),
    .i1(\u_EXU_LSU/n55 [4]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [4]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b5  (
    .i0(\u_EXU_LSU/n74 [5]),
    .i1(\u_EXU_LSU/n55 [5]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [5]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b6  (
    .i0(\u_EXU_LSU/n74 [6]),
    .i1(\u_EXU_LSU/n55 [6]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [6]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b7  (
    .i0(\u_EXU_LSU/n74 [7]),
    .i1(\u_EXU_LSU/n55 [7]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [7]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b8  (
    .i0(\u_EXU_LSU/n74 [8]),
    .i1(\u_EXU_LSU/n55 [8]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [8]));  // ../RTL/core/exu_lsu.v(160)
  binary_mux_s1_w1 \u_EXU_LSU/mux22_b9  (
    .i0(\u_EXU_LSU/n74 [9]),
    .i1(\u_EXU_LSU/n55 [9]),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n79 [9]));  // ../RTL/core/exu_lsu.v(160)
  AL_MUX \u_EXU_LSU/mux27_b16  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/access2_data [15]),
    .sel(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .o(\u_EXU_LSU/n136 [16]));
  and \u_EXU_LSU/mux27_b16_sel_is_1  (\u_EXU_LSU/mux27_b16_sel_is_1_o , \u_EXU_LSU/lsuinfo [3], \u_EXU_LSU/lsuinfo[5]_neg );
  AL_MUX \u_EXU_LSU/mux28_b0  (
    .i0(\u_EXU_LSU/access2_data [0]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [0]));
  AL_MUX \u_EXU_LSU/mux28_b1  (
    .i0(\u_EXU_LSU/access2_data [1]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [1]));
  AL_MUX \u_EXU_LSU/mux28_b10  (
    .i0(\u_EXU_LSU/access2_data [10]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [10]));
  AL_MUX \u_EXU_LSU/mux28_b11  (
    .i0(\u_EXU_LSU/access2_data [11]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [11]));
  AL_MUX \u_EXU_LSU/mux28_b12  (
    .i0(\u_EXU_LSU/access2_data [12]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [12]));
  AL_MUX \u_EXU_LSU/mux28_b13  (
    .i0(\u_EXU_LSU/access2_data [13]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [13]));
  AL_MUX \u_EXU_LSU/mux28_b14  (
    .i0(\u_EXU_LSU/access2_data [14]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [14]));
  AL_MUX \u_EXU_LSU/mux28_b15  (
    .i0(\u_EXU_LSU/access2_data [15]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [15]));
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b16  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [16]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [16]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b17  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [17]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [17]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b18  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [18]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [18]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b19  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [19]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [19]));  // ../RTL/core/exu_lsu.v(215)
  AL_MUX \u_EXU_LSU/mux28_b2  (
    .i0(\u_EXU_LSU/access2_data [2]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [2]));
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b20  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [20]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [20]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b21  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [21]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [21]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b22  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [22]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [22]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b23  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [23]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [23]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b24  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [24]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [24]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b25  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [25]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [25]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b26  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [26]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [26]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b27  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [27]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [27]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b28  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [28]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [28]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b29  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [29]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [29]));  // ../RTL/core/exu_lsu.v(215)
  AL_MUX \u_EXU_LSU/mux28_b3  (
    .i0(\u_EXU_LSU/access2_data [3]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [3]));
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b30  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [30]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [30]));  // ../RTL/core/exu_lsu.v(215)
  binary_mux_s1_w1 \u_EXU_LSU/mux28_b31  (
    .i0(\u_EXU_LSU/n136 [16]),
    .i1(\u_EXU_LSU/access2_data [31]),
    .sel(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n137 [31]));  // ../RTL/core/exu_lsu.v(215)
  AL_MUX \u_EXU_LSU/mux28_b4  (
    .i0(\u_EXU_LSU/access2_data [4]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [4]));
  AL_MUX \u_EXU_LSU/mux28_b5  (
    .i0(\u_EXU_LSU/access2_data [5]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [5]));
  AL_MUX \u_EXU_LSU/mux28_b6  (
    .i0(\u_EXU_LSU/access2_data [6]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [6]));
  AL_MUX \u_EXU_LSU/mux28_b7  (
    .i0(\u_EXU_LSU/access2_data [7]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [7]));
  AL_MUX \u_EXU_LSU/mux28_b8  (
    .i0(\u_EXU_LSU/access2_data [8]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [8]));
  AL_MUX \u_EXU_LSU/mux28_b9  (
    .i0(\u_EXU_LSU/access2_data [9]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/mux16_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n137 [9]));
  binary_mux_s1_w1 \u_EXU_LSU/mux29_b0  (
    .i0(\u_EXU_LSU/access_data [15]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/lsuinfo [5]),
    .o(\u_EXU_LSU/n138 [0]));  // ../RTL/core/exu_lsu.v(222)
  binary_mux_s1_w1 \u_EXU_LSU/mux30_b0  (
    .i0(\u_EXU_LSU/access2_data [39]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/lsuinfo [5]),
    .o(\u_EXU_LSU/n139 [0]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b10  (
    .i0(i_ribm_rdata[10]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [10]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b11  (
    .i0(i_ribm_rdata[11]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [11]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b12  (
    .i0(i_ribm_rdata[12]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [12]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b13  (
    .i0(i_ribm_rdata[13]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [13]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b14  (
    .i0(i_ribm_rdata[14]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [14]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b15  (
    .i0(i_ribm_rdata[15]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [15]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b16  (
    .i0(i_ribm_rdata[16]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [16]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b17  (
    .i0(i_ribm_rdata[17]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [17]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b18  (
    .i0(i_ribm_rdata[18]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [18]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b19  (
    .i0(i_ribm_rdata[19]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [19]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b20  (
    .i0(i_ribm_rdata[20]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [20]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b21  (
    .i0(i_ribm_rdata[21]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [21]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b22  (
    .i0(i_ribm_rdata[22]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [22]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b23  (
    .i0(i_ribm_rdata[23]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [23]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b24  (
    .i0(i_ribm_rdata[24]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [24]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b25  (
    .i0(i_ribm_rdata[25]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [25]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b26  (
    .i0(i_ribm_rdata[26]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [26]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b27  (
    .i0(i_ribm_rdata[27]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [27]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b28  (
    .i0(i_ribm_rdata[28]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [28]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b29  (
    .i0(i_ribm_rdata[29]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [29]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b30  (
    .i0(i_ribm_rdata[30]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [30]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b31  (
    .i0(i_ribm_rdata[31]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [31]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b8  (
    .i0(i_ribm_rdata[8]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [8]));  // ../RTL/core/exu_lsu.v(223)
  binary_mux_s1_w1 \u_EXU_LSU/mux31_b9  (
    .i0(i_ribm_rdata[9]),
    .i1(\u_EXU_LSU/n139 [0]),
    .sel(\u_EXU_LSU/lsuinfo [2]),
    .o(\u_EXU_LSU/n140 [9]));  // ../RTL/core/exu_lsu.v(223)
  AL_MUX \u_EXU_LSU/mux32_b0  (
    .i0(\u_EXU_LSU/access2_data [32]),
    .i1(i_ribm_rdata[0]),
    .sel(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n141 [0]));
  and \u_EXU_LSU/mux32_b0_sel_is_0  (\u_EXU_LSU/mux32_b0_sel_is_0_o , \u_EXU_LSU/lsuinfo[3]_neg , \u_EXU_LSU/lsuinfo[2]_neg );
  AL_MUX \u_EXU_LSU/mux32_b1  (
    .i0(\u_EXU_LSU/access2_data [33]),
    .i1(i_ribm_rdata[1]),
    .sel(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n141 [1]));
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b10  (
    .i0(\u_EXU_LSU/n140 [10]),
    .i1(\u_EXU_LSU/access2_data [42]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [10]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b11  (
    .i0(\u_EXU_LSU/n140 [11]),
    .i1(\u_EXU_LSU/access2_data [43]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [11]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b12  (
    .i0(\u_EXU_LSU/n140 [12]),
    .i1(\u_EXU_LSU/access_data [12]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [12]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b13  (
    .i0(\u_EXU_LSU/n140 [13]),
    .i1(\u_EXU_LSU/access_data [13]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [13]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b14  (
    .i0(\u_EXU_LSU/n140 [14]),
    .i1(\u_EXU_LSU/access_data [14]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [14]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b15  (
    .i0(\u_EXU_LSU/n140 [15]),
    .i1(\u_EXU_LSU/access_data [15]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [15]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b16  (
    .i0(\u_EXU_LSU/n140 [16]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [16]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b17  (
    .i0(\u_EXU_LSU/n140 [17]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [17]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b18  (
    .i0(\u_EXU_LSU/n140 [18]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [18]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b19  (
    .i0(\u_EXU_LSU/n140 [19]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [19]));  // ../RTL/core/exu_lsu.v(221)
  AL_MUX \u_EXU_LSU/mux32_b2  (
    .i0(\u_EXU_LSU/access2_data [34]),
    .i1(i_ribm_rdata[2]),
    .sel(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n141 [2]));
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b20  (
    .i0(\u_EXU_LSU/n140 [20]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [20]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b21  (
    .i0(\u_EXU_LSU/n140 [21]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [21]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b22  (
    .i0(\u_EXU_LSU/n140 [22]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [22]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b23  (
    .i0(\u_EXU_LSU/n140 [23]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [23]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b24  (
    .i0(\u_EXU_LSU/n140 [24]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [24]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b25  (
    .i0(\u_EXU_LSU/n140 [25]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [25]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b26  (
    .i0(\u_EXU_LSU/n140 [26]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [26]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b27  (
    .i0(\u_EXU_LSU/n140 [27]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [27]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b28  (
    .i0(\u_EXU_LSU/n140 [28]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [28]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b29  (
    .i0(\u_EXU_LSU/n140 [29]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [29]));  // ../RTL/core/exu_lsu.v(221)
  AL_MUX \u_EXU_LSU/mux32_b3  (
    .i0(\u_EXU_LSU/access2_data [35]),
    .i1(i_ribm_rdata[3]),
    .sel(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n141 [3]));
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b30  (
    .i0(\u_EXU_LSU/n140 [30]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [30]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b31  (
    .i0(\u_EXU_LSU/n140 [31]),
    .i1(\u_EXU_LSU/n138 [0]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [31]));  // ../RTL/core/exu_lsu.v(221)
  AL_MUX \u_EXU_LSU/mux32_b4  (
    .i0(\u_EXU_LSU/access2_data [36]),
    .i1(i_ribm_rdata[4]),
    .sel(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n141 [4]));
  AL_MUX \u_EXU_LSU/mux32_b5  (
    .i0(\u_EXU_LSU/access2_data [37]),
    .i1(i_ribm_rdata[5]),
    .sel(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n141 [5]));
  AL_MUX \u_EXU_LSU/mux32_b6  (
    .i0(\u_EXU_LSU/access2_data [38]),
    .i1(i_ribm_rdata[6]),
    .sel(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n141 [6]));
  AL_MUX \u_EXU_LSU/mux32_b7  (
    .i0(\u_EXU_LSU/access2_data [39]),
    .i1(i_ribm_rdata[7]),
    .sel(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n141 [7]));
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b8  (
    .i0(\u_EXU_LSU/n140 [8]),
    .i1(\u_EXU_LSU/access2_data [40]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [8]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux32_b9  (
    .i0(\u_EXU_LSU/n140 [9]),
    .i1(\u_EXU_LSU/access2_data [41]),
    .sel(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/n141 [9]));  // ../RTL/core/exu_lsu.v(221)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b0  (
    .i0(\u_EXU_LSU/n141 [0]),
    .i1(\u_EXU_LSU/n137 [0]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[0]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b1  (
    .i0(\u_EXU_LSU/n141 [1]),
    .i1(\u_EXU_LSU/n137 [1]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[1]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b10  (
    .i0(\u_EXU_LSU/n141 [10]),
    .i1(\u_EXU_LSU/n137 [10]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[10]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b11  (
    .i0(\u_EXU_LSU/n141 [11]),
    .i1(\u_EXU_LSU/n137 [11]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[11]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b12  (
    .i0(\u_EXU_LSU/n141 [12]),
    .i1(\u_EXU_LSU/n137 [12]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[12]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b13  (
    .i0(\u_EXU_LSU/n141 [13]),
    .i1(\u_EXU_LSU/n137 [13]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[13]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b14  (
    .i0(\u_EXU_LSU/n141 [14]),
    .i1(\u_EXU_LSU/n137 [14]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[14]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b15  (
    .i0(\u_EXU_LSU/n141 [15]),
    .i1(\u_EXU_LSU/n137 [15]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[15]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b16  (
    .i0(\u_EXU_LSU/n141 [16]),
    .i1(\u_EXU_LSU/n137 [16]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[16]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b17  (
    .i0(\u_EXU_LSU/n141 [17]),
    .i1(\u_EXU_LSU/n137 [17]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[17]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b18  (
    .i0(\u_EXU_LSU/n141 [18]),
    .i1(\u_EXU_LSU/n137 [18]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[18]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b19  (
    .i0(\u_EXU_LSU/n141 [19]),
    .i1(\u_EXU_LSU/n137 [19]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[19]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b2  (
    .i0(\u_EXU_LSU/n141 [2]),
    .i1(\u_EXU_LSU/n137 [2]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[2]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b20  (
    .i0(\u_EXU_LSU/n141 [20]),
    .i1(\u_EXU_LSU/n137 [20]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[20]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b21  (
    .i0(\u_EXU_LSU/n141 [21]),
    .i1(\u_EXU_LSU/n137 [21]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[21]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b22  (
    .i0(\u_EXU_LSU/n141 [22]),
    .i1(\u_EXU_LSU/n137 [22]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[22]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b23  (
    .i0(\u_EXU_LSU/n141 [23]),
    .i1(\u_EXU_LSU/n137 [23]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[23]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b24  (
    .i0(\u_EXU_LSU/n141 [24]),
    .i1(\u_EXU_LSU/n137 [24]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[24]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b25  (
    .i0(\u_EXU_LSU/n141 [25]),
    .i1(\u_EXU_LSU/n137 [25]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[25]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b26  (
    .i0(\u_EXU_LSU/n141 [26]),
    .i1(\u_EXU_LSU/n137 [26]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[26]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b27  (
    .i0(\u_EXU_LSU/n141 [27]),
    .i1(\u_EXU_LSU/n137 [27]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[27]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b28  (
    .i0(\u_EXU_LSU/n141 [28]),
    .i1(\u_EXU_LSU/n137 [28]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[28]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b29  (
    .i0(\u_EXU_LSU/n141 [29]),
    .i1(\u_EXU_LSU/n137 [29]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[29]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b3  (
    .i0(\u_EXU_LSU/n141 [3]),
    .i1(\u_EXU_LSU/n137 [3]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[3]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b30  (
    .i0(\u_EXU_LSU/n141 [30]),
    .i1(\u_EXU_LSU/n137 [30]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[30]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b31  (
    .i0(\u_EXU_LSU/n141 [31]),
    .i1(\u_EXU_LSU/n137 [31]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[31]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b4  (
    .i0(\u_EXU_LSU/n141 [4]),
    .i1(\u_EXU_LSU/n137 [4]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[4]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b5  (
    .i0(\u_EXU_LSU/n141 [5]),
    .i1(\u_EXU_LSU/n137 [5]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[5]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b6  (
    .i0(\u_EXU_LSU/n141 [6]),
    .i1(\u_EXU_LSU/n137 [6]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[6]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b7  (
    .i0(\u_EXU_LSU/n141 [7]),
    .i1(\u_EXU_LSU/n137 [7]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[7]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b8  (
    .i0(\u_EXU_LSU/n141 [8]),
    .i1(\u_EXU_LSU/n137 [8]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[8]));  // ../RTL/core/exu_lsu.v(214)
  binary_mux_s1_w1 \u_EXU_LSU/mux33_b9  (
    .i0(\u_EXU_LSU/n141 [9]),
    .i1(\u_EXU_LSU/n137 [9]),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[9]));  // ../RTL/core/exu_lsu.v(214)
  and \u_EXU_LSU/mux6_b0_sel_is_2  (\u_EXU_LSU/mux6_b0_sel_is_2_o , \u_EXU_LSU/lsu_vld_neg , \u_EXU_LSU/mux1_b0_sel_is_2_o );
  not \u_EXU_LSU/n13_inv  (\u_EXU_LSU/n13_neg , \u_EXU_LSU/n13 );
  not \u_EXU_LSU/n58_inv  (\u_EXU_LSU/n58_neg , \u_EXU_LSU/n58 );
  not \u_EXU_LSU/n66[1]_inv  (\u_EXU_LSU/n66[1]_neg , \u_EXU_LSU/n66 [1]);
  ne_w2 \u_EXU_LSU/neq0  (
    .i0(alu2lsu_result[1:0]),
    .i1(2'b00),
    .o(\u_EXU_LSU/n9 ));  // ../RTL/core/exu_lsu.v(120)
  AL_DFF_X \u_EXU_LSU/o_ribm_req_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n75 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_req));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/o_ribm_wrcs_reg  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_decinfo[1]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wrcs));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/rdwen_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n23 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_exu_rdwen2));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg0_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_rdidx0[0]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_rdidx2[0]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg0_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_rdidx0[1]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_rdidx2[1]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg0_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_rdidx0[2]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_rdidx2[2]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg0_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_rdidx0[3]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_rdidx2[3]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg0_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(o_rdidx0[4]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_rdidx2[4]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg1_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(alu2lsu_result[0]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/align_mode_reg [0]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg1_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(alu2lsu_result[1]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/align_mode_reg [1]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[0]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [0]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[1]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [1]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[10]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [10]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[11]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [11]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[12]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [12]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[13]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [13]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[14]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [14]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[15]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [15]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[16]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [16]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[17]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [17]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[18]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [18]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[19]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [19]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[2]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [2]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[20]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [20]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[21]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [21]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[22]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [22]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[23]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [23]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[24]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [24]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[25]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [25]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[26]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [26]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[27]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [27]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[28]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [28]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[29]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [29]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[3]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [3]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[30]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [30]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[31]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [31]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[4]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [4]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[5]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [5]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[6]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [6]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[7]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [7]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[8]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [8]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg2_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rs2rdata[9]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/rs2rdata_reg [9]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg3_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_decinfo[2]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/lsuinfo [2]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg3_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_decinfo[3]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/lsuinfo [3]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg3_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_decinfo[4]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/lsuinfo [4]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg3_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_decinfo[5]),
    .en(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/lsuinfo [5]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[0]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [0]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[1]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [1]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[10]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [10]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[11]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [11]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[12]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [12]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[13]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [13]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[14]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [14]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[15]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [15]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[16]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [16]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[17]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [17]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[18]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [18]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[19]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [19]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[2]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [2]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[20]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [20]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[21]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [21]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[22]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [22]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[23]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [23]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[24]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [24]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[25]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [25]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[26]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [26]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[27]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [27]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[28]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [28]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[29]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [29]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[3]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [3]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[30]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [30]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[31]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [31]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[4]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [4]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[5]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [5]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[6]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [6]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[7]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [7]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[8]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [8]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg4_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_ribm_rdata[9]),
    .en(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/overleft_buffer [9]));  // ../RTL/core/exu_lsu.v(105)
  AL_DFF_X \u_EXU_LSU/reg5_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [10]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[10]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [11]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[11]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [12]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[12]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [13]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[13]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [14]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[14]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [15]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[15]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [16]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[16]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [17]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[17]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [18]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[18]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [19]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[19]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [2]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[2]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [20]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[20]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [21]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[21]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [22]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[22]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [23]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[23]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [24]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[24]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [25]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[25]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [26]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[26]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [27]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[27]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [28]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[28]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [29]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[29]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [3]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[3]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [30]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[30]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [31]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[31]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [4]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[4]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [5]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[5]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [6]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[6]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [7]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[7]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [8]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[8]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg5_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [9]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_addr[9]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg6_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n78 [0]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_mask[0]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg6_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n78 [1]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_mask[1]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg6_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n78 [2]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_mask[2]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg6_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n78 [3]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_mask[3]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [0]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[0]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b1  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [1]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[1]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [10]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[10]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b11  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [11]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[11]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b12  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [12]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[12]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b13  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [13]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[13]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b14  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [14]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[14]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b15  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [15]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[15]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b16  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [16]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[16]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b17  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [17]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[17]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b18  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [18]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[18]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b19  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [19]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[19]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b2  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [2]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[2]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [20]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[20]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b21  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [21]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[21]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b22  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [22]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[22]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b23  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [23]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[23]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b24  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [24]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[24]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b25  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [25]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[25]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b26  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [26]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[26]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b27  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [27]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[27]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b28  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [28]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[28]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b29  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [29]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[29]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b3  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [3]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[3]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [30]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[30]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b31  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [31]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[31]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b4  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [4]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[4]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b5  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [5]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[5]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b6  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [6]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[6]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b7  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [7]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[7]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b8  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [8]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[8]));  // ../RTL/core/exu_lsu.v(156)
  AL_DFF_X \u_EXU_LSU/reg7_b9  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [9]),
    .en(i_rstn),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_ribm_wdata[9]));  // ../RTL/core/exu_lsu.v(156)
  add_pu2_mu2_o3 \u_EXU_LSU/sub0_2  (
    .i0(2'b00),
    .i1(\u_EXU_LSU/align_mode_reg ),
    .o({\u_EXU_LSU/sub0_2_co ,\u_EXU_LSU/n66 [1:0]}));  // ../RTL/core/exu_lsu.v(194)
  not \u_EXU_LSU/sub0_2_co_inv  (\u_EXU_LSU/sub0_2_co_neg , \u_EXU_LSU/sub0_2_co );
  not \u_EXU_LSU/u10  (\u_EXU_LSU/n3 , o_lsu_working);  // ../RTL/core/exu_lsu.v(101)
  AL_MUX \u_EXU_LSU/u100  (
    .i0(\u_EXU_LSU/n101 ),
    .i1(\u_EXU_LSU/n178 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access_data [12]));  // ../RTL/core/exu_lsu.v(210)
  AL_MUX \u_EXU_LSU/u101  (
    .i0(\u_EXU_LSU/n100 ),
    .i1(\u_EXU_LSU/n179 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access_data [13]));  // ../RTL/core/exu_lsu.v(210)
  AL_MUX \u_EXU_LSU/u102  (
    .i0(\u_EXU_LSU/n99 ),
    .i1(\u_EXU_LSU/n180 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access_data [14]));  // ../RTL/core/exu_lsu.v(210)
  AL_MUX \u_EXU_LSU/u103  (
    .i0(\u_EXU_LSU/n98 ),
    .i1(\u_EXU_LSU/n181 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access_data [15]));  // ../RTL/core/exu_lsu.v(210)
  and \u_EXU_LSU/u11  (\u_EXU_LSU/n4 , i_decinfo_grp[1], \u_EXU_LSU/n3 );  // ../RTL/core/exu_lsu.v(101)
  and \u_EXU_LSU/u12  (\u_EXU_LSU/lsu_vld , \u_EXU_LSU/n4 , i_vld);  // ../RTL/core/exu_lsu.v(101)
  AL_MUX \u_EXU_LSU/u120  (
    .i0(\u_EXU_LSU/overleft_buffer [0]),
    .i1(\u_EXU_LSU/overleft_buffer [8]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n91 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u121  (
    .i0(\u_EXU_LSU/overleft_buffer [1]),
    .i1(\u_EXU_LSU/overleft_buffer [9]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n90 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u122  (
    .i0(\u_EXU_LSU/overleft_buffer [2]),
    .i1(\u_EXU_LSU/overleft_buffer [10]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n89 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u123  (
    .i0(\u_EXU_LSU/overleft_buffer [3]),
    .i1(\u_EXU_LSU/overleft_buffer [11]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n88 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u124  (
    .i0(\u_EXU_LSU/overleft_buffer [4]),
    .i1(\u_EXU_LSU/overleft_buffer [12]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n87 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u125  (
    .i0(\u_EXU_LSU/overleft_buffer [5]),
    .i1(\u_EXU_LSU/overleft_buffer [13]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n86 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u126  (
    .i0(\u_EXU_LSU/overleft_buffer [6]),
    .i1(\u_EXU_LSU/overleft_buffer [14]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n85 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u127  (
    .i0(\u_EXU_LSU/overleft_buffer [7]),
    .i1(\u_EXU_LSU/overleft_buffer [15]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n84 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u128  (
    .i0(\u_EXU_LSU/overleft_buffer [8]),
    .i1(\u_EXU_LSU/overleft_buffer [16]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n83 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u129  (
    .i0(\u_EXU_LSU/overleft_buffer [9]),
    .i1(\u_EXU_LSU/overleft_buffer [17]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n82 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u13  (
    .i0(1'b1),
    .i1(\u_EXU_LSU/access2_once ),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(\u_EXU_LSU/n5 ));  // ../RTL/core/exu_lsu.v(103)
  AL_MUX \u_EXU_LSU/u130  (
    .i0(\u_EXU_LSU/overleft_buffer [10]),
    .i1(\u_EXU_LSU/overleft_buffer [18]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n81 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u131  (
    .i0(\u_EXU_LSU/overleft_buffer [11]),
    .i1(\u_EXU_LSU/overleft_buffer [19]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n173 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u132  (
    .i0(\u_EXU_LSU/overleft_buffer [12]),
    .i1(\u_EXU_LSU/overleft_buffer [20]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n172 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u133  (
    .i0(\u_EXU_LSU/overleft_buffer [13]),
    .i1(\u_EXU_LSU/overleft_buffer [21]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n171 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u134  (
    .i0(\u_EXU_LSU/overleft_buffer [14]),
    .i1(\u_EXU_LSU/overleft_buffer [22]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n170 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u135  (
    .i0(\u_EXU_LSU/overleft_buffer [15]),
    .i1(\u_EXU_LSU/overleft_buffer [23]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n169 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u136  (
    .i0(\u_EXU_LSU/overleft_buffer [16]),
    .i1(\u_EXU_LSU/overleft_buffer [24]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n168 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u137  (
    .i0(\u_EXU_LSU/overleft_buffer [17]),
    .i1(\u_EXU_LSU/overleft_buffer [25]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n167 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u138  (
    .i0(\u_EXU_LSU/overleft_buffer [18]),
    .i1(\u_EXU_LSU/overleft_buffer [26]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n166 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u139  (
    .i0(\u_EXU_LSU/overleft_buffer [19]),
    .i1(\u_EXU_LSU/overleft_buffer [27]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n165 ));  // ../RTL/core/exu_lsu.v(209)
  not \u_EXU_LSU/u14  (\u_EXU_LSU/n7 , i_decinfo[1]);  // ../RTL/core/exu_lsu.v(113)
  AL_MUX \u_EXU_LSU/u140  (
    .i0(\u_EXU_LSU/overleft_buffer [20]),
    .i1(\u_EXU_LSU/overleft_buffer [28]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n164 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u141  (
    .i0(\u_EXU_LSU/overleft_buffer [21]),
    .i1(\u_EXU_LSU/overleft_buffer [29]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n163 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u142  (
    .i0(\u_EXU_LSU/overleft_buffer [22]),
    .i1(\u_EXU_LSU/overleft_buffer [30]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n162 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u143  (
    .i0(\u_EXU_LSU/overleft_buffer [23]),
    .i1(\u_EXU_LSU/overleft_buffer [31]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n161 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u144  (
    .i0(\u_EXU_LSU/overleft_buffer [24]),
    .i1(i_ribm_rdata[0]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n160 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u145  (
    .i0(\u_EXU_LSU/overleft_buffer [25]),
    .i1(i_ribm_rdata[1]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n159 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u146  (
    .i0(\u_EXU_LSU/overleft_buffer [26]),
    .i1(i_ribm_rdata[2]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n158 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u147  (
    .i0(\u_EXU_LSU/overleft_buffer [27]),
    .i1(i_ribm_rdata[3]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n157 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u148  (
    .i0(\u_EXU_LSU/overleft_buffer [28]),
    .i1(i_ribm_rdata[4]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n156 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u149  (
    .i0(\u_EXU_LSU/overleft_buffer [29]),
    .i1(i_ribm_rdata[5]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n155 ));  // ../RTL/core/exu_lsu.v(209)
  and \u_EXU_LSU/u15  (\u_EXU_LSU/n8 , \u_EXU_LSU/n7 , o_exu_rdwen0);  // ../RTL/core/exu_lsu.v(113)
  AL_MUX \u_EXU_LSU/u150  (
    .i0(\u_EXU_LSU/overleft_buffer [30]),
    .i1(i_ribm_rdata[6]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n154 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u151  (
    .i0(\u_EXU_LSU/overleft_buffer [31]),
    .i1(i_ribm_rdata[7]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n153 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u152  (
    .i0(i_ribm_rdata[0]),
    .i1(i_ribm_rdata[8]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n152 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u153  (
    .i0(i_ribm_rdata[1]),
    .i1(i_ribm_rdata[9]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n151 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u154  (
    .i0(i_ribm_rdata[2]),
    .i1(i_ribm_rdata[10]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n150 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u155  (
    .i0(i_ribm_rdata[3]),
    .i1(i_ribm_rdata[11]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n149 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u156  (
    .i0(i_ribm_rdata[4]),
    .i1(i_ribm_rdata[12]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n148 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u157  (
    .i0(i_ribm_rdata[5]),
    .i1(i_ribm_rdata[13]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n147 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u158  (
    .i0(i_ribm_rdata[6]),
    .i1(i_ribm_rdata[14]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n146 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u159  (
    .i0(i_ribm_rdata[7]),
    .i1(i_ribm_rdata[15]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n145 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u16  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n10 ),
    .sel(i_decinfo[3]),
    .o(\u_EXU_LSU/n11 ));  // ../RTL/core/exu_lsu.v(121)
  AL_MUX \u_EXU_LSU/u160  (
    .i0(i_ribm_rdata[8]),
    .i1(i_ribm_rdata[16]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n144 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u161  (
    .i0(i_ribm_rdata[9]),
    .i1(i_ribm_rdata[17]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n143 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u162  (
    .i0(i_ribm_rdata[10]),
    .i1(i_ribm_rdata[18]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n142 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u163  (
    .i0(i_ribm_rdata[11]),
    .i1(i_ribm_rdata[19]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n102 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u164  (
    .i0(i_ribm_rdata[12]),
    .i1(i_ribm_rdata[20]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n101 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u165  (
    .i0(i_ribm_rdata[13]),
    .i1(i_ribm_rdata[21]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n100 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u166  (
    .i0(i_ribm_rdata[14]),
    .i1(i_ribm_rdata[22]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n99 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u167  (
    .i0(i_ribm_rdata[15]),
    .i1(i_ribm_rdata[23]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n98 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u168  (
    .i0(i_ribm_rdata[16]),
    .i1(i_ribm_rdata[24]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n97 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u169  (
    .i0(i_ribm_rdata[17]),
    .i1(i_ribm_rdata[25]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n48 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u17  (
    .i0(\u_EXU_LSU/n11 ),
    .i1(\u_EXU_LSU/n9 ),
    .sel(i_decinfo[4]),
    .o(\u_EXU_LSU/n12 ));  // ../RTL/core/exu_lsu.v(120)
  AL_MUX \u_EXU_LSU/u170  (
    .i0(i_ribm_rdata[18]),
    .i1(i_ribm_rdata[26]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n47 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u171  (
    .i0(i_ribm_rdata[19]),
    .i1(i_ribm_rdata[27]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n46 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u172  (
    .i0(i_ribm_rdata[20]),
    .i1(i_ribm_rdata[28]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n45 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u173  (
    .i0(i_ribm_rdata[21]),
    .i1(i_ribm_rdata[29]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n44 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u174  (
    .i0(i_ribm_rdata[22]),
    .i1(i_ribm_rdata[30]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n43 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u175  (
    .i0(i_ribm_rdata[23]),
    .i1(i_ribm_rdata[31]),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n42 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u176  (
    .i0(i_ribm_rdata[24]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n174 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u177  (
    .i0(i_ribm_rdata[25]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n175 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u178  (
    .i0(i_ribm_rdata[26]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n176 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u179  (
    .i0(i_ribm_rdata[27]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n177 ));  // ../RTL/core/exu_lsu.v(209)
  and \u_EXU_LSU/u18  (\u_EXU_LSU/n13 , \u_EXU_LSU/access2_vld , \u_EXU_LSU/trans_finish );  // ../RTL/core/exu_lsu.v(135)
  AL_MUX \u_EXU_LSU/u180  (
    .i0(i_ribm_rdata[28]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n178 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u181  (
    .i0(i_ribm_rdata[29]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n179 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u182  (
    .i0(i_ribm_rdata[30]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n180 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u183  (
    .i0(i_ribm_rdata[31]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/n181 ));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u184  (
    .i0(\u_EXU_LSU/n91 ),
    .i1(\u_EXU_LSU/n168 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [0]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u185  (
    .i0(\u_EXU_LSU/n90 ),
    .i1(\u_EXU_LSU/n167 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [1]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u186  (
    .i0(\u_EXU_LSU/n89 ),
    .i1(\u_EXU_LSU/n166 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [2]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u187  (
    .i0(\u_EXU_LSU/n88 ),
    .i1(\u_EXU_LSU/n165 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [3]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u188  (
    .i0(\u_EXU_LSU/n87 ),
    .i1(\u_EXU_LSU/n164 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [4]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u189  (
    .i0(\u_EXU_LSU/n86 ),
    .i1(\u_EXU_LSU/n163 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [5]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u190  (
    .i0(\u_EXU_LSU/n85 ),
    .i1(\u_EXU_LSU/n162 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [6]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u191  (
    .i0(\u_EXU_LSU/n84 ),
    .i1(\u_EXU_LSU/n161 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [7]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u192  (
    .i0(\u_EXU_LSU/n83 ),
    .i1(\u_EXU_LSU/n160 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [8]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u193  (
    .i0(\u_EXU_LSU/n82 ),
    .i1(\u_EXU_LSU/n159 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [9]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u194  (
    .i0(\u_EXU_LSU/n81 ),
    .i1(\u_EXU_LSU/n158 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [10]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u195  (
    .i0(\u_EXU_LSU/n173 ),
    .i1(\u_EXU_LSU/n157 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [11]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u196  (
    .i0(\u_EXU_LSU/n172 ),
    .i1(\u_EXU_LSU/n156 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [12]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u197  (
    .i0(\u_EXU_LSU/n171 ),
    .i1(\u_EXU_LSU/n155 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [13]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u198  (
    .i0(\u_EXU_LSU/n170 ),
    .i1(\u_EXU_LSU/n154 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [14]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u199  (
    .i0(\u_EXU_LSU/n169 ),
    .i1(\u_EXU_LSU/n153 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [15]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u20  (
    .i0(\u_EXU_LSU/access2_once ),
    .i1(1'b1),
    .sel(\u_EXU_LSU/n13 ),
    .o(\u_EXU_LSU/n16 ));  // ../RTL/core/exu_lsu.v(135)
  AL_MUX \u_EXU_LSU/u200  (
    .i0(\u_EXU_LSU/n168 ),
    .i1(\u_EXU_LSU/n152 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [16]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u201  (
    .i0(\u_EXU_LSU/n167 ),
    .i1(\u_EXU_LSU/n151 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [17]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u202  (
    .i0(\u_EXU_LSU/n166 ),
    .i1(\u_EXU_LSU/n150 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [18]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u203  (
    .i0(\u_EXU_LSU/n165 ),
    .i1(\u_EXU_LSU/n149 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [19]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u204  (
    .i0(\u_EXU_LSU/n164 ),
    .i1(\u_EXU_LSU/n148 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [20]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u205  (
    .i0(\u_EXU_LSU/n163 ),
    .i1(\u_EXU_LSU/n147 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [21]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u206  (
    .i0(\u_EXU_LSU/n162 ),
    .i1(\u_EXU_LSU/n146 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [22]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u207  (
    .i0(\u_EXU_LSU/n161 ),
    .i1(\u_EXU_LSU/n145 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [23]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u208  (
    .i0(\u_EXU_LSU/n160 ),
    .i1(\u_EXU_LSU/n144 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [24]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u209  (
    .i0(\u_EXU_LSU/n159 ),
    .i1(\u_EXU_LSU/n143 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [25]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u210  (
    .i0(\u_EXU_LSU/n158 ),
    .i1(\u_EXU_LSU/n142 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [26]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u211  (
    .i0(\u_EXU_LSU/n157 ),
    .i1(\u_EXU_LSU/n102 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [27]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u212  (
    .i0(\u_EXU_LSU/n156 ),
    .i1(\u_EXU_LSU/n101 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [28]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u213  (
    .i0(\u_EXU_LSU/n155 ),
    .i1(\u_EXU_LSU/n100 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [29]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u214  (
    .i0(\u_EXU_LSU/n154 ),
    .i1(\u_EXU_LSU/n99 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [30]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u215  (
    .i0(\u_EXU_LSU/n153 ),
    .i1(\u_EXU_LSU/n98 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [31]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u216  (
    .i0(\u_EXU_LSU/n152 ),
    .i1(\u_EXU_LSU/n97 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [32]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u217  (
    .i0(\u_EXU_LSU/n151 ),
    .i1(\u_EXU_LSU/n48 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [33]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u218  (
    .i0(\u_EXU_LSU/n150 ),
    .i1(\u_EXU_LSU/n47 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [34]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u219  (
    .i0(\u_EXU_LSU/n149 ),
    .i1(\u_EXU_LSU/n46 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [35]));  // ../RTL/core/exu_lsu.v(209)
  and \u_EXU_LSU/u21_sel_is_2  (\u_EXU_LSU/u21_sel_is_2_o , \u_EXU_LSU/n13_neg , lsu_flush);
  not \u_EXU_LSU/u21_sel_is_2_o_inv  (\u_EXU_LSU/u21_sel_is_2_o_neg , \u_EXU_LSU/u21_sel_is_2_o );
  AL_MUX \u_EXU_LSU/u22  (
    .i0(1'b0),
    .i1(o_exu_rdwen2),
    .sel(\u_EXU_LSU/u22_sel_is_0_o ),
    .o(\u_EXU_LSU/n18 ));
  AL_MUX \u_EXU_LSU/u220  (
    .i0(\u_EXU_LSU/n148 ),
    .i1(\u_EXU_LSU/n45 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [36]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u221  (
    .i0(\u_EXU_LSU/n147 ),
    .i1(\u_EXU_LSU/n44 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [37]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u222  (
    .i0(\u_EXU_LSU/n146 ),
    .i1(\u_EXU_LSU/n43 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [38]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u223  (
    .i0(\u_EXU_LSU/n145 ),
    .i1(\u_EXU_LSU/n42 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [39]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u224  (
    .i0(\u_EXU_LSU/n144 ),
    .i1(\u_EXU_LSU/n174 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [40]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u225  (
    .i0(\u_EXU_LSU/n143 ),
    .i1(\u_EXU_LSU/n175 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [41]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u226  (
    .i0(\u_EXU_LSU/n142 ),
    .i1(\u_EXU_LSU/n176 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [42]));  // ../RTL/core/exu_lsu.v(209)
  AL_MUX \u_EXU_LSU/u227  (
    .i0(\u_EXU_LSU/n102 ),
    .i1(\u_EXU_LSU/n177 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [43]));  // ../RTL/core/exu_lsu.v(209)
  and \u_EXU_LSU/u22_sel_is_0  (\u_EXU_LSU/u22_sel_is_0_o , \u_EXU_LSU/lsu_finish_neg , \u_EXU_LSU/u21_sel_is_2_o_neg );
  AL_MUX \u_EXU_LSU/u23  (
    .i0(\u_EXU_LSU/working ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/lsu_finish ),
    .o(\u_EXU_LSU/n19 ));  // ../RTL/core/exu_lsu.v(129)
  AL_MUX \u_EXU_LSU/u24  (
    .i0(\u_EXU_LSU/access2_vld ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/lsu_finish ),
    .o(\u_EXU_LSU/n20 ));  // ../RTL/core/exu_lsu.v(129)
  AL_MUX \u_EXU_LSU/u252  (
    .i0(\u_EXU_LSU/rs2rdata_reg [0]),
    .i1(\u_EXU_LSU/rs2rdata_reg [8]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n182 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u253  (
    .i0(\u_EXU_LSU/rs2rdata_reg [1]),
    .i1(\u_EXU_LSU/rs2rdata_reg [9]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n183 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u254  (
    .i0(\u_EXU_LSU/rs2rdata_reg [2]),
    .i1(\u_EXU_LSU/rs2rdata_reg [10]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n184 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u255  (
    .i0(\u_EXU_LSU/rs2rdata_reg [3]),
    .i1(\u_EXU_LSU/rs2rdata_reg [11]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n185 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u256  (
    .i0(\u_EXU_LSU/rs2rdata_reg [4]),
    .i1(\u_EXU_LSU/rs2rdata_reg [12]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n186 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u257  (
    .i0(\u_EXU_LSU/rs2rdata_reg [5]),
    .i1(\u_EXU_LSU/rs2rdata_reg [13]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n187 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u258  (
    .i0(\u_EXU_LSU/rs2rdata_reg [6]),
    .i1(\u_EXU_LSU/rs2rdata_reg [14]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n188 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u259  (
    .i0(\u_EXU_LSU/rs2rdata_reg [7]),
    .i1(\u_EXU_LSU/rs2rdata_reg [15]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n189 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u26  (
    .i0(\u_EXU_LSU/n18 ),
    .i1(\u_EXU_LSU/n8 ),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n23 ));  // ../RTL/core/exu_lsu.v(111)
  AL_MUX \u_EXU_LSU/u260  (
    .i0(\u_EXU_LSU/rs2rdata_reg [8]),
    .i1(\u_EXU_LSU/rs2rdata_reg [16]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n190 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u261  (
    .i0(\u_EXU_LSU/rs2rdata_reg [9]),
    .i1(\u_EXU_LSU/rs2rdata_reg [17]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n191 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u262  (
    .i0(\u_EXU_LSU/rs2rdata_reg [10]),
    .i1(\u_EXU_LSU/rs2rdata_reg [18]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n192 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u263  (
    .i0(\u_EXU_LSU/rs2rdata_reg [11]),
    .i1(\u_EXU_LSU/rs2rdata_reg [19]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n193 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u264  (
    .i0(\u_EXU_LSU/rs2rdata_reg [12]),
    .i1(\u_EXU_LSU/rs2rdata_reg [20]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n194 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u265  (
    .i0(\u_EXU_LSU/rs2rdata_reg [13]),
    .i1(\u_EXU_LSU/rs2rdata_reg [21]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n195 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u266  (
    .i0(\u_EXU_LSU/rs2rdata_reg [14]),
    .i1(\u_EXU_LSU/rs2rdata_reg [22]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n196 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u267  (
    .i0(\u_EXU_LSU/rs2rdata_reg [15]),
    .i1(\u_EXU_LSU/rs2rdata_reg [23]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n197 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u268  (
    .i0(\u_EXU_LSU/rs2rdata_reg [16]),
    .i1(\u_EXU_LSU/rs2rdata_reg [24]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n198 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u269  (
    .i0(\u_EXU_LSU/rs2rdata_reg [17]),
    .i1(\u_EXU_LSU/rs2rdata_reg [25]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n199 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u27  (
    .i0(\u_EXU_LSU/n19 ),
    .i1(1'b1),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n25 ));  // ../RTL/core/exu_lsu.v(111)
  AL_MUX \u_EXU_LSU/u270  (
    .i0(\u_EXU_LSU/rs2rdata_reg [18]),
    .i1(\u_EXU_LSU/rs2rdata_reg [26]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n200 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u271  (
    .i0(\u_EXU_LSU/rs2rdata_reg [19]),
    .i1(\u_EXU_LSU/rs2rdata_reg [27]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n201 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u272  (
    .i0(\u_EXU_LSU/rs2rdata_reg [20]),
    .i1(\u_EXU_LSU/rs2rdata_reg [28]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n202 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u273  (
    .i0(\u_EXU_LSU/rs2rdata_reg [21]),
    .i1(\u_EXU_LSU/rs2rdata_reg [29]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n203 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u274  (
    .i0(\u_EXU_LSU/rs2rdata_reg [22]),
    .i1(\u_EXU_LSU/rs2rdata_reg [30]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n204 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u275  (
    .i0(\u_EXU_LSU/rs2rdata_reg [23]),
    .i1(\u_EXU_LSU/rs2rdata_reg [31]),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n205 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u276  (
    .i0(\u_EXU_LSU/rs2rdata_reg [24]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n206 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u277  (
    .i0(\u_EXU_LSU/rs2rdata_reg [25]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n207 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u278  (
    .i0(\u_EXU_LSU/rs2rdata_reg [26]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n208 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u279  (
    .i0(\u_EXU_LSU/rs2rdata_reg [27]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n209 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u28  (
    .i0(\u_EXU_LSU/n20 ),
    .i1(\u_EXU_LSU/n12 ),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n26 ));  // ../RTL/core/exu_lsu.v(111)
  AL_MUX \u_EXU_LSU/u280  (
    .i0(\u_EXU_LSU/rs2rdata_reg [28]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n210 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u281  (
    .i0(\u_EXU_LSU/rs2rdata_reg [29]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n211 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u282  (
    .i0(\u_EXU_LSU/rs2rdata_reg [30]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n212 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u283  (
    .i0(\u_EXU_LSU/rs2rdata_reg [31]),
    .i1(1'b0),
    .sel(\u_EXU_LSU/n66 [0]),
    .o(\u_EXU_LSU/n213 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u284  (
    .i0(\u_EXU_LSU/n182 ),
    .i1(\u_EXU_LSU/n198 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n214 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u285  (
    .i0(\u_EXU_LSU/n183 ),
    .i1(\u_EXU_LSU/n199 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n215 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u286  (
    .i0(\u_EXU_LSU/n184 ),
    .i1(\u_EXU_LSU/n200 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n216 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u287  (
    .i0(\u_EXU_LSU/n185 ),
    .i1(\u_EXU_LSU/n201 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n217 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u288  (
    .i0(\u_EXU_LSU/n186 ),
    .i1(\u_EXU_LSU/n202 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n218 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u289  (
    .i0(\u_EXU_LSU/n187 ),
    .i1(\u_EXU_LSU/n203 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n219 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u29  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n16 ),
    .sel(\u_EXU_LSU/u29_sel_is_0_o ),
    .o(\u_EXU_LSU/n30 ));
  AL_MUX \u_EXU_LSU/u290  (
    .i0(\u_EXU_LSU/n188 ),
    .i1(\u_EXU_LSU/n204 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n220 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u291  (
    .i0(\u_EXU_LSU/n189 ),
    .i1(\u_EXU_LSU/n205 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n221 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u292  (
    .i0(\u_EXU_LSU/n190 ),
    .i1(\u_EXU_LSU/n206 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n222 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u293  (
    .i0(\u_EXU_LSU/n191 ),
    .i1(\u_EXU_LSU/n207 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n223 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u294  (
    .i0(\u_EXU_LSU/n192 ),
    .i1(\u_EXU_LSU/n208 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n224 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u295  (
    .i0(\u_EXU_LSU/n193 ),
    .i1(\u_EXU_LSU/n209 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n225 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u296  (
    .i0(\u_EXU_LSU/n194 ),
    .i1(\u_EXU_LSU/n210 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n226 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u297  (
    .i0(\u_EXU_LSU/n195 ),
    .i1(\u_EXU_LSU/n211 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n227 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u298  (
    .i0(\u_EXU_LSU/n196 ),
    .i1(\u_EXU_LSU/n212 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n228 ));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u299  (
    .i0(\u_EXU_LSU/n197 ),
    .i1(\u_EXU_LSU/n213 ),
    .sel(\u_EXU_LSU/n66 [1]),
    .o(\u_EXU_LSU/n229 ));  // ../RTL/core/exu_lsu.v(194)
  and \u_EXU_LSU/u29_sel_is_0  (\u_EXU_LSU/u29_sel_is_0_o , \u_EXU_LSU/lsu_vld_neg , \u_EXU_LSU/lsu_finish_neg );
  and \u_EXU_LSU/u3  (\u_EXU_LSU/handshake_rdy , o_ribm_req, i_ribm_gnt);  // ../RTL/core/exu_lsu.v(66)
  and \u_EXU_LSU/u30  (\u_EXU_LSU/n37 , \u_EXU_LSU/trans_finish , \u_EXU_LSU/access2_once );  // ../RTL/core/exu_lsu.v(145)
  not \u_EXU_LSU/u31  (\u_EXU_LSU/n38 , \u_EXU_LSU/n37 );  // ../RTL/core/exu_lsu.v(145)
  and \u_EXU_LSU/u32  (\u_EXU_LSU/n39 , \u_EXU_LSU/working , \u_EXU_LSU/n38 );  // ../RTL/core/exu_lsu.v(145)
  AL_MUX \u_EXU_LSU/u320  (
    .i0(\u_EXU_LSU/n214 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [0]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u321  (
    .i0(\u_EXU_LSU/n215 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [1]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u322  (
    .i0(\u_EXU_LSU/n216 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [2]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u323  (
    .i0(\u_EXU_LSU/n217 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [3]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u324  (
    .i0(\u_EXU_LSU/n218 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [4]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u325  (
    .i0(\u_EXU_LSU/n219 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [5]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u326  (
    .i0(\u_EXU_LSU/n220 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [6]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u327  (
    .i0(\u_EXU_LSU/n221 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [7]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u328  (
    .i0(\u_EXU_LSU/n222 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [8]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u329  (
    .i0(\u_EXU_LSU/n223 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [9]));  // ../RTL/core/exu_lsu.v(194)
  not \u_EXU_LSU/u33  (\u_EXU_LSU/n40 , \u_EXU_LSU/trans_finish );  // ../RTL/core/exu_lsu.v(145)
  AL_MUX \u_EXU_LSU/u330  (
    .i0(\u_EXU_LSU/n224 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [10]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u331  (
    .i0(\u_EXU_LSU/n225 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [11]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u332  (
    .i0(\u_EXU_LSU/n226 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [12]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u333  (
    .i0(\u_EXU_LSU/n227 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [13]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u334  (
    .i0(\u_EXU_LSU/n228 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [14]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u335  (
    .i0(\u_EXU_LSU/n229 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/sub0_2_co_neg ),
    .o(\u_EXU_LSU/n67 [15]));  // ../RTL/core/exu_lsu.v(194)
  AL_MUX \u_EXU_LSU/u336  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n198 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [16]));
  and \u_EXU_LSU/u336_sel_is_0  (\u_EXU_LSU/u336_sel_is_0_o , \u_EXU_LSU/sub0_2_co , \u_EXU_LSU/n66[1]_neg );
  AL_MUX \u_EXU_LSU/u337  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n199 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [17]));
  AL_MUX \u_EXU_LSU/u338  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n200 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [18]));
  AL_MUX \u_EXU_LSU/u339  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n201 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [19]));
  and \u_EXU_LSU/u34  (\u_EXU_LSU/n41 , \u_EXU_LSU/working , \u_EXU_LSU/n40 );  // ../RTL/core/exu_lsu.v(145)
  AL_MUX \u_EXU_LSU/u340  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n202 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [20]));
  AL_MUX \u_EXU_LSU/u341  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n203 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [21]));
  AL_MUX \u_EXU_LSU/u342  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n204 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [22]));
  AL_MUX \u_EXU_LSU/u343  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n205 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [23]));
  AL_MUX \u_EXU_LSU/u344  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n206 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [24]));
  AL_MUX \u_EXU_LSU/u345  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n207 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [25]));
  AL_MUX \u_EXU_LSU/u346  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n208 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [26]));
  AL_MUX \u_EXU_LSU/u347  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n209 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [27]));
  AL_MUX \u_EXU_LSU/u348  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n210 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [28]));
  AL_MUX \u_EXU_LSU/u349  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n211 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [29]));
  AL_MUX \u_EXU_LSU/u35  (
    .i0(\u_EXU_LSU/n41 ),
    .i1(\u_EXU_LSU/n39 ),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(o_lsu_working));  // ../RTL/core/exu_lsu.v(145)
  AL_MUX \u_EXU_LSU/u350  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n212 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [30]));
  AL_MUX \u_EXU_LSU/u351  (
    .i0(1'b0),
    .i1(\u_EXU_LSU/n213 ),
    .sel(\u_EXU_LSU/u336_sel_is_0_o ),
    .o(\u_EXU_LSU/n67 [31]));
  not \u_EXU_LSU/u352  (\u_EXU_LSU/n63 [2], \u_EXU_LSU/n62 [2]);  // ../RTL/core/exu_lsu.v(191)
  not \u_EXU_LSU/u353  (\u_EXU_LSU/n63 [3], \u_EXU_LSU/align_mode_reg [1]);  // ../RTL/core/exu_lsu.v(191)
  not \u_EXU_LSU/u354  (\u_EXU_LSU/n250 , \u_EXU_LSU/align_mode_reg [0]);  // ../RTL/core/exu_lsu.v(191)
  AL_MUX \u_EXU_LSU/u355  (
    .i0(\u_EXU_LSU/align_mode_reg [0]),
    .i1(\u_EXU_LSU/n250 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/n62 [2]));  // ../RTL/core/exu_lsu.v(191)
  AL_MUX \u_EXU_LSU/u356  (
    .i0(\u_EXU_LSU/n250 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/n62 [0]));  // ../RTL/core/exu_lsu.v(191)
  not \u_EXU_LSU/u357  (\u_EXU_LSU/n61 [2], \u_EXU_LSU/n60 [2]);  // ../RTL/core/exu_lsu.v(190)
  AL_MUX \u_EXU_LSU/u359  (
    .i0(1'b1),
    .i1(\u_EXU_LSU/n250 ),
    .sel(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/n60 [2]));  // ../RTL/core/exu_lsu.v(190)
  AL_MUX \u_EXU_LSU/u361  (
    .i0(i_rs2rdata[31]),
    .i1(i_rs2rdata[23]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n252 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u362  (
    .i0(i_rs2rdata[30]),
    .i1(i_rs2rdata[22]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n253 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u363  (
    .i0(i_rs2rdata[29]),
    .i1(i_rs2rdata[21]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n254 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u364  (
    .i0(i_rs2rdata[28]),
    .i1(i_rs2rdata[20]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n255 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u365  (
    .i0(i_rs2rdata[27]),
    .i1(i_rs2rdata[19]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n256 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u366  (
    .i0(i_rs2rdata[26]),
    .i1(i_rs2rdata[18]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n257 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u367  (
    .i0(i_rs2rdata[25]),
    .i1(i_rs2rdata[17]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n258 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u368  (
    .i0(i_rs2rdata[24]),
    .i1(i_rs2rdata[16]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n259 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u369  (
    .i0(i_rs2rdata[23]),
    .i1(i_rs2rdata[15]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n260 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u370  (
    .i0(i_rs2rdata[22]),
    .i1(i_rs2rdata[14]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n261 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u371  (
    .i0(i_rs2rdata[21]),
    .i1(i_rs2rdata[13]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n262 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u372  (
    .i0(i_rs2rdata[20]),
    .i1(i_rs2rdata[12]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n263 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u373  (
    .i0(i_rs2rdata[19]),
    .i1(i_rs2rdata[11]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n264 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u374  (
    .i0(i_rs2rdata[18]),
    .i1(i_rs2rdata[10]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n265 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u375  (
    .i0(i_rs2rdata[17]),
    .i1(i_rs2rdata[9]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n266 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u376  (
    .i0(i_rs2rdata[16]),
    .i1(i_rs2rdata[8]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n267 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u377  (
    .i0(i_rs2rdata[15]),
    .i1(i_rs2rdata[7]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n268 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u378  (
    .i0(i_rs2rdata[14]),
    .i1(i_rs2rdata[6]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n269 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u379  (
    .i0(i_rs2rdata[13]),
    .i1(i_rs2rdata[5]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n270 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u380  (
    .i0(i_rs2rdata[12]),
    .i1(i_rs2rdata[4]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n271 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u381  (
    .i0(i_rs2rdata[11]),
    .i1(i_rs2rdata[3]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n272 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u382  (
    .i0(i_rs2rdata[10]),
    .i1(i_rs2rdata[2]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n273 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u383  (
    .i0(i_rs2rdata[9]),
    .i1(i_rs2rdata[1]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n274 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u384  (
    .i0(i_rs2rdata[8]),
    .i1(i_rs2rdata[0]),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n275 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u385  (
    .i0(i_rs2rdata[7]),
    .i1(1'b0),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n276 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u386  (
    .i0(i_rs2rdata[6]),
    .i1(1'b0),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n277 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u387  (
    .i0(i_rs2rdata[5]),
    .i1(1'b0),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n278 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u388  (
    .i0(i_rs2rdata[4]),
    .i1(1'b0),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n279 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u389  (
    .i0(i_rs2rdata[3]),
    .i1(1'b0),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n280 ));  // ../RTL/core/exu_lsu.v(174)
  and \u_EXU_LSU/u39  (\u_EXU_LSU/lsu_finish , \u_EXU_LSU/n5 , \u_EXU_LSU/trans_finish );  // ../RTL/core/exu_lsu.v(103)
  AL_MUX \u_EXU_LSU/u390  (
    .i0(i_rs2rdata[2]),
    .i1(1'b0),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n281 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u391  (
    .i0(i_rs2rdata[1]),
    .i1(1'b0),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n282 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u392  (
    .i0(i_rs2rdata[0]),
    .i1(1'b0),
    .sel(alu2lsu_result[0]),
    .o(\u_EXU_LSU/n283 ));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u393  (
    .i0(\u_EXU_LSU/n252 ),
    .i1(\u_EXU_LSU/n268 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [31]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u394  (
    .i0(\u_EXU_LSU/n253 ),
    .i1(\u_EXU_LSU/n269 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [30]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u395  (
    .i0(\u_EXU_LSU/n254 ),
    .i1(\u_EXU_LSU/n270 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [29]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u396  (
    .i0(\u_EXU_LSU/n255 ),
    .i1(\u_EXU_LSU/n271 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [28]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u397  (
    .i0(\u_EXU_LSU/n256 ),
    .i1(\u_EXU_LSU/n272 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [27]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u398  (
    .i0(\u_EXU_LSU/n257 ),
    .i1(\u_EXU_LSU/n273 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [26]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u399  (
    .i0(\u_EXU_LSU/n258 ),
    .i1(\u_EXU_LSU/n274 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [25]));  // ../RTL/core/exu_lsu.v(174)
  not \u_EXU_LSU/u40  (\u_EXU_LSU/n56 , \u_EXU_LSU/handshake_once );  // ../RTL/core/exu_lsu.v(179)
  AL_MUX \u_EXU_LSU/u400  (
    .i0(\u_EXU_LSU/n259 ),
    .i1(\u_EXU_LSU/n275 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [24]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u401  (
    .i0(\u_EXU_LSU/n260 ),
    .i1(\u_EXU_LSU/n276 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [23]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u402  (
    .i0(\u_EXU_LSU/n261 ),
    .i1(\u_EXU_LSU/n277 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [22]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u403  (
    .i0(\u_EXU_LSU/n262 ),
    .i1(\u_EXU_LSU/n278 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [21]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u404  (
    .i0(\u_EXU_LSU/n263 ),
    .i1(\u_EXU_LSU/n279 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [20]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u405  (
    .i0(\u_EXU_LSU/n264 ),
    .i1(\u_EXU_LSU/n280 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [19]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u406  (
    .i0(\u_EXU_LSU/n265 ),
    .i1(\u_EXU_LSU/n281 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [18]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u407  (
    .i0(\u_EXU_LSU/n266 ),
    .i1(\u_EXU_LSU/n282 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [17]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u408  (
    .i0(\u_EXU_LSU/n267 ),
    .i1(\u_EXU_LSU/n283 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [16]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u409  (
    .i0(\u_EXU_LSU/n268 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [15]));  // ../RTL/core/exu_lsu.v(174)
  and \u_EXU_LSU/u41  (\u_EXU_LSU/n57 , \u_EXU_LSU/n56 , \u_EXU_LSU/access2_vld );  // ../RTL/core/exu_lsu.v(179)
  AL_MUX \u_EXU_LSU/u410  (
    .i0(\u_EXU_LSU/n269 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [14]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u411  (
    .i0(\u_EXU_LSU/n270 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [13]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u412  (
    .i0(\u_EXU_LSU/n271 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [12]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u413  (
    .i0(\u_EXU_LSU/n272 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [11]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u414  (
    .i0(\u_EXU_LSU/n273 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [10]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u415  (
    .i0(\u_EXU_LSU/n274 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [9]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u416  (
    .i0(\u_EXU_LSU/n275 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [8]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u417  (
    .i0(\u_EXU_LSU/n276 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [7]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u418  (
    .i0(\u_EXU_LSU/n277 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [6]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u419  (
    .i0(\u_EXU_LSU/n278 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [5]));  // ../RTL/core/exu_lsu.v(174)
  and \u_EXU_LSU/u42  (\u_EXU_LSU/n58 , \u_EXU_LSU/n57 , \u_EXU_LSU/handshake_rdy );  // ../RTL/core/exu_lsu.v(179)
  AL_MUX \u_EXU_LSU/u420  (
    .i0(\u_EXU_LSU/n279 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [4]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u421  (
    .i0(\u_EXU_LSU/n280 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [3]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u422  (
    .i0(\u_EXU_LSU/n281 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [2]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u423  (
    .i0(\u_EXU_LSU/n282 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [1]));  // ../RTL/core/exu_lsu.v(174)
  AL_MUX \u_EXU_LSU/u424  (
    .i0(\u_EXU_LSU/n283 ),
    .i1(1'b0),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n55 [0]));  // ../RTL/core/exu_lsu.v(174)
  not \u_EXU_LSU/u425  (\u_EXU_LSU/n284 , alu2lsu_result[0]);  // ../RTL/core/exu_lsu.v(171)
  not \u_EXU_LSU/u43  (\u_EXU_LSU/n61 [0], \u_EXU_LSU/n62 [0]);  // ../RTL/core/exu_lsu.v(190)
  AL_MUX \u_EXU_LSU/u433  (
    .i0(alu2lsu_result[0]),
    .i1(\u_EXU_LSU/n284 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n50 [2]));  // ../RTL/core/exu_lsu.v(170)
  AL_MUX \u_EXU_LSU/u439  (
    .i0(1'b1),
    .i1(\u_EXU_LSU/n284 ),
    .sel(alu2lsu_result[1]),
    .o(\u_EXU_LSU/n49 [2]));  // ../RTL/core/exu_lsu.v(169)
  AL_MUX \u_EXU_LSU/u45  (
    .i0(o_ribm_req),
    .i1(1'b0),
    .sel(\u_EXU_LSU/handshake_rdy ),
    .o(\u_EXU_LSU/n68 ));  // ../RTL/core/exu_lsu.v(197)
  AL_MUX \u_EXU_LSU/u46  (
    .i0(\u_EXU_LSU/handshake_once ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/handshake_rdy ),
    .o(\u_EXU_LSU/n69 ));  // ../RTL/core/exu_lsu.v(197)
  AL_MUX \u_EXU_LSU/u47  (
    .i0(\u_EXU_LSU/n69 ),
    .i1(1'b1),
    .sel(\u_EXU_LSU/n58 ),
    .o(\u_EXU_LSU/n70 ));  // ../RTL/core/exu_lsu.v(179)
  AL_MUX \u_EXU_LSU/u49  (
    .i0(1'b1),
    .i1(\u_EXU_LSU/n68 ),
    .sel(\u_EXU_LSU/mux20_b0_sel_is_0_o ),
    .o(\u_EXU_LSU/n75 ));
  and \u_EXU_LSU/u5  (\u_EXU_LSU/trans_finish , \u_EXU_LSU/handshake_rdy_last , i_ribm_rsp);  // ../RTL/core/exu_lsu.v(71)
  AL_MUX \u_EXU_LSU/u51  (
    .i0(\u_EXU_LSU/n70 ),
    .i1(1'b0),
    .sel(\u_EXU_LSU/lsu_vld ),
    .o(\u_EXU_LSU/n80 ));  // ../RTL/core/exu_lsu.v(160)
  AL_MUX \u_EXU_LSU/u53  (
    .i0(o_exu_rdwen2),
    .i1(\u_EXU_LSU/access2_once ),
    .sel(\u_EXU_LSU/access2_vld ),
    .o(\u_EXU_LSU/n96 ));  // ../RTL/core/exu_lsu.v(206)
  and \u_EXU_LSU/u54  (o_rdwen2, \u_EXU_LSU/n96 , \u_EXU_LSU/trans_finish );  // ../RTL/core/exu_lsu.v(206)
  not \u_EXU_LSU/u7  (\u_EXU_LSU/n0 , \u_EXU_LSU/handshake_rdy_last );  // ../RTL/core/exu_lsu.v(78)
  or \u_EXU_LSU/u8  (\u_EXU_LSU/n1 , i_ribm_rsp, \u_EXU_LSU/n0 );  // ../RTL/core/exu_lsu.v(78)
  AL_DFF_X \u_EXU_LSU/working_reg  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_EXU_LSU/n25 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_EXU_LSU/working ));  // ../RTL/core/exu_lsu.v(105)
  EXU_MDU u_EXU_MDU (
    .i_clk(i_clk),
    .i_decinfo_grp(i_decinfo_grp),
    .i_flush(mdu_flush),
    .i_mdu_op1(i_exu_op1),
    .i_mdu_op2(i_exu_op2),
    .i_mdu_rdidx(o_rdidx0),
    .i_mdu_rdwen(o_exu_rdwen0),
    .i_mduinfo({i_decinfo[9:1],1'b0}),
    .i_rstn(i_rstn),
    .i_vld(i_vld),
    .o_mdu_rdidx(o_rdidx1),
    .o_mdu_rdwdata(o_rdwdata1),
    .o_mdu_rdwen(o_rdwen1),
    .o_will_rdidx(o_exu_rdidx1),
    .o_will_rdwen(o_exu_rdwen1),
    .o_working(o_mdu_working));  // ../RTL/core/exu.v(176)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b0  (
    .i0(i_exu_op1[0]),
    .i1(i_csr_zimm[0]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [0]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b1  (
    .i0(i_exu_op1[1]),
    .i1(i_csr_zimm[1]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [1]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b10  (
    .i0(i_exu_op1[10]),
    .i1(i_csr_zimm[10]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [10]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b11  (
    .i0(i_exu_op1[11]),
    .i1(i_csr_zimm[11]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [11]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b12  (
    .i0(i_exu_op1[12]),
    .i1(i_csr_zimm[12]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [12]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b13  (
    .i0(i_exu_op1[13]),
    .i1(i_csr_zimm[13]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [13]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b14  (
    .i0(i_exu_op1[14]),
    .i1(i_csr_zimm[14]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [14]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b15  (
    .i0(i_exu_op1[15]),
    .i1(i_csr_zimm[15]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [15]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b16  (
    .i0(i_exu_op1[16]),
    .i1(i_csr_zimm[16]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [16]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b17  (
    .i0(i_exu_op1[17]),
    .i1(i_csr_zimm[17]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [17]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b18  (
    .i0(i_exu_op1[18]),
    .i1(i_csr_zimm[18]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [18]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b19  (
    .i0(i_exu_op1[19]),
    .i1(i_csr_zimm[19]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [19]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b2  (
    .i0(i_exu_op1[2]),
    .i1(i_csr_zimm[2]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [2]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b20  (
    .i0(i_exu_op1[20]),
    .i1(i_csr_zimm[20]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [20]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b21  (
    .i0(i_exu_op1[21]),
    .i1(i_csr_zimm[21]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [21]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b22  (
    .i0(i_exu_op1[22]),
    .i1(i_csr_zimm[22]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [22]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b23  (
    .i0(i_exu_op1[23]),
    .i1(i_csr_zimm[23]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [23]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b24  (
    .i0(i_exu_op1[24]),
    .i1(i_csr_zimm[24]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [24]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b25  (
    .i0(i_exu_op1[25]),
    .i1(i_csr_zimm[25]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [25]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b26  (
    .i0(i_exu_op1[26]),
    .i1(i_csr_zimm[26]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [26]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b27  (
    .i0(i_exu_op1[27]),
    .i1(i_csr_zimm[27]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [27]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b28  (
    .i0(i_exu_op1[28]),
    .i1(i_csr_zimm[28]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [28]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b29  (
    .i0(i_exu_op1[29]),
    .i1(i_csr_zimm[29]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [29]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b3  (
    .i0(i_exu_op1[3]),
    .i1(i_csr_zimm[3]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [3]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b30  (
    .i0(i_exu_op1[30]),
    .i1(i_csr_zimm[30]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [30]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b31  (
    .i0(i_exu_op1[31]),
    .i1(i_csr_zimm[31]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [31]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b4  (
    .i0(i_exu_op1[4]),
    .i1(i_csr_zimm[4]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [4]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b5  (
    .i0(i_exu_op1[5]),
    .i1(i_csr_zimm[5]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [5]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b6  (
    .i0(i_exu_op1[6]),
    .i1(i_csr_zimm[6]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [6]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b7  (
    .i0(i_exu_op1[7]),
    .i1(i_csr_zimm[7]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [7]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b8  (
    .i0(i_exu_op1[8]),
    .i1(i_csr_zimm[8]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [8]));  // ../RTL/core/exu_scu.v(47)
  binary_mux_s1_w1 \u_EXU_SCU/mux0_b9  (
    .i0(i_exu_op1[9]),
    .i1(i_csr_zimm[9]),
    .sel(i_decinfo[6]),
    .o(\u_EXU_SCU/csr_rw [9]));  // ../RTL/core/exu_scu.v(47)
  and \u_EXU_SCU/u0  (\u_EXU_SCU/n2 [5], i_decinfo[4], \u_EXU_SCU/csr_rs [5]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u1  (\u_EXU_SCU/n2 [4], i_decinfo[4], \u_EXU_SCU/csr_rs [4]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u10  (\u_EXU_SCU/n2 [7], i_decinfo[4], \u_EXU_SCU/csr_rs [7]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u104  (o_csr_wdata[1], \u_EXU_SCU/n3 [1], \u_EXU_SCU/n4 [1]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u105  (o_csr_wdata[2], \u_EXU_SCU/n3 [2], \u_EXU_SCU/n4 [2]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u106  (o_csr_wdata[3], \u_EXU_SCU/n3 [3], \u_EXU_SCU/n4 [3]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u107  (o_csr_wdata[4], \u_EXU_SCU/n3 [4], \u_EXU_SCU/n4 [4]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u108  (o_csr_wdata[5], \u_EXU_SCU/n3 [5], \u_EXU_SCU/n4 [5]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u109  (o_csr_wdata[6], \u_EXU_SCU/n3 [6], \u_EXU_SCU/n4 [6]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u11  (\u_EXU_SCU/csr_rc [0], i_csr_rdata[0], \u_EXU_SCU/n0 [0]);  // ../RTL/core/exu_scu.v(49)
  or \u_EXU_SCU/u110  (o_csr_wdata[7], \u_EXU_SCU/n3 [7], \u_EXU_SCU/n4 [7]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u111  (o_csr_wdata[8], \u_EXU_SCU/n3 [8], \u_EXU_SCU/n4 [8]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u112  (o_csr_wdata[9], \u_EXU_SCU/n3 [9], \u_EXU_SCU/n4 [9]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u113  (o_csr_wdata[10], \u_EXU_SCU/n3 [10], \u_EXU_SCU/n4 [10]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u114  (o_csr_wdata[11], \u_EXU_SCU/n3 [11], \u_EXU_SCU/n4 [11]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u115  (o_csr_wdata[12], \u_EXU_SCU/n3 [12], \u_EXU_SCU/n4 [12]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u116  (o_csr_wdata[13], \u_EXU_SCU/n3 [13], \u_EXU_SCU/n4 [13]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u117  (o_csr_wdata[14], \u_EXU_SCU/n3 [14], \u_EXU_SCU/n4 [14]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u118  (o_csr_wdata[15], \u_EXU_SCU/n3 [15], \u_EXU_SCU/n4 [15]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u119  (o_csr_wdata[16], \u_EXU_SCU/n3 [16], \u_EXU_SCU/n4 [16]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u12  (\u_EXU_SCU/n3 [0], \u_EXU_SCU/n1 [0], \u_EXU_SCU/n2 [0]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u120  (o_csr_wdata[17], \u_EXU_SCU/n3 [17], \u_EXU_SCU/n4 [17]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u121  (o_csr_wdata[18], \u_EXU_SCU/n3 [18], \u_EXU_SCU/n4 [18]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u122  (o_csr_wdata[19], \u_EXU_SCU/n3 [19], \u_EXU_SCU/n4 [19]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u123  (o_csr_wdata[20], \u_EXU_SCU/n3 [20], \u_EXU_SCU/n4 [20]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u124  (o_csr_wdata[21], \u_EXU_SCU/n3 [21], \u_EXU_SCU/n4 [21]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u125  (o_csr_wdata[22], \u_EXU_SCU/n3 [22], \u_EXU_SCU/n4 [22]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u126  (o_csr_wdata[23], \u_EXU_SCU/n3 [23], \u_EXU_SCU/n4 [23]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u127  (o_csr_wdata[24], \u_EXU_SCU/n3 [24], \u_EXU_SCU/n4 [24]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u128  (o_csr_wdata[25], \u_EXU_SCU/n3 [25], \u_EXU_SCU/n4 [25]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u129  (o_csr_wdata[26], \u_EXU_SCU/n3 [26], \u_EXU_SCU/n4 [26]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u13  (\u_EXU_SCU/n4 [0], i_decinfo[5], \u_EXU_SCU/csr_rc [0]);  // ../RTL/core/exu_scu.v(57)
  or \u_EXU_SCU/u130  (o_csr_wdata[27], \u_EXU_SCU/n3 [27], \u_EXU_SCU/n4 [27]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u131  (o_csr_wdata[28], \u_EXU_SCU/n3 [28], \u_EXU_SCU/n4 [28]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u132  (o_csr_wdata[29], \u_EXU_SCU/n3 [29], \u_EXU_SCU/n4 [29]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u133  (o_csr_wdata[30], \u_EXU_SCU/n3 [30], \u_EXU_SCU/n4 [30]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u134  (o_csr_wdata[31], \u_EXU_SCU/n3 [31], \u_EXU_SCU/n4 [31]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u135  (\u_EXU_SCU/n4 [1], i_decinfo[5], \u_EXU_SCU/csr_rc [1]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u136  (\u_EXU_SCU/n4 [2], i_decinfo[5], \u_EXU_SCU/csr_rc [2]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u137  (\u_EXU_SCU/n4 [3], i_decinfo[5], \u_EXU_SCU/csr_rc [3]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u138  (\u_EXU_SCU/n4 [4], i_decinfo[5], \u_EXU_SCU/csr_rc [4]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u139  (\u_EXU_SCU/n4 [5], i_decinfo[5], \u_EXU_SCU/csr_rc [5]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u140  (\u_EXU_SCU/n4 [6], i_decinfo[5], \u_EXU_SCU/csr_rc [6]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u141  (\u_EXU_SCU/n4 [7], i_decinfo[5], \u_EXU_SCU/csr_rc [7]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u142  (\u_EXU_SCU/n4 [8], i_decinfo[5], \u_EXU_SCU/csr_rc [8]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u143  (\u_EXU_SCU/n4 [9], i_decinfo[5], \u_EXU_SCU/csr_rc [9]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u144  (\u_EXU_SCU/n4 [10], i_decinfo[5], \u_EXU_SCU/csr_rc [10]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u145  (\u_EXU_SCU/n4 [11], i_decinfo[5], \u_EXU_SCU/csr_rc [11]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u146  (\u_EXU_SCU/n4 [12], i_decinfo[5], \u_EXU_SCU/csr_rc [12]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u147  (\u_EXU_SCU/n4 [13], i_decinfo[5], \u_EXU_SCU/csr_rc [13]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u148  (\u_EXU_SCU/n4 [14], i_decinfo[5], \u_EXU_SCU/csr_rc [14]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u149  (\u_EXU_SCU/n4 [15], i_decinfo[5], \u_EXU_SCU/csr_rc [15]);  // ../RTL/core/exu_scu.v(57)
  or \u_EXU_SCU/u15  (o_csr_wdata[0], \u_EXU_SCU/n3 [0], \u_EXU_SCU/n4 [0]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u150  (\u_EXU_SCU/n4 [16], i_decinfo[5], \u_EXU_SCU/csr_rc [16]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u151  (\u_EXU_SCU/n4 [17], i_decinfo[5], \u_EXU_SCU/csr_rc [17]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u152  (\u_EXU_SCU/n4 [18], i_decinfo[5], \u_EXU_SCU/csr_rc [18]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u153  (\u_EXU_SCU/n4 [19], i_decinfo[5], \u_EXU_SCU/csr_rc [19]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u154  (\u_EXU_SCU/n4 [20], i_decinfo[5], \u_EXU_SCU/csr_rc [20]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u155  (\u_EXU_SCU/n4 [21], i_decinfo[5], \u_EXU_SCU/csr_rc [21]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u156  (\u_EXU_SCU/n4 [22], i_decinfo[5], \u_EXU_SCU/csr_rc [22]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u157  (\u_EXU_SCU/n4 [23], i_decinfo[5], \u_EXU_SCU/csr_rc [23]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u158  (\u_EXU_SCU/n4 [24], i_decinfo[5], \u_EXU_SCU/csr_rc [24]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u159  (\u_EXU_SCU/n4 [25], i_decinfo[5], \u_EXU_SCU/csr_rc [25]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u160  (\u_EXU_SCU/n4 [26], i_decinfo[5], \u_EXU_SCU/csr_rc [26]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u161  (\u_EXU_SCU/n4 [27], i_decinfo[5], \u_EXU_SCU/csr_rc [27]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u162  (\u_EXU_SCU/n4 [28], i_decinfo[5], \u_EXU_SCU/csr_rc [28]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u163  (\u_EXU_SCU/n4 [29], i_decinfo[5], \u_EXU_SCU/csr_rc [29]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u164  (\u_EXU_SCU/n4 [30], i_decinfo[5], \u_EXU_SCU/csr_rc [30]);  // ../RTL/core/exu_scu.v(57)
  and \u_EXU_SCU/u165  (\u_EXU_SCU/n4 [31], i_decinfo[5], \u_EXU_SCU/csr_rc [31]);  // ../RTL/core/exu_scu.v(57)
  or \u_EXU_SCU/u166  (\u_EXU_SCU/n3 [1], \u_EXU_SCU/n1 [1], \u_EXU_SCU/n2 [1]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u167  (\u_EXU_SCU/n3 [2], \u_EXU_SCU/n1 [2], \u_EXU_SCU/n2 [2]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u168  (\u_EXU_SCU/n3 [3], \u_EXU_SCU/n1 [3], \u_EXU_SCU/n2 [3]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u169  (\u_EXU_SCU/n3 [4], \u_EXU_SCU/n1 [4], \u_EXU_SCU/n2 [4]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u17  (\u_EXU_SCU/n2 [8], i_decinfo[4], \u_EXU_SCU/csr_rs [8]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u170  (\u_EXU_SCU/n3 [5], \u_EXU_SCU/n1 [5], \u_EXU_SCU/n2 [5]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u171  (\u_EXU_SCU/n3 [6], \u_EXU_SCU/n1 [6], \u_EXU_SCU/n2 [6]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u172  (\u_EXU_SCU/n3 [7], \u_EXU_SCU/n1 [7], \u_EXU_SCU/n2 [7]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u173  (\u_EXU_SCU/n3 [8], \u_EXU_SCU/n1 [8], \u_EXU_SCU/n2 [8]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u174  (\u_EXU_SCU/n3 [9], \u_EXU_SCU/n1 [9], \u_EXU_SCU/n2 [9]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u175  (\u_EXU_SCU/n3 [10], \u_EXU_SCU/n1 [10], \u_EXU_SCU/n2 [10]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u176  (\u_EXU_SCU/n3 [11], \u_EXU_SCU/n1 [11], \u_EXU_SCU/n2 [11]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u177  (\u_EXU_SCU/n3 [12], \u_EXU_SCU/n1 [12], \u_EXU_SCU/n2 [12]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u178  (\u_EXU_SCU/n3 [13], \u_EXU_SCU/n1 [13], \u_EXU_SCU/n2 [13]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u179  (\u_EXU_SCU/n3 [14], \u_EXU_SCU/n1 [14], \u_EXU_SCU/n2 [14]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u18  (\u_EXU_SCU/n2 [9], i_decinfo[4], \u_EXU_SCU/csr_rs [9]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u180  (\u_EXU_SCU/n3 [15], \u_EXU_SCU/n1 [15], \u_EXU_SCU/n2 [15]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u181  (\u_EXU_SCU/n3 [16], \u_EXU_SCU/n1 [16], \u_EXU_SCU/n2 [16]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u182  (\u_EXU_SCU/n3 [17], \u_EXU_SCU/n1 [17], \u_EXU_SCU/n2 [17]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u183  (\u_EXU_SCU/n3 [18], \u_EXU_SCU/n1 [18], \u_EXU_SCU/n2 [18]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u184  (\u_EXU_SCU/n3 [19], \u_EXU_SCU/n1 [19], \u_EXU_SCU/n2 [19]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u185  (\u_EXU_SCU/n3 [20], \u_EXU_SCU/n1 [20], \u_EXU_SCU/n2 [20]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u186  (\u_EXU_SCU/n3 [21], \u_EXU_SCU/n1 [21], \u_EXU_SCU/n2 [21]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u187  (\u_EXU_SCU/n3 [22], \u_EXU_SCU/n1 [22], \u_EXU_SCU/n2 [22]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u188  (\u_EXU_SCU/n3 [23], \u_EXU_SCU/n1 [23], \u_EXU_SCU/n2 [23]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u189  (\u_EXU_SCU/n3 [24], \u_EXU_SCU/n1 [24], \u_EXU_SCU/n2 [24]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u19  (\u_EXU_SCU/n2 [10], i_decinfo[4], \u_EXU_SCU/csr_rs [10]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u190  (\u_EXU_SCU/n3 [25], \u_EXU_SCU/n1 [25], \u_EXU_SCU/n2 [25]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u191  (\u_EXU_SCU/n3 [26], \u_EXU_SCU/n1 [26], \u_EXU_SCU/n2 [26]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u192  (\u_EXU_SCU/n3 [27], \u_EXU_SCU/n1 [27], \u_EXU_SCU/n2 [27]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u193  (\u_EXU_SCU/n3 [28], \u_EXU_SCU/n1 [28], \u_EXU_SCU/n2 [28]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u194  (\u_EXU_SCU/n3 [29], \u_EXU_SCU/n1 [29], \u_EXU_SCU/n2 [29]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u195  (\u_EXU_SCU/n3 [30], \u_EXU_SCU/n1 [30], \u_EXU_SCU/n2 [30]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u196  (\u_EXU_SCU/n3 [31], \u_EXU_SCU/n1 [31], \u_EXU_SCU/n2 [31]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u197  (\u_EXU_SCU/csr_rc [1], i_csr_rdata[1], \u_EXU_SCU/n0 [1]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u198  (\u_EXU_SCU/csr_rc [2], i_csr_rdata[2], \u_EXU_SCU/n0 [2]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u199  (\u_EXU_SCU/csr_rc [3], i_csr_rdata[3], \u_EXU_SCU/n0 [3]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u2  (\u_EXU_SCU/n2 [3], i_decinfo[4], \u_EXU_SCU/csr_rs [3]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u20  (\u_EXU_SCU/n2 [11], i_decinfo[4], \u_EXU_SCU/csr_rs [11]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u200  (\u_EXU_SCU/csr_rc [4], i_csr_rdata[4], \u_EXU_SCU/n0 [4]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u201  (\u_EXU_SCU/csr_rc [5], i_csr_rdata[5], \u_EXU_SCU/n0 [5]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u202  (\u_EXU_SCU/csr_rc [6], i_csr_rdata[6], \u_EXU_SCU/n0 [6]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u203  (\u_EXU_SCU/csr_rc [7], i_csr_rdata[7], \u_EXU_SCU/n0 [7]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u204  (\u_EXU_SCU/csr_rc [8], i_csr_rdata[8], \u_EXU_SCU/n0 [8]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u205  (\u_EXU_SCU/csr_rc [9], i_csr_rdata[9], \u_EXU_SCU/n0 [9]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u206  (\u_EXU_SCU/csr_rc [10], i_csr_rdata[10], \u_EXU_SCU/n0 [10]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u207  (\u_EXU_SCU/csr_rc [11], i_csr_rdata[11], \u_EXU_SCU/n0 [11]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u208  (\u_EXU_SCU/csr_rc [12], i_csr_rdata[12], \u_EXU_SCU/n0 [12]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u209  (\u_EXU_SCU/csr_rc [13], i_csr_rdata[13], \u_EXU_SCU/n0 [13]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u21  (\u_EXU_SCU/n2 [12], i_decinfo[4], \u_EXU_SCU/csr_rs [12]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u210  (\u_EXU_SCU/csr_rc [14], i_csr_rdata[14], \u_EXU_SCU/n0 [14]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u211  (\u_EXU_SCU/csr_rc [15], i_csr_rdata[15], \u_EXU_SCU/n0 [15]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u212  (\u_EXU_SCU/csr_rc [16], i_csr_rdata[16], \u_EXU_SCU/n0 [16]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u213  (\u_EXU_SCU/csr_rc [17], i_csr_rdata[17], \u_EXU_SCU/n0 [17]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u214  (\u_EXU_SCU/csr_rc [18], i_csr_rdata[18], \u_EXU_SCU/n0 [18]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u215  (\u_EXU_SCU/csr_rc [19], i_csr_rdata[19], \u_EXU_SCU/n0 [19]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u216  (\u_EXU_SCU/csr_rc [20], i_csr_rdata[20], \u_EXU_SCU/n0 [20]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u217  (\u_EXU_SCU/csr_rc [21], i_csr_rdata[21], \u_EXU_SCU/n0 [21]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u218  (\u_EXU_SCU/csr_rc [22], i_csr_rdata[22], \u_EXU_SCU/n0 [22]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u219  (\u_EXU_SCU/csr_rc [23], i_csr_rdata[23], \u_EXU_SCU/n0 [23]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u22  (\u_EXU_SCU/n2 [13], i_decinfo[4], \u_EXU_SCU/csr_rs [13]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u220  (\u_EXU_SCU/csr_rc [24], i_csr_rdata[24], \u_EXU_SCU/n0 [24]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u221  (\u_EXU_SCU/csr_rc [25], i_csr_rdata[25], \u_EXU_SCU/n0 [25]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u222  (\u_EXU_SCU/csr_rc [26], i_csr_rdata[26], \u_EXU_SCU/n0 [26]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u223  (\u_EXU_SCU/csr_rc [27], i_csr_rdata[27], \u_EXU_SCU/n0 [27]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u224  (\u_EXU_SCU/csr_rc [28], i_csr_rdata[28], \u_EXU_SCU/n0 [28]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u225  (\u_EXU_SCU/csr_rc [29], i_csr_rdata[29], \u_EXU_SCU/n0 [29]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u226  (\u_EXU_SCU/csr_rc [30], i_csr_rdata[30], \u_EXU_SCU/n0 [30]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u227  (\u_EXU_SCU/csr_rc [31], i_csr_rdata[31], \u_EXU_SCU/n0 [31]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u228  (\u_EXU_SCU/n0 [1], \u_EXU_SCU/csr_rw [1]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u229  (\u_EXU_SCU/n0 [2], \u_EXU_SCU/csr_rw [2]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u23  (\u_EXU_SCU/n2 [14], i_decinfo[4], \u_EXU_SCU/csr_rs [14]);  // ../RTL/core/exu_scu.v(55)
  not \u_EXU_SCU/u230  (\u_EXU_SCU/n0 [3], \u_EXU_SCU/csr_rw [3]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u231  (\u_EXU_SCU/n0 [4], \u_EXU_SCU/csr_rw [4]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u232  (\u_EXU_SCU/n0 [5], \u_EXU_SCU/csr_rw [5]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u233  (\u_EXU_SCU/n0 [6], \u_EXU_SCU/csr_rw [6]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u234  (\u_EXU_SCU/n0 [7], \u_EXU_SCU/csr_rw [7]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u235  (\u_EXU_SCU/n0 [8], \u_EXU_SCU/csr_rw [8]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u236  (\u_EXU_SCU/n0 [9], \u_EXU_SCU/csr_rw [9]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u237  (\u_EXU_SCU/n0 [10], \u_EXU_SCU/csr_rw [10]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u238  (\u_EXU_SCU/n0 [11], \u_EXU_SCU/csr_rw [11]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u239  (\u_EXU_SCU/n0 [12], \u_EXU_SCU/csr_rw [12]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u24  (\u_EXU_SCU/n2 [15], i_decinfo[4], \u_EXU_SCU/csr_rs [15]);  // ../RTL/core/exu_scu.v(55)
  not \u_EXU_SCU/u240  (\u_EXU_SCU/n0 [13], \u_EXU_SCU/csr_rw [13]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u241  (\u_EXU_SCU/n0 [14], \u_EXU_SCU/csr_rw [14]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u242  (\u_EXU_SCU/n0 [15], \u_EXU_SCU/csr_rw [15]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u243  (\u_EXU_SCU/n0 [16], \u_EXU_SCU/csr_rw [16]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u244  (\u_EXU_SCU/n0 [17], \u_EXU_SCU/csr_rw [17]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u245  (\u_EXU_SCU/n0 [18], \u_EXU_SCU/csr_rw [18]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u246  (\u_EXU_SCU/n0 [19], \u_EXU_SCU/csr_rw [19]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u247  (\u_EXU_SCU/n0 [20], \u_EXU_SCU/csr_rw [20]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u248  (\u_EXU_SCU/n0 [21], \u_EXU_SCU/csr_rw [21]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u249  (\u_EXU_SCU/n0 [22], \u_EXU_SCU/csr_rw [22]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u25  (\u_EXU_SCU/n2 [16], i_decinfo[4], \u_EXU_SCU/csr_rs [16]);  // ../RTL/core/exu_scu.v(55)
  not \u_EXU_SCU/u250  (\u_EXU_SCU/n0 [23], \u_EXU_SCU/csr_rw [23]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u251  (\u_EXU_SCU/n0 [24], \u_EXU_SCU/csr_rw [24]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u252  (\u_EXU_SCU/n0 [25], \u_EXU_SCU/csr_rw [25]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u253  (\u_EXU_SCU/n0 [26], \u_EXU_SCU/csr_rw [26]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u254  (\u_EXU_SCU/n0 [27], \u_EXU_SCU/csr_rw [27]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u255  (\u_EXU_SCU/n0 [28], \u_EXU_SCU/csr_rw [28]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u256  (\u_EXU_SCU/n0 [29], \u_EXU_SCU/csr_rw [29]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u257  (\u_EXU_SCU/n0 [30], \u_EXU_SCU/csr_rw [30]);  // ../RTL/core/exu_scu.v(49)
  not \u_EXU_SCU/u258  (\u_EXU_SCU/n0 [31], \u_EXU_SCU/csr_rw [31]);  // ../RTL/core/exu_scu.v(49)
  or \u_EXU_SCU/u259  (\u_EXU_SCU/csr_rs [1], i_csr_rdata[1], \u_EXU_SCU/csr_rw [1]);  // ../RTL/core/exu_scu.v(48)
  and \u_EXU_SCU/u26  (\u_EXU_SCU/n2 [17], i_decinfo[4], \u_EXU_SCU/csr_rs [17]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u260  (\u_EXU_SCU/csr_rs [2], i_csr_rdata[2], \u_EXU_SCU/csr_rw [2]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u261  (\u_EXU_SCU/csr_rs [3], i_csr_rdata[3], \u_EXU_SCU/csr_rw [3]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u262  (\u_EXU_SCU/csr_rs [4], i_csr_rdata[4], \u_EXU_SCU/csr_rw [4]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u263  (\u_EXU_SCU/csr_rs [5], i_csr_rdata[5], \u_EXU_SCU/csr_rw [5]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u264  (\u_EXU_SCU/csr_rs [6], i_csr_rdata[6], \u_EXU_SCU/csr_rw [6]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u265  (\u_EXU_SCU/csr_rs [7], i_csr_rdata[7], \u_EXU_SCU/csr_rw [7]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u266  (\u_EXU_SCU/csr_rs [8], i_csr_rdata[8], \u_EXU_SCU/csr_rw [8]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u267  (\u_EXU_SCU/csr_rs [9], i_csr_rdata[9], \u_EXU_SCU/csr_rw [9]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u268  (\u_EXU_SCU/csr_rs [10], i_csr_rdata[10], \u_EXU_SCU/csr_rw [10]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u269  (\u_EXU_SCU/csr_rs [11], i_csr_rdata[11], \u_EXU_SCU/csr_rw [11]);  // ../RTL/core/exu_scu.v(48)
  and \u_EXU_SCU/u27  (\u_EXU_SCU/n2 [18], i_decinfo[4], \u_EXU_SCU/csr_rs [18]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u270  (\u_EXU_SCU/csr_rs [12], i_csr_rdata[12], \u_EXU_SCU/csr_rw [12]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u271  (\u_EXU_SCU/csr_rs [13], i_csr_rdata[13], \u_EXU_SCU/csr_rw [13]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u272  (\u_EXU_SCU/csr_rs [14], i_csr_rdata[14], \u_EXU_SCU/csr_rw [14]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u273  (\u_EXU_SCU/csr_rs [15], i_csr_rdata[15], \u_EXU_SCU/csr_rw [15]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u274  (\u_EXU_SCU/csr_rs [16], i_csr_rdata[16], \u_EXU_SCU/csr_rw [16]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u275  (\u_EXU_SCU/csr_rs [17], i_csr_rdata[17], \u_EXU_SCU/csr_rw [17]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u276  (\u_EXU_SCU/csr_rs [18], i_csr_rdata[18], \u_EXU_SCU/csr_rw [18]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u277  (\u_EXU_SCU/csr_rs [19], i_csr_rdata[19], \u_EXU_SCU/csr_rw [19]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u278  (\u_EXU_SCU/csr_rs [20], i_csr_rdata[20], \u_EXU_SCU/csr_rw [20]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u279  (\u_EXU_SCU/csr_rs [21], i_csr_rdata[21], \u_EXU_SCU/csr_rw [21]);  // ../RTL/core/exu_scu.v(48)
  and \u_EXU_SCU/u28  (\u_EXU_SCU/n2 [19], i_decinfo[4], \u_EXU_SCU/csr_rs [19]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u280  (\u_EXU_SCU/csr_rs [22], i_csr_rdata[22], \u_EXU_SCU/csr_rw [22]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u281  (\u_EXU_SCU/csr_rs [23], i_csr_rdata[23], \u_EXU_SCU/csr_rw [23]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u282  (\u_EXU_SCU/csr_rs [24], i_csr_rdata[24], \u_EXU_SCU/csr_rw [24]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u283  (\u_EXU_SCU/csr_rs [25], i_csr_rdata[25], \u_EXU_SCU/csr_rw [25]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u284  (\u_EXU_SCU/csr_rs [26], i_csr_rdata[26], \u_EXU_SCU/csr_rw [26]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u285  (\u_EXU_SCU/csr_rs [27], i_csr_rdata[27], \u_EXU_SCU/csr_rw [27]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u286  (\u_EXU_SCU/csr_rs [28], i_csr_rdata[28], \u_EXU_SCU/csr_rw [28]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u287  (\u_EXU_SCU/csr_rs [29], i_csr_rdata[29], \u_EXU_SCU/csr_rw [29]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u288  (\u_EXU_SCU/csr_rs [30], i_csr_rdata[30], \u_EXU_SCU/csr_rw [30]);  // ../RTL/core/exu_scu.v(48)
  or \u_EXU_SCU/u289  (\u_EXU_SCU/csr_rs [31], i_csr_rdata[31], \u_EXU_SCU/csr_rw [31]);  // ../RTL/core/exu_scu.v(48)
  and \u_EXU_SCU/u29  (\u_EXU_SCU/n2 [20], i_decinfo[4], \u_EXU_SCU/csr_rs [20]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u3  (\u_EXU_SCU/n2 [2], i_decinfo[4], \u_EXU_SCU/csr_rs [2]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u30  (\u_EXU_SCU/n2 [21], i_decinfo[4], \u_EXU_SCU/csr_rs [21]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u31  (\u_EXU_SCU/n2 [22], i_decinfo[4], \u_EXU_SCU/csr_rs [22]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u32  (\u_EXU_SCU/n2 [23], i_decinfo[4], \u_EXU_SCU/csr_rs [23]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u33  (\u_EXU_SCU/n2 [24], i_decinfo[4], \u_EXU_SCU/csr_rs [24]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u34  (\u_EXU_SCU/n2 [25], i_decinfo[4], \u_EXU_SCU/csr_rs [25]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u35  (\u_EXU_SCU/n2 [26], i_decinfo[4], \u_EXU_SCU/csr_rs [26]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u36  (\u_EXU_SCU/n2 [27], i_decinfo[4], \u_EXU_SCU/csr_rs [27]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u37  (\u_EXU_SCU/n2 [28], i_decinfo[4], \u_EXU_SCU/csr_rs [28]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u38  (\u_EXU_SCU/n2 [29], i_decinfo[4], \u_EXU_SCU/csr_rs [29]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u39  (\u_EXU_SCU/n2 [30], i_decinfo[4], \u_EXU_SCU/csr_rs [30]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u4  (\u_EXU_SCU/n2 [1], i_decinfo[4], \u_EXU_SCU/csr_rs [1]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u40  (\u_EXU_SCU/n2 [31], i_decinfo[4], \u_EXU_SCU/csr_rs [31]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u41  (\u_EXU_SCU/n1 [0], i_decinfo[3], \u_EXU_SCU/csr_rw [0]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u42  (\u_EXU_SCU/n1 [1], i_decinfo[3], \u_EXU_SCU/csr_rw [1]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u43  (\u_EXU_SCU/n1 [2], i_decinfo[3], \u_EXU_SCU/csr_rw [2]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u44  (\u_EXU_SCU/n1 [3], i_decinfo[3], \u_EXU_SCU/csr_rw [3]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u45  (\u_EXU_SCU/n1 [4], i_decinfo[3], \u_EXU_SCU/csr_rw [4]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u46  (\u_EXU_SCU/n1 [5], i_decinfo[3], \u_EXU_SCU/csr_rw [5]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u47  (\u_EXU_SCU/n1 [6], i_decinfo[3], \u_EXU_SCU/csr_rw [6]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u48  (\u_EXU_SCU/n1 [7], i_decinfo[3], \u_EXU_SCU/csr_rw [7]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u49  (\u_EXU_SCU/n1 [8], i_decinfo[3], \u_EXU_SCU/csr_rw [8]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u5  (\u_EXU_SCU/n2 [0], i_decinfo[4], \u_EXU_SCU/csr_rs [0]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u50  (\u_EXU_SCU/n1 [9], i_decinfo[3], \u_EXU_SCU/csr_rw [9]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u51  (\u_EXU_SCU/n1 [10], i_decinfo[3], \u_EXU_SCU/csr_rw [10]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u52  (\u_EXU_SCU/n1 [11], i_decinfo[3], \u_EXU_SCU/csr_rw [11]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u53  (\u_EXU_SCU/n1 [12], i_decinfo[3], \u_EXU_SCU/csr_rw [12]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u54  (\u_EXU_SCU/n1 [13], i_decinfo[3], \u_EXU_SCU/csr_rw [13]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u55  (\u_EXU_SCU/n1 [14], i_decinfo[3], \u_EXU_SCU/csr_rw [14]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u56  (\u_EXU_SCU/n1 [15], i_decinfo[3], \u_EXU_SCU/csr_rw [15]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u57  (\u_EXU_SCU/n1 [16], i_decinfo[3], \u_EXU_SCU/csr_rw [16]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u58  (\u_EXU_SCU/n1 [17], i_decinfo[3], \u_EXU_SCU/csr_rw [17]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u59  (\u_EXU_SCU/n1 [18], i_decinfo[3], \u_EXU_SCU/csr_rw [18]);  // ../RTL/core/exu_scu.v(55)
  or \u_EXU_SCU/u6  (\u_EXU_SCU/csr_rs [0], i_csr_rdata[0], \u_EXU_SCU/csr_rw [0]);  // ../RTL/core/exu_scu.v(48)
  and \u_EXU_SCU/u60  (\u_EXU_SCU/n1 [19], i_decinfo[3], \u_EXU_SCU/csr_rw [19]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u61  (\u_EXU_SCU/n1 [20], i_decinfo[3], \u_EXU_SCU/csr_rw [20]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u62  (\u_EXU_SCU/n1 [21], i_decinfo[3], \u_EXU_SCU/csr_rw [21]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u63  (\u_EXU_SCU/n1 [22], i_decinfo[3], \u_EXU_SCU/csr_rw [22]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u64  (\u_EXU_SCU/n1 [23], i_decinfo[3], \u_EXU_SCU/csr_rw [23]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u65  (\u_EXU_SCU/n1 [24], i_decinfo[3], \u_EXU_SCU/csr_rw [24]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u66  (\u_EXU_SCU/n1 [25], i_decinfo[3], \u_EXU_SCU/csr_rw [25]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u67  (\u_EXU_SCU/n1 [26], i_decinfo[3], \u_EXU_SCU/csr_rw [26]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u68  (\u_EXU_SCU/n1 [27], i_decinfo[3], \u_EXU_SCU/csr_rw [27]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u69  (\u_EXU_SCU/n1 [28], i_decinfo[3], \u_EXU_SCU/csr_rw [28]);  // ../RTL/core/exu_scu.v(55)
  not \u_EXU_SCU/u7  (\u_EXU_SCU/n0 [0], \u_EXU_SCU/csr_rw [0]);  // ../RTL/core/exu_scu.v(49)
  and \u_EXU_SCU/u70  (\u_EXU_SCU/n1 [29], i_decinfo[3], \u_EXU_SCU/csr_rw [29]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u71  (\u_EXU_SCU/n1 [30], i_decinfo[3], \u_EXU_SCU/csr_rw [30]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u72  (\u_EXU_SCU/n1 [31], i_decinfo[3], \u_EXU_SCU/csr_rw [31]);  // ../RTL/core/exu_scu.v(55)
  and \u_EXU_SCU/u8  (o_csr_wen, i_decinfo_grp[4], i_decinfo[7]);  // ../RTL/core/exu_scu.v(54)
  and \u_EXU_SCU/u9  (\u_EXU_SCU/n2 [6], i_decinfo[4], \u_EXU_SCU/csr_rs [6]);  // ../RTL/core/exu_scu.v(55)

endmodule 

module add_pu1_pu1_o1
  (
  i0,
  i1,
  o
  );

  input i0;
  input i1;
  output o;

  wire net_a0;
  wire net_cin;
  wire net_cout0;
  wire net_sum0;

  assign net_a0 = i0;
  assign net_cin = i1;
  assign o = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(1'b0),
    .c(net_cin),
    .cout(net_cout0),
    .sum(net_sum0));

endmodule 

module add_pu1_mu1_o1
  (
  i0,
  i1,
  o
  );

  input i0;
  input i1;
  output o;

  wire net_a0;
  wire net_cin;
  wire net_cout0;
  wire net_ncin;
  wire net_sum0;

  assign net_a0 = i0;
  assign net_cin = i1;
  assign o = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(1'b1),
    .c(net_ncin),
    .cout(net_cout0),
    .sum(net_sum0));
  not inv_cin (net_ncin, net_cin);

endmodule 

module add_pu30_pu30_o30
  (
  i0,
  i1,
  o
  );

  input [29:0] i0;
  input [29:0] i1;
  output [29:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module add_pu4_pu4_o4
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output [3:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;

  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));

endmodule 

module eq_w4
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output o;

  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;

  not none_diff (o, \or_or_xor_i0[0]_i1[0_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \xor_i0[3]_i1[3]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);

endmodule 

module add_pu4_mu4_o4
  (
  i0,
  i1,
  o
  );

  input [3:0] i0;
  input [3:0] i1;
  output [3:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_nb0;
  wire net_nb1;
  wire net_nb2;
  wire net_nb3;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;

  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b2 (net_nb2, net_b2);
  not inv_b3 (net_nb3, net_b3);

endmodule 

module eq_w5
  (
  i0,
  i1,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  output o;

  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;

  not none_diff (o, \or_or_xor_i0[0]_i1[0_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \xor_i0[4]_i1[4]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);

endmodule 

module ne_w5
  (
  i0,
  i1,
  o
  );

  input [4:0] i0;
  input [4:0] i1;
  output o;

  wire [4:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2], diff[3], diff[4]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_4 (diff[4], i0[4], i1[4]);

endmodule 

module add_pu32_pu32_o32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output [31:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_b23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_b24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_b25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_b26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_b27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_b28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_b29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_b30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_b31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module eq_w3
  (
  i0,
  i1,
  o
  );

  input [2:0] i0;
  input [2:0] i1;
  output o;

  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;

  not none_diff (o, \or_xor_i0[0]_i1[0]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);

endmodule 

module eq_w7
  (
  i0,
  i1,
  o
  );

  input [6:0] i0;
  input [6:0] i1;
  output o;

  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[3]_i1[3_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[5]_i1[5]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;

  not none_diff (o, \or_or_xor_i0[0]_i1[0_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_or_xor_i0[3]_i1[3_o );
  or \or_or_xor_i0[3]_i1[3  (\or_or_xor_i0[3]_i1[3_o , \or_xor_i0[3]_i1[3]_o_o , \or_xor_i0[5]_i1[5]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \xor_i0[4]_i1[4]_o );
  or \or_xor_i0[5]_i1[5]_o  (\or_xor_i0[5]_i1[5]_o_o , \xor_i0[5]_i1[5]_o , \xor_i0[6]_i1[6]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);

endmodule 

module eq_w12
  (
  i0,
  i1,
  o
  );

  input [11:0] i0;
  input [11:0] i1;
  output o;

  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[6]_i1[6_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[10]_i1[10]_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[7]_i1[7]_o_o ;
  wire \or_xor_i0[9]_i1[9]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, \or_or_or_xor_i0[0]_i_o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[6]_i1[6_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_or_xor_i0[6]_i1[6  (\or_or_xor_i0[6]_i1[6_o , \or_xor_i0[6]_i1[6]_o_o , \or_xor_i0[9]_i1[9]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[10]_i1[10]  (\or_xor_i0[10]_i1[10]_o , \xor_i0[10]_i1[10]_o , \xor_i0[11]_i1[11]_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \or_xor_i0[4]_i1[4]_o_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \or_xor_i0[7]_i1[7]_o_o );
  or \or_xor_i0[7]_i1[7]_o  (\or_xor_i0[7]_i1[7]_o_o , \xor_i0[7]_i1[7]_o , \xor_i0[8]_i1[8]_o );
  or \or_xor_i0[9]_i1[9]_o  (\or_xor_i0[9]_i1[9]_o_o , \xor_i0[9]_i1[9]_o , \or_xor_i0[10]_i1[10]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module REGFILE  // ../RTL/core/regfile.v(12)
  (
  i_clk,
  i_rd_wdata,
  i_rdidx,
  i_rdwen,
  i_rs1idx,
  i_rs1ren,
  i_rs2idx,
  i_rs2ren,
  i_rstn,
  o_rs1_rdata,
  o_rs2_rdata
  );

  input i_clk;  // ../RTL/core/regfile.v(13)
  input [31:0] i_rd_wdata;  // ../RTL/core/regfile.v(17)
  input [4:0] i_rdidx;  // ../RTL/core/regfile.v(16)
  input i_rdwen;  // ../RTL/core/regfile.v(15)
  input [4:0] i_rs1idx;  // ../RTL/core/regfile.v(19)
  input i_rs1ren;  // ../RTL/core/regfile.v(18)
  input [4:0] i_rs2idx;  // ../RTL/core/regfile.v(22)
  input i_rs2ren;  // ../RTL/core/regfile.v(21)
  input i_rstn;  // ../RTL/core/regfile.v(14)
  output [31:0] o_rs1_rdata;  // ../RTL/core/regfile.v(20)
  output [31:0] o_rs2_rdata;  // ../RTL/core/regfile.v(23)

  // localparam gen_regfile_rd[0].i = 0;
  // localparam gen_regfile_rd[10].i = 10;
  // localparam gen_regfile_rd[11].i = 11;
  // localparam gen_regfile_rd[12].i = 12;
  // localparam gen_regfile_rd[13].i = 13;
  // localparam gen_regfile_rd[14].i = 14;
  // localparam gen_regfile_rd[15].i = 15;
  // localparam gen_regfile_rd[16].i = 16;
  // localparam gen_regfile_rd[17].i = 17;
  // localparam gen_regfile_rd[18].i = 18;
  // localparam gen_regfile_rd[19].i = 19;
  // localparam gen_regfile_rd[1].i = 1;
  // localparam gen_regfile_rd[20].i = 20;
  // localparam gen_regfile_rd[21].i = 21;
  // localparam gen_regfile_rd[22].i = 22;
  // localparam gen_regfile_rd[23].i = 23;
  // localparam gen_regfile_rd[24].i = 24;
  // localparam gen_regfile_rd[25].i = 25;
  // localparam gen_regfile_rd[26].i = 26;
  // localparam gen_regfile_rd[27].i = 27;
  // localparam gen_regfile_rd[28].i = 28;
  // localparam gen_regfile_rd[29].i = 29;
  // localparam gen_regfile_rd[2].i = 2;
  // localparam gen_regfile_rd[30].i = 30;
  // localparam gen_regfile_rd[31].i = 31;
  // localparam gen_regfile_rd[3].i = 3;
  // localparam gen_regfile_rd[4].i = 4;
  // localparam gen_regfile_rd[5].i = 5;
  // localparam gen_regfile_rd[6].i = 6;
  // localparam gen_regfile_rd[7].i = 7;
  // localparam gen_regfile_rd[8].i = 8;
  // localparam gen_regfile_rd[9].i = 9;
  wire [31:0] n100;
  wire [31:0] n95;
  wire [31:0] n96;
  wire [31:0] n99;
  wire [31:0] \rfxs[10] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[11] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[12] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[13] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[14] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[15] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[16] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[17] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[18] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[19] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[1] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[20] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[21] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[22] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[23] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[24] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[25] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[26] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[27] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[28] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[29] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[2] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[30] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[31] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[3] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[4] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[5] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[6] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[7] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[8] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[9] ;  // ../RTL/core/regfile.v(27)
  wire n0;
  wire n1;
  wire n10;
  wire n12;
  wire n13;
  wire n15;
  wire n16;
  wire n18;
  wire n19;
  wire n21;
  wire n22;
  wire n24;
  wire n25;
  wire n27;
  wire n28;
  wire n3;
  wire n30;
  wire n31;
  wire n33;
  wire n34;
  wire n36;
  wire n37;
  wire n39;
  wire n4;
  wire n40;
  wire n42;
  wire n43;
  wire n45;
  wire n46;
  wire n48;
  wire n49;
  wire n51;
  wire n52;
  wire n54;
  wire n55;
  wire n57;
  wire n58;
  wire n6;
  wire n60;
  wire n61;
  wire n63;
  wire n64;
  wire n66;
  wire n67;
  wire n69;
  wire n7;
  wire n70;
  wire n72;
  wire n73;
  wire n75;
  wire n76;
  wire n78;
  wire n79;
  wire n81;
  wire n82;
  wire n84;
  wire n85;
  wire n87;
  wire n88;
  wire n9;
  wire n90;
  wire n91;
  wire n93;
  wire n94;
  wire n97;
  wire n98;

  eq_w5 eq0 (
    .i0(i_rdidx),
    .i1(5'b00001),
    .o(n0));  // ../RTL/core/regfile.v(37)
  eq_w5 eq1 (
    .i0(i_rdidx),
    .i1(5'b00010),
    .o(n3));  // ../RTL/core/regfile.v(37)
  eq_w5 eq10 (
    .i0(i_rdidx),
    .i1(5'b01011),
    .o(n30));  // ../RTL/core/regfile.v(37)
  eq_w5 eq11 (
    .i0(i_rdidx),
    .i1(5'b01100),
    .o(n33));  // ../RTL/core/regfile.v(37)
  eq_w5 eq12 (
    .i0(i_rdidx),
    .i1(5'b01101),
    .o(n36));  // ../RTL/core/regfile.v(37)
  eq_w5 eq13 (
    .i0(i_rdidx),
    .i1(5'b01110),
    .o(n39));  // ../RTL/core/regfile.v(37)
  eq_w5 eq14 (
    .i0(i_rdidx),
    .i1(5'b01111),
    .o(n42));  // ../RTL/core/regfile.v(37)
  eq_w5 eq15 (
    .i0(i_rdidx),
    .i1(5'b10000),
    .o(n45));  // ../RTL/core/regfile.v(37)
  eq_w5 eq16 (
    .i0(i_rdidx),
    .i1(5'b10001),
    .o(n48));  // ../RTL/core/regfile.v(37)
  eq_w5 eq17 (
    .i0(i_rdidx),
    .i1(5'b10010),
    .o(n51));  // ../RTL/core/regfile.v(37)
  eq_w5 eq18 (
    .i0(i_rdidx),
    .i1(5'b10011),
    .o(n54));  // ../RTL/core/regfile.v(37)
  eq_w5 eq19 (
    .i0(i_rdidx),
    .i1(5'b10100),
    .o(n57));  // ../RTL/core/regfile.v(37)
  eq_w5 eq2 (
    .i0(i_rdidx),
    .i1(5'b00011),
    .o(n6));  // ../RTL/core/regfile.v(37)
  eq_w5 eq20 (
    .i0(i_rdidx),
    .i1(5'b10101),
    .o(n60));  // ../RTL/core/regfile.v(37)
  eq_w5 eq21 (
    .i0(i_rdidx),
    .i1(5'b10110),
    .o(n63));  // ../RTL/core/regfile.v(37)
  eq_w5 eq22 (
    .i0(i_rdidx),
    .i1(5'b10111),
    .o(n66));  // ../RTL/core/regfile.v(37)
  eq_w5 eq23 (
    .i0(i_rdidx),
    .i1(5'b11000),
    .o(n69));  // ../RTL/core/regfile.v(37)
  eq_w5 eq24 (
    .i0(i_rdidx),
    .i1(5'b11001),
    .o(n72));  // ../RTL/core/regfile.v(37)
  eq_w5 eq25 (
    .i0(i_rdidx),
    .i1(5'b11010),
    .o(n75));  // ../RTL/core/regfile.v(37)
  eq_w5 eq26 (
    .i0(i_rdidx),
    .i1(5'b11011),
    .o(n78));  // ../RTL/core/regfile.v(37)
  eq_w5 eq27 (
    .i0(i_rdidx),
    .i1(5'b11100),
    .o(n81));  // ../RTL/core/regfile.v(37)
  eq_w5 eq28 (
    .i0(i_rdidx),
    .i1(5'b11101),
    .o(n84));  // ../RTL/core/regfile.v(37)
  eq_w5 eq29 (
    .i0(i_rdidx),
    .i1(5'b11110),
    .o(n87));  // ../RTL/core/regfile.v(37)
  eq_w5 eq3 (
    .i0(i_rdidx),
    .i1(5'b00100),
    .o(n9));  // ../RTL/core/regfile.v(37)
  eq_w5 eq30 (
    .i0(i_rdidx),
    .i1(5'b11111),
    .o(n90));  // ../RTL/core/regfile.v(37)
  eq_w5 eq31 (
    .i0(i_rs1idx),
    .i1(i_rdidx),
    .o(n93));  // ../RTL/core/regfile.v(46)
  eq_w5 eq32 (
    .i0(i_rs2idx),
    .i1(i_rdidx),
    .o(n97));  // ../RTL/core/regfile.v(47)
  eq_w5 eq4 (
    .i0(i_rdidx),
    .i1(5'b00101),
    .o(n12));  // ../RTL/core/regfile.v(37)
  eq_w5 eq5 (
    .i0(i_rdidx),
    .i1(5'b00110),
    .o(n15));  // ../RTL/core/regfile.v(37)
  eq_w5 eq6 (
    .i0(i_rdidx),
    .i1(5'b00111),
    .o(n18));  // ../RTL/core/regfile.v(37)
  eq_w5 eq7 (
    .i0(i_rdidx),
    .i1(5'b01000),
    .o(n21));  // ../RTL/core/regfile.v(37)
  eq_w5 eq8 (
    .i0(i_rdidx),
    .i1(5'b01001),
    .o(n24));  // ../RTL/core/regfile.v(37)
  eq_w5 eq9 (
    .i0(i_rdidx),
    .i1(5'b01010),
    .o(n27));  // ../RTL/core/regfile.v(37)
  binary_mux_s5_w1 mux31_b0 (
    .i0(1'b0),
    .i1(\rfxs[1] [0]),
    .i10(\rfxs[10] [0]),
    .i11(\rfxs[11] [0]),
    .i12(\rfxs[12] [0]),
    .i13(\rfxs[13] [0]),
    .i14(\rfxs[14] [0]),
    .i15(\rfxs[15] [0]),
    .i16(\rfxs[16] [0]),
    .i17(\rfxs[17] [0]),
    .i18(\rfxs[18] [0]),
    .i19(\rfxs[19] [0]),
    .i2(\rfxs[2] [0]),
    .i20(\rfxs[20] [0]),
    .i21(\rfxs[21] [0]),
    .i22(\rfxs[22] [0]),
    .i23(\rfxs[23] [0]),
    .i24(\rfxs[24] [0]),
    .i25(\rfxs[25] [0]),
    .i26(\rfxs[26] [0]),
    .i27(\rfxs[27] [0]),
    .i28(\rfxs[28] [0]),
    .i29(\rfxs[29] [0]),
    .i3(\rfxs[3] [0]),
    .i30(\rfxs[30] [0]),
    .i31(\rfxs[31] [0]),
    .i4(\rfxs[4] [0]),
    .i5(\rfxs[5] [0]),
    .i6(\rfxs[6] [0]),
    .i7(\rfxs[7] [0]),
    .i8(\rfxs[8] [0]),
    .i9(\rfxs[9] [0]),
    .sel(i_rs1idx),
    .o(n95[0]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b1 (
    .i0(1'b0),
    .i1(\rfxs[1] [1]),
    .i10(\rfxs[10] [1]),
    .i11(\rfxs[11] [1]),
    .i12(\rfxs[12] [1]),
    .i13(\rfxs[13] [1]),
    .i14(\rfxs[14] [1]),
    .i15(\rfxs[15] [1]),
    .i16(\rfxs[16] [1]),
    .i17(\rfxs[17] [1]),
    .i18(\rfxs[18] [1]),
    .i19(\rfxs[19] [1]),
    .i2(\rfxs[2] [1]),
    .i20(\rfxs[20] [1]),
    .i21(\rfxs[21] [1]),
    .i22(\rfxs[22] [1]),
    .i23(\rfxs[23] [1]),
    .i24(\rfxs[24] [1]),
    .i25(\rfxs[25] [1]),
    .i26(\rfxs[26] [1]),
    .i27(\rfxs[27] [1]),
    .i28(\rfxs[28] [1]),
    .i29(\rfxs[29] [1]),
    .i3(\rfxs[3] [1]),
    .i30(\rfxs[30] [1]),
    .i31(\rfxs[31] [1]),
    .i4(\rfxs[4] [1]),
    .i5(\rfxs[5] [1]),
    .i6(\rfxs[6] [1]),
    .i7(\rfxs[7] [1]),
    .i8(\rfxs[8] [1]),
    .i9(\rfxs[9] [1]),
    .sel(i_rs1idx),
    .o(n95[1]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b10 (
    .i0(1'b0),
    .i1(\rfxs[1] [10]),
    .i10(\rfxs[10] [10]),
    .i11(\rfxs[11] [10]),
    .i12(\rfxs[12] [10]),
    .i13(\rfxs[13] [10]),
    .i14(\rfxs[14] [10]),
    .i15(\rfxs[15] [10]),
    .i16(\rfxs[16] [10]),
    .i17(\rfxs[17] [10]),
    .i18(\rfxs[18] [10]),
    .i19(\rfxs[19] [10]),
    .i2(\rfxs[2] [10]),
    .i20(\rfxs[20] [10]),
    .i21(\rfxs[21] [10]),
    .i22(\rfxs[22] [10]),
    .i23(\rfxs[23] [10]),
    .i24(\rfxs[24] [10]),
    .i25(\rfxs[25] [10]),
    .i26(\rfxs[26] [10]),
    .i27(\rfxs[27] [10]),
    .i28(\rfxs[28] [10]),
    .i29(\rfxs[29] [10]),
    .i3(\rfxs[3] [10]),
    .i30(\rfxs[30] [10]),
    .i31(\rfxs[31] [10]),
    .i4(\rfxs[4] [10]),
    .i5(\rfxs[5] [10]),
    .i6(\rfxs[6] [10]),
    .i7(\rfxs[7] [10]),
    .i8(\rfxs[8] [10]),
    .i9(\rfxs[9] [10]),
    .sel(i_rs1idx),
    .o(n95[10]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b11 (
    .i0(1'b0),
    .i1(\rfxs[1] [11]),
    .i10(\rfxs[10] [11]),
    .i11(\rfxs[11] [11]),
    .i12(\rfxs[12] [11]),
    .i13(\rfxs[13] [11]),
    .i14(\rfxs[14] [11]),
    .i15(\rfxs[15] [11]),
    .i16(\rfxs[16] [11]),
    .i17(\rfxs[17] [11]),
    .i18(\rfxs[18] [11]),
    .i19(\rfxs[19] [11]),
    .i2(\rfxs[2] [11]),
    .i20(\rfxs[20] [11]),
    .i21(\rfxs[21] [11]),
    .i22(\rfxs[22] [11]),
    .i23(\rfxs[23] [11]),
    .i24(\rfxs[24] [11]),
    .i25(\rfxs[25] [11]),
    .i26(\rfxs[26] [11]),
    .i27(\rfxs[27] [11]),
    .i28(\rfxs[28] [11]),
    .i29(\rfxs[29] [11]),
    .i3(\rfxs[3] [11]),
    .i30(\rfxs[30] [11]),
    .i31(\rfxs[31] [11]),
    .i4(\rfxs[4] [11]),
    .i5(\rfxs[5] [11]),
    .i6(\rfxs[6] [11]),
    .i7(\rfxs[7] [11]),
    .i8(\rfxs[8] [11]),
    .i9(\rfxs[9] [11]),
    .sel(i_rs1idx),
    .o(n95[11]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b12 (
    .i0(1'b0),
    .i1(\rfxs[1] [12]),
    .i10(\rfxs[10] [12]),
    .i11(\rfxs[11] [12]),
    .i12(\rfxs[12] [12]),
    .i13(\rfxs[13] [12]),
    .i14(\rfxs[14] [12]),
    .i15(\rfxs[15] [12]),
    .i16(\rfxs[16] [12]),
    .i17(\rfxs[17] [12]),
    .i18(\rfxs[18] [12]),
    .i19(\rfxs[19] [12]),
    .i2(\rfxs[2] [12]),
    .i20(\rfxs[20] [12]),
    .i21(\rfxs[21] [12]),
    .i22(\rfxs[22] [12]),
    .i23(\rfxs[23] [12]),
    .i24(\rfxs[24] [12]),
    .i25(\rfxs[25] [12]),
    .i26(\rfxs[26] [12]),
    .i27(\rfxs[27] [12]),
    .i28(\rfxs[28] [12]),
    .i29(\rfxs[29] [12]),
    .i3(\rfxs[3] [12]),
    .i30(\rfxs[30] [12]),
    .i31(\rfxs[31] [12]),
    .i4(\rfxs[4] [12]),
    .i5(\rfxs[5] [12]),
    .i6(\rfxs[6] [12]),
    .i7(\rfxs[7] [12]),
    .i8(\rfxs[8] [12]),
    .i9(\rfxs[9] [12]),
    .sel(i_rs1idx),
    .o(n95[12]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b13 (
    .i0(1'b0),
    .i1(\rfxs[1] [13]),
    .i10(\rfxs[10] [13]),
    .i11(\rfxs[11] [13]),
    .i12(\rfxs[12] [13]),
    .i13(\rfxs[13] [13]),
    .i14(\rfxs[14] [13]),
    .i15(\rfxs[15] [13]),
    .i16(\rfxs[16] [13]),
    .i17(\rfxs[17] [13]),
    .i18(\rfxs[18] [13]),
    .i19(\rfxs[19] [13]),
    .i2(\rfxs[2] [13]),
    .i20(\rfxs[20] [13]),
    .i21(\rfxs[21] [13]),
    .i22(\rfxs[22] [13]),
    .i23(\rfxs[23] [13]),
    .i24(\rfxs[24] [13]),
    .i25(\rfxs[25] [13]),
    .i26(\rfxs[26] [13]),
    .i27(\rfxs[27] [13]),
    .i28(\rfxs[28] [13]),
    .i29(\rfxs[29] [13]),
    .i3(\rfxs[3] [13]),
    .i30(\rfxs[30] [13]),
    .i31(\rfxs[31] [13]),
    .i4(\rfxs[4] [13]),
    .i5(\rfxs[5] [13]),
    .i6(\rfxs[6] [13]),
    .i7(\rfxs[7] [13]),
    .i8(\rfxs[8] [13]),
    .i9(\rfxs[9] [13]),
    .sel(i_rs1idx),
    .o(n95[13]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b14 (
    .i0(1'b0),
    .i1(\rfxs[1] [14]),
    .i10(\rfxs[10] [14]),
    .i11(\rfxs[11] [14]),
    .i12(\rfxs[12] [14]),
    .i13(\rfxs[13] [14]),
    .i14(\rfxs[14] [14]),
    .i15(\rfxs[15] [14]),
    .i16(\rfxs[16] [14]),
    .i17(\rfxs[17] [14]),
    .i18(\rfxs[18] [14]),
    .i19(\rfxs[19] [14]),
    .i2(\rfxs[2] [14]),
    .i20(\rfxs[20] [14]),
    .i21(\rfxs[21] [14]),
    .i22(\rfxs[22] [14]),
    .i23(\rfxs[23] [14]),
    .i24(\rfxs[24] [14]),
    .i25(\rfxs[25] [14]),
    .i26(\rfxs[26] [14]),
    .i27(\rfxs[27] [14]),
    .i28(\rfxs[28] [14]),
    .i29(\rfxs[29] [14]),
    .i3(\rfxs[3] [14]),
    .i30(\rfxs[30] [14]),
    .i31(\rfxs[31] [14]),
    .i4(\rfxs[4] [14]),
    .i5(\rfxs[5] [14]),
    .i6(\rfxs[6] [14]),
    .i7(\rfxs[7] [14]),
    .i8(\rfxs[8] [14]),
    .i9(\rfxs[9] [14]),
    .sel(i_rs1idx),
    .o(n95[14]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b15 (
    .i0(1'b0),
    .i1(\rfxs[1] [15]),
    .i10(\rfxs[10] [15]),
    .i11(\rfxs[11] [15]),
    .i12(\rfxs[12] [15]),
    .i13(\rfxs[13] [15]),
    .i14(\rfxs[14] [15]),
    .i15(\rfxs[15] [15]),
    .i16(\rfxs[16] [15]),
    .i17(\rfxs[17] [15]),
    .i18(\rfxs[18] [15]),
    .i19(\rfxs[19] [15]),
    .i2(\rfxs[2] [15]),
    .i20(\rfxs[20] [15]),
    .i21(\rfxs[21] [15]),
    .i22(\rfxs[22] [15]),
    .i23(\rfxs[23] [15]),
    .i24(\rfxs[24] [15]),
    .i25(\rfxs[25] [15]),
    .i26(\rfxs[26] [15]),
    .i27(\rfxs[27] [15]),
    .i28(\rfxs[28] [15]),
    .i29(\rfxs[29] [15]),
    .i3(\rfxs[3] [15]),
    .i30(\rfxs[30] [15]),
    .i31(\rfxs[31] [15]),
    .i4(\rfxs[4] [15]),
    .i5(\rfxs[5] [15]),
    .i6(\rfxs[6] [15]),
    .i7(\rfxs[7] [15]),
    .i8(\rfxs[8] [15]),
    .i9(\rfxs[9] [15]),
    .sel(i_rs1idx),
    .o(n95[15]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b16 (
    .i0(1'b0),
    .i1(\rfxs[1] [16]),
    .i10(\rfxs[10] [16]),
    .i11(\rfxs[11] [16]),
    .i12(\rfxs[12] [16]),
    .i13(\rfxs[13] [16]),
    .i14(\rfxs[14] [16]),
    .i15(\rfxs[15] [16]),
    .i16(\rfxs[16] [16]),
    .i17(\rfxs[17] [16]),
    .i18(\rfxs[18] [16]),
    .i19(\rfxs[19] [16]),
    .i2(\rfxs[2] [16]),
    .i20(\rfxs[20] [16]),
    .i21(\rfxs[21] [16]),
    .i22(\rfxs[22] [16]),
    .i23(\rfxs[23] [16]),
    .i24(\rfxs[24] [16]),
    .i25(\rfxs[25] [16]),
    .i26(\rfxs[26] [16]),
    .i27(\rfxs[27] [16]),
    .i28(\rfxs[28] [16]),
    .i29(\rfxs[29] [16]),
    .i3(\rfxs[3] [16]),
    .i30(\rfxs[30] [16]),
    .i31(\rfxs[31] [16]),
    .i4(\rfxs[4] [16]),
    .i5(\rfxs[5] [16]),
    .i6(\rfxs[6] [16]),
    .i7(\rfxs[7] [16]),
    .i8(\rfxs[8] [16]),
    .i9(\rfxs[9] [16]),
    .sel(i_rs1idx),
    .o(n95[16]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b17 (
    .i0(1'b0),
    .i1(\rfxs[1] [17]),
    .i10(\rfxs[10] [17]),
    .i11(\rfxs[11] [17]),
    .i12(\rfxs[12] [17]),
    .i13(\rfxs[13] [17]),
    .i14(\rfxs[14] [17]),
    .i15(\rfxs[15] [17]),
    .i16(\rfxs[16] [17]),
    .i17(\rfxs[17] [17]),
    .i18(\rfxs[18] [17]),
    .i19(\rfxs[19] [17]),
    .i2(\rfxs[2] [17]),
    .i20(\rfxs[20] [17]),
    .i21(\rfxs[21] [17]),
    .i22(\rfxs[22] [17]),
    .i23(\rfxs[23] [17]),
    .i24(\rfxs[24] [17]),
    .i25(\rfxs[25] [17]),
    .i26(\rfxs[26] [17]),
    .i27(\rfxs[27] [17]),
    .i28(\rfxs[28] [17]),
    .i29(\rfxs[29] [17]),
    .i3(\rfxs[3] [17]),
    .i30(\rfxs[30] [17]),
    .i31(\rfxs[31] [17]),
    .i4(\rfxs[4] [17]),
    .i5(\rfxs[5] [17]),
    .i6(\rfxs[6] [17]),
    .i7(\rfxs[7] [17]),
    .i8(\rfxs[8] [17]),
    .i9(\rfxs[9] [17]),
    .sel(i_rs1idx),
    .o(n95[17]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b18 (
    .i0(1'b0),
    .i1(\rfxs[1] [18]),
    .i10(\rfxs[10] [18]),
    .i11(\rfxs[11] [18]),
    .i12(\rfxs[12] [18]),
    .i13(\rfxs[13] [18]),
    .i14(\rfxs[14] [18]),
    .i15(\rfxs[15] [18]),
    .i16(\rfxs[16] [18]),
    .i17(\rfxs[17] [18]),
    .i18(\rfxs[18] [18]),
    .i19(\rfxs[19] [18]),
    .i2(\rfxs[2] [18]),
    .i20(\rfxs[20] [18]),
    .i21(\rfxs[21] [18]),
    .i22(\rfxs[22] [18]),
    .i23(\rfxs[23] [18]),
    .i24(\rfxs[24] [18]),
    .i25(\rfxs[25] [18]),
    .i26(\rfxs[26] [18]),
    .i27(\rfxs[27] [18]),
    .i28(\rfxs[28] [18]),
    .i29(\rfxs[29] [18]),
    .i3(\rfxs[3] [18]),
    .i30(\rfxs[30] [18]),
    .i31(\rfxs[31] [18]),
    .i4(\rfxs[4] [18]),
    .i5(\rfxs[5] [18]),
    .i6(\rfxs[6] [18]),
    .i7(\rfxs[7] [18]),
    .i8(\rfxs[8] [18]),
    .i9(\rfxs[9] [18]),
    .sel(i_rs1idx),
    .o(n95[18]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b19 (
    .i0(1'b0),
    .i1(\rfxs[1] [19]),
    .i10(\rfxs[10] [19]),
    .i11(\rfxs[11] [19]),
    .i12(\rfxs[12] [19]),
    .i13(\rfxs[13] [19]),
    .i14(\rfxs[14] [19]),
    .i15(\rfxs[15] [19]),
    .i16(\rfxs[16] [19]),
    .i17(\rfxs[17] [19]),
    .i18(\rfxs[18] [19]),
    .i19(\rfxs[19] [19]),
    .i2(\rfxs[2] [19]),
    .i20(\rfxs[20] [19]),
    .i21(\rfxs[21] [19]),
    .i22(\rfxs[22] [19]),
    .i23(\rfxs[23] [19]),
    .i24(\rfxs[24] [19]),
    .i25(\rfxs[25] [19]),
    .i26(\rfxs[26] [19]),
    .i27(\rfxs[27] [19]),
    .i28(\rfxs[28] [19]),
    .i29(\rfxs[29] [19]),
    .i3(\rfxs[3] [19]),
    .i30(\rfxs[30] [19]),
    .i31(\rfxs[31] [19]),
    .i4(\rfxs[4] [19]),
    .i5(\rfxs[5] [19]),
    .i6(\rfxs[6] [19]),
    .i7(\rfxs[7] [19]),
    .i8(\rfxs[8] [19]),
    .i9(\rfxs[9] [19]),
    .sel(i_rs1idx),
    .o(n95[19]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b2 (
    .i0(1'b0),
    .i1(\rfxs[1] [2]),
    .i10(\rfxs[10] [2]),
    .i11(\rfxs[11] [2]),
    .i12(\rfxs[12] [2]),
    .i13(\rfxs[13] [2]),
    .i14(\rfxs[14] [2]),
    .i15(\rfxs[15] [2]),
    .i16(\rfxs[16] [2]),
    .i17(\rfxs[17] [2]),
    .i18(\rfxs[18] [2]),
    .i19(\rfxs[19] [2]),
    .i2(\rfxs[2] [2]),
    .i20(\rfxs[20] [2]),
    .i21(\rfxs[21] [2]),
    .i22(\rfxs[22] [2]),
    .i23(\rfxs[23] [2]),
    .i24(\rfxs[24] [2]),
    .i25(\rfxs[25] [2]),
    .i26(\rfxs[26] [2]),
    .i27(\rfxs[27] [2]),
    .i28(\rfxs[28] [2]),
    .i29(\rfxs[29] [2]),
    .i3(\rfxs[3] [2]),
    .i30(\rfxs[30] [2]),
    .i31(\rfxs[31] [2]),
    .i4(\rfxs[4] [2]),
    .i5(\rfxs[5] [2]),
    .i6(\rfxs[6] [2]),
    .i7(\rfxs[7] [2]),
    .i8(\rfxs[8] [2]),
    .i9(\rfxs[9] [2]),
    .sel(i_rs1idx),
    .o(n95[2]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b20 (
    .i0(1'b0),
    .i1(\rfxs[1] [20]),
    .i10(\rfxs[10] [20]),
    .i11(\rfxs[11] [20]),
    .i12(\rfxs[12] [20]),
    .i13(\rfxs[13] [20]),
    .i14(\rfxs[14] [20]),
    .i15(\rfxs[15] [20]),
    .i16(\rfxs[16] [20]),
    .i17(\rfxs[17] [20]),
    .i18(\rfxs[18] [20]),
    .i19(\rfxs[19] [20]),
    .i2(\rfxs[2] [20]),
    .i20(\rfxs[20] [20]),
    .i21(\rfxs[21] [20]),
    .i22(\rfxs[22] [20]),
    .i23(\rfxs[23] [20]),
    .i24(\rfxs[24] [20]),
    .i25(\rfxs[25] [20]),
    .i26(\rfxs[26] [20]),
    .i27(\rfxs[27] [20]),
    .i28(\rfxs[28] [20]),
    .i29(\rfxs[29] [20]),
    .i3(\rfxs[3] [20]),
    .i30(\rfxs[30] [20]),
    .i31(\rfxs[31] [20]),
    .i4(\rfxs[4] [20]),
    .i5(\rfxs[5] [20]),
    .i6(\rfxs[6] [20]),
    .i7(\rfxs[7] [20]),
    .i8(\rfxs[8] [20]),
    .i9(\rfxs[9] [20]),
    .sel(i_rs1idx),
    .o(n95[20]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b21 (
    .i0(1'b0),
    .i1(\rfxs[1] [21]),
    .i10(\rfxs[10] [21]),
    .i11(\rfxs[11] [21]),
    .i12(\rfxs[12] [21]),
    .i13(\rfxs[13] [21]),
    .i14(\rfxs[14] [21]),
    .i15(\rfxs[15] [21]),
    .i16(\rfxs[16] [21]),
    .i17(\rfxs[17] [21]),
    .i18(\rfxs[18] [21]),
    .i19(\rfxs[19] [21]),
    .i2(\rfxs[2] [21]),
    .i20(\rfxs[20] [21]),
    .i21(\rfxs[21] [21]),
    .i22(\rfxs[22] [21]),
    .i23(\rfxs[23] [21]),
    .i24(\rfxs[24] [21]),
    .i25(\rfxs[25] [21]),
    .i26(\rfxs[26] [21]),
    .i27(\rfxs[27] [21]),
    .i28(\rfxs[28] [21]),
    .i29(\rfxs[29] [21]),
    .i3(\rfxs[3] [21]),
    .i30(\rfxs[30] [21]),
    .i31(\rfxs[31] [21]),
    .i4(\rfxs[4] [21]),
    .i5(\rfxs[5] [21]),
    .i6(\rfxs[6] [21]),
    .i7(\rfxs[7] [21]),
    .i8(\rfxs[8] [21]),
    .i9(\rfxs[9] [21]),
    .sel(i_rs1idx),
    .o(n95[21]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b22 (
    .i0(1'b0),
    .i1(\rfxs[1] [22]),
    .i10(\rfxs[10] [22]),
    .i11(\rfxs[11] [22]),
    .i12(\rfxs[12] [22]),
    .i13(\rfxs[13] [22]),
    .i14(\rfxs[14] [22]),
    .i15(\rfxs[15] [22]),
    .i16(\rfxs[16] [22]),
    .i17(\rfxs[17] [22]),
    .i18(\rfxs[18] [22]),
    .i19(\rfxs[19] [22]),
    .i2(\rfxs[2] [22]),
    .i20(\rfxs[20] [22]),
    .i21(\rfxs[21] [22]),
    .i22(\rfxs[22] [22]),
    .i23(\rfxs[23] [22]),
    .i24(\rfxs[24] [22]),
    .i25(\rfxs[25] [22]),
    .i26(\rfxs[26] [22]),
    .i27(\rfxs[27] [22]),
    .i28(\rfxs[28] [22]),
    .i29(\rfxs[29] [22]),
    .i3(\rfxs[3] [22]),
    .i30(\rfxs[30] [22]),
    .i31(\rfxs[31] [22]),
    .i4(\rfxs[4] [22]),
    .i5(\rfxs[5] [22]),
    .i6(\rfxs[6] [22]),
    .i7(\rfxs[7] [22]),
    .i8(\rfxs[8] [22]),
    .i9(\rfxs[9] [22]),
    .sel(i_rs1idx),
    .o(n95[22]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b23 (
    .i0(1'b0),
    .i1(\rfxs[1] [23]),
    .i10(\rfxs[10] [23]),
    .i11(\rfxs[11] [23]),
    .i12(\rfxs[12] [23]),
    .i13(\rfxs[13] [23]),
    .i14(\rfxs[14] [23]),
    .i15(\rfxs[15] [23]),
    .i16(\rfxs[16] [23]),
    .i17(\rfxs[17] [23]),
    .i18(\rfxs[18] [23]),
    .i19(\rfxs[19] [23]),
    .i2(\rfxs[2] [23]),
    .i20(\rfxs[20] [23]),
    .i21(\rfxs[21] [23]),
    .i22(\rfxs[22] [23]),
    .i23(\rfxs[23] [23]),
    .i24(\rfxs[24] [23]),
    .i25(\rfxs[25] [23]),
    .i26(\rfxs[26] [23]),
    .i27(\rfxs[27] [23]),
    .i28(\rfxs[28] [23]),
    .i29(\rfxs[29] [23]),
    .i3(\rfxs[3] [23]),
    .i30(\rfxs[30] [23]),
    .i31(\rfxs[31] [23]),
    .i4(\rfxs[4] [23]),
    .i5(\rfxs[5] [23]),
    .i6(\rfxs[6] [23]),
    .i7(\rfxs[7] [23]),
    .i8(\rfxs[8] [23]),
    .i9(\rfxs[9] [23]),
    .sel(i_rs1idx),
    .o(n95[23]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b24 (
    .i0(1'b0),
    .i1(\rfxs[1] [24]),
    .i10(\rfxs[10] [24]),
    .i11(\rfxs[11] [24]),
    .i12(\rfxs[12] [24]),
    .i13(\rfxs[13] [24]),
    .i14(\rfxs[14] [24]),
    .i15(\rfxs[15] [24]),
    .i16(\rfxs[16] [24]),
    .i17(\rfxs[17] [24]),
    .i18(\rfxs[18] [24]),
    .i19(\rfxs[19] [24]),
    .i2(\rfxs[2] [24]),
    .i20(\rfxs[20] [24]),
    .i21(\rfxs[21] [24]),
    .i22(\rfxs[22] [24]),
    .i23(\rfxs[23] [24]),
    .i24(\rfxs[24] [24]),
    .i25(\rfxs[25] [24]),
    .i26(\rfxs[26] [24]),
    .i27(\rfxs[27] [24]),
    .i28(\rfxs[28] [24]),
    .i29(\rfxs[29] [24]),
    .i3(\rfxs[3] [24]),
    .i30(\rfxs[30] [24]),
    .i31(\rfxs[31] [24]),
    .i4(\rfxs[4] [24]),
    .i5(\rfxs[5] [24]),
    .i6(\rfxs[6] [24]),
    .i7(\rfxs[7] [24]),
    .i8(\rfxs[8] [24]),
    .i9(\rfxs[9] [24]),
    .sel(i_rs1idx),
    .o(n95[24]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b25 (
    .i0(1'b0),
    .i1(\rfxs[1] [25]),
    .i10(\rfxs[10] [25]),
    .i11(\rfxs[11] [25]),
    .i12(\rfxs[12] [25]),
    .i13(\rfxs[13] [25]),
    .i14(\rfxs[14] [25]),
    .i15(\rfxs[15] [25]),
    .i16(\rfxs[16] [25]),
    .i17(\rfxs[17] [25]),
    .i18(\rfxs[18] [25]),
    .i19(\rfxs[19] [25]),
    .i2(\rfxs[2] [25]),
    .i20(\rfxs[20] [25]),
    .i21(\rfxs[21] [25]),
    .i22(\rfxs[22] [25]),
    .i23(\rfxs[23] [25]),
    .i24(\rfxs[24] [25]),
    .i25(\rfxs[25] [25]),
    .i26(\rfxs[26] [25]),
    .i27(\rfxs[27] [25]),
    .i28(\rfxs[28] [25]),
    .i29(\rfxs[29] [25]),
    .i3(\rfxs[3] [25]),
    .i30(\rfxs[30] [25]),
    .i31(\rfxs[31] [25]),
    .i4(\rfxs[4] [25]),
    .i5(\rfxs[5] [25]),
    .i6(\rfxs[6] [25]),
    .i7(\rfxs[7] [25]),
    .i8(\rfxs[8] [25]),
    .i9(\rfxs[9] [25]),
    .sel(i_rs1idx),
    .o(n95[25]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b26 (
    .i0(1'b0),
    .i1(\rfxs[1] [26]),
    .i10(\rfxs[10] [26]),
    .i11(\rfxs[11] [26]),
    .i12(\rfxs[12] [26]),
    .i13(\rfxs[13] [26]),
    .i14(\rfxs[14] [26]),
    .i15(\rfxs[15] [26]),
    .i16(\rfxs[16] [26]),
    .i17(\rfxs[17] [26]),
    .i18(\rfxs[18] [26]),
    .i19(\rfxs[19] [26]),
    .i2(\rfxs[2] [26]),
    .i20(\rfxs[20] [26]),
    .i21(\rfxs[21] [26]),
    .i22(\rfxs[22] [26]),
    .i23(\rfxs[23] [26]),
    .i24(\rfxs[24] [26]),
    .i25(\rfxs[25] [26]),
    .i26(\rfxs[26] [26]),
    .i27(\rfxs[27] [26]),
    .i28(\rfxs[28] [26]),
    .i29(\rfxs[29] [26]),
    .i3(\rfxs[3] [26]),
    .i30(\rfxs[30] [26]),
    .i31(\rfxs[31] [26]),
    .i4(\rfxs[4] [26]),
    .i5(\rfxs[5] [26]),
    .i6(\rfxs[6] [26]),
    .i7(\rfxs[7] [26]),
    .i8(\rfxs[8] [26]),
    .i9(\rfxs[9] [26]),
    .sel(i_rs1idx),
    .o(n95[26]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b27 (
    .i0(1'b0),
    .i1(\rfxs[1] [27]),
    .i10(\rfxs[10] [27]),
    .i11(\rfxs[11] [27]),
    .i12(\rfxs[12] [27]),
    .i13(\rfxs[13] [27]),
    .i14(\rfxs[14] [27]),
    .i15(\rfxs[15] [27]),
    .i16(\rfxs[16] [27]),
    .i17(\rfxs[17] [27]),
    .i18(\rfxs[18] [27]),
    .i19(\rfxs[19] [27]),
    .i2(\rfxs[2] [27]),
    .i20(\rfxs[20] [27]),
    .i21(\rfxs[21] [27]),
    .i22(\rfxs[22] [27]),
    .i23(\rfxs[23] [27]),
    .i24(\rfxs[24] [27]),
    .i25(\rfxs[25] [27]),
    .i26(\rfxs[26] [27]),
    .i27(\rfxs[27] [27]),
    .i28(\rfxs[28] [27]),
    .i29(\rfxs[29] [27]),
    .i3(\rfxs[3] [27]),
    .i30(\rfxs[30] [27]),
    .i31(\rfxs[31] [27]),
    .i4(\rfxs[4] [27]),
    .i5(\rfxs[5] [27]),
    .i6(\rfxs[6] [27]),
    .i7(\rfxs[7] [27]),
    .i8(\rfxs[8] [27]),
    .i9(\rfxs[9] [27]),
    .sel(i_rs1idx),
    .o(n95[27]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b28 (
    .i0(1'b0),
    .i1(\rfxs[1] [28]),
    .i10(\rfxs[10] [28]),
    .i11(\rfxs[11] [28]),
    .i12(\rfxs[12] [28]),
    .i13(\rfxs[13] [28]),
    .i14(\rfxs[14] [28]),
    .i15(\rfxs[15] [28]),
    .i16(\rfxs[16] [28]),
    .i17(\rfxs[17] [28]),
    .i18(\rfxs[18] [28]),
    .i19(\rfxs[19] [28]),
    .i2(\rfxs[2] [28]),
    .i20(\rfxs[20] [28]),
    .i21(\rfxs[21] [28]),
    .i22(\rfxs[22] [28]),
    .i23(\rfxs[23] [28]),
    .i24(\rfxs[24] [28]),
    .i25(\rfxs[25] [28]),
    .i26(\rfxs[26] [28]),
    .i27(\rfxs[27] [28]),
    .i28(\rfxs[28] [28]),
    .i29(\rfxs[29] [28]),
    .i3(\rfxs[3] [28]),
    .i30(\rfxs[30] [28]),
    .i31(\rfxs[31] [28]),
    .i4(\rfxs[4] [28]),
    .i5(\rfxs[5] [28]),
    .i6(\rfxs[6] [28]),
    .i7(\rfxs[7] [28]),
    .i8(\rfxs[8] [28]),
    .i9(\rfxs[9] [28]),
    .sel(i_rs1idx),
    .o(n95[28]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b29 (
    .i0(1'b0),
    .i1(\rfxs[1] [29]),
    .i10(\rfxs[10] [29]),
    .i11(\rfxs[11] [29]),
    .i12(\rfxs[12] [29]),
    .i13(\rfxs[13] [29]),
    .i14(\rfxs[14] [29]),
    .i15(\rfxs[15] [29]),
    .i16(\rfxs[16] [29]),
    .i17(\rfxs[17] [29]),
    .i18(\rfxs[18] [29]),
    .i19(\rfxs[19] [29]),
    .i2(\rfxs[2] [29]),
    .i20(\rfxs[20] [29]),
    .i21(\rfxs[21] [29]),
    .i22(\rfxs[22] [29]),
    .i23(\rfxs[23] [29]),
    .i24(\rfxs[24] [29]),
    .i25(\rfxs[25] [29]),
    .i26(\rfxs[26] [29]),
    .i27(\rfxs[27] [29]),
    .i28(\rfxs[28] [29]),
    .i29(\rfxs[29] [29]),
    .i3(\rfxs[3] [29]),
    .i30(\rfxs[30] [29]),
    .i31(\rfxs[31] [29]),
    .i4(\rfxs[4] [29]),
    .i5(\rfxs[5] [29]),
    .i6(\rfxs[6] [29]),
    .i7(\rfxs[7] [29]),
    .i8(\rfxs[8] [29]),
    .i9(\rfxs[9] [29]),
    .sel(i_rs1idx),
    .o(n95[29]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b3 (
    .i0(1'b0),
    .i1(\rfxs[1] [3]),
    .i10(\rfxs[10] [3]),
    .i11(\rfxs[11] [3]),
    .i12(\rfxs[12] [3]),
    .i13(\rfxs[13] [3]),
    .i14(\rfxs[14] [3]),
    .i15(\rfxs[15] [3]),
    .i16(\rfxs[16] [3]),
    .i17(\rfxs[17] [3]),
    .i18(\rfxs[18] [3]),
    .i19(\rfxs[19] [3]),
    .i2(\rfxs[2] [3]),
    .i20(\rfxs[20] [3]),
    .i21(\rfxs[21] [3]),
    .i22(\rfxs[22] [3]),
    .i23(\rfxs[23] [3]),
    .i24(\rfxs[24] [3]),
    .i25(\rfxs[25] [3]),
    .i26(\rfxs[26] [3]),
    .i27(\rfxs[27] [3]),
    .i28(\rfxs[28] [3]),
    .i29(\rfxs[29] [3]),
    .i3(\rfxs[3] [3]),
    .i30(\rfxs[30] [3]),
    .i31(\rfxs[31] [3]),
    .i4(\rfxs[4] [3]),
    .i5(\rfxs[5] [3]),
    .i6(\rfxs[6] [3]),
    .i7(\rfxs[7] [3]),
    .i8(\rfxs[8] [3]),
    .i9(\rfxs[9] [3]),
    .sel(i_rs1idx),
    .o(n95[3]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b30 (
    .i0(1'b0),
    .i1(\rfxs[1] [30]),
    .i10(\rfxs[10] [30]),
    .i11(\rfxs[11] [30]),
    .i12(\rfxs[12] [30]),
    .i13(\rfxs[13] [30]),
    .i14(\rfxs[14] [30]),
    .i15(\rfxs[15] [30]),
    .i16(\rfxs[16] [30]),
    .i17(\rfxs[17] [30]),
    .i18(\rfxs[18] [30]),
    .i19(\rfxs[19] [30]),
    .i2(\rfxs[2] [30]),
    .i20(\rfxs[20] [30]),
    .i21(\rfxs[21] [30]),
    .i22(\rfxs[22] [30]),
    .i23(\rfxs[23] [30]),
    .i24(\rfxs[24] [30]),
    .i25(\rfxs[25] [30]),
    .i26(\rfxs[26] [30]),
    .i27(\rfxs[27] [30]),
    .i28(\rfxs[28] [30]),
    .i29(\rfxs[29] [30]),
    .i3(\rfxs[3] [30]),
    .i30(\rfxs[30] [30]),
    .i31(\rfxs[31] [30]),
    .i4(\rfxs[4] [30]),
    .i5(\rfxs[5] [30]),
    .i6(\rfxs[6] [30]),
    .i7(\rfxs[7] [30]),
    .i8(\rfxs[8] [30]),
    .i9(\rfxs[9] [30]),
    .sel(i_rs1idx),
    .o(n95[30]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b31 (
    .i0(1'b0),
    .i1(\rfxs[1] [31]),
    .i10(\rfxs[10] [31]),
    .i11(\rfxs[11] [31]),
    .i12(\rfxs[12] [31]),
    .i13(\rfxs[13] [31]),
    .i14(\rfxs[14] [31]),
    .i15(\rfxs[15] [31]),
    .i16(\rfxs[16] [31]),
    .i17(\rfxs[17] [31]),
    .i18(\rfxs[18] [31]),
    .i19(\rfxs[19] [31]),
    .i2(\rfxs[2] [31]),
    .i20(\rfxs[20] [31]),
    .i21(\rfxs[21] [31]),
    .i22(\rfxs[22] [31]),
    .i23(\rfxs[23] [31]),
    .i24(\rfxs[24] [31]),
    .i25(\rfxs[25] [31]),
    .i26(\rfxs[26] [31]),
    .i27(\rfxs[27] [31]),
    .i28(\rfxs[28] [31]),
    .i29(\rfxs[29] [31]),
    .i3(\rfxs[3] [31]),
    .i30(\rfxs[30] [31]),
    .i31(\rfxs[31] [31]),
    .i4(\rfxs[4] [31]),
    .i5(\rfxs[5] [31]),
    .i6(\rfxs[6] [31]),
    .i7(\rfxs[7] [31]),
    .i8(\rfxs[8] [31]),
    .i9(\rfxs[9] [31]),
    .sel(i_rs1idx),
    .o(n95[31]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b4 (
    .i0(1'b0),
    .i1(\rfxs[1] [4]),
    .i10(\rfxs[10] [4]),
    .i11(\rfxs[11] [4]),
    .i12(\rfxs[12] [4]),
    .i13(\rfxs[13] [4]),
    .i14(\rfxs[14] [4]),
    .i15(\rfxs[15] [4]),
    .i16(\rfxs[16] [4]),
    .i17(\rfxs[17] [4]),
    .i18(\rfxs[18] [4]),
    .i19(\rfxs[19] [4]),
    .i2(\rfxs[2] [4]),
    .i20(\rfxs[20] [4]),
    .i21(\rfxs[21] [4]),
    .i22(\rfxs[22] [4]),
    .i23(\rfxs[23] [4]),
    .i24(\rfxs[24] [4]),
    .i25(\rfxs[25] [4]),
    .i26(\rfxs[26] [4]),
    .i27(\rfxs[27] [4]),
    .i28(\rfxs[28] [4]),
    .i29(\rfxs[29] [4]),
    .i3(\rfxs[3] [4]),
    .i30(\rfxs[30] [4]),
    .i31(\rfxs[31] [4]),
    .i4(\rfxs[4] [4]),
    .i5(\rfxs[5] [4]),
    .i6(\rfxs[6] [4]),
    .i7(\rfxs[7] [4]),
    .i8(\rfxs[8] [4]),
    .i9(\rfxs[9] [4]),
    .sel(i_rs1idx),
    .o(n95[4]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b5 (
    .i0(1'b0),
    .i1(\rfxs[1] [5]),
    .i10(\rfxs[10] [5]),
    .i11(\rfxs[11] [5]),
    .i12(\rfxs[12] [5]),
    .i13(\rfxs[13] [5]),
    .i14(\rfxs[14] [5]),
    .i15(\rfxs[15] [5]),
    .i16(\rfxs[16] [5]),
    .i17(\rfxs[17] [5]),
    .i18(\rfxs[18] [5]),
    .i19(\rfxs[19] [5]),
    .i2(\rfxs[2] [5]),
    .i20(\rfxs[20] [5]),
    .i21(\rfxs[21] [5]),
    .i22(\rfxs[22] [5]),
    .i23(\rfxs[23] [5]),
    .i24(\rfxs[24] [5]),
    .i25(\rfxs[25] [5]),
    .i26(\rfxs[26] [5]),
    .i27(\rfxs[27] [5]),
    .i28(\rfxs[28] [5]),
    .i29(\rfxs[29] [5]),
    .i3(\rfxs[3] [5]),
    .i30(\rfxs[30] [5]),
    .i31(\rfxs[31] [5]),
    .i4(\rfxs[4] [5]),
    .i5(\rfxs[5] [5]),
    .i6(\rfxs[6] [5]),
    .i7(\rfxs[7] [5]),
    .i8(\rfxs[8] [5]),
    .i9(\rfxs[9] [5]),
    .sel(i_rs1idx),
    .o(n95[5]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b6 (
    .i0(1'b0),
    .i1(\rfxs[1] [6]),
    .i10(\rfxs[10] [6]),
    .i11(\rfxs[11] [6]),
    .i12(\rfxs[12] [6]),
    .i13(\rfxs[13] [6]),
    .i14(\rfxs[14] [6]),
    .i15(\rfxs[15] [6]),
    .i16(\rfxs[16] [6]),
    .i17(\rfxs[17] [6]),
    .i18(\rfxs[18] [6]),
    .i19(\rfxs[19] [6]),
    .i2(\rfxs[2] [6]),
    .i20(\rfxs[20] [6]),
    .i21(\rfxs[21] [6]),
    .i22(\rfxs[22] [6]),
    .i23(\rfxs[23] [6]),
    .i24(\rfxs[24] [6]),
    .i25(\rfxs[25] [6]),
    .i26(\rfxs[26] [6]),
    .i27(\rfxs[27] [6]),
    .i28(\rfxs[28] [6]),
    .i29(\rfxs[29] [6]),
    .i3(\rfxs[3] [6]),
    .i30(\rfxs[30] [6]),
    .i31(\rfxs[31] [6]),
    .i4(\rfxs[4] [6]),
    .i5(\rfxs[5] [6]),
    .i6(\rfxs[6] [6]),
    .i7(\rfxs[7] [6]),
    .i8(\rfxs[8] [6]),
    .i9(\rfxs[9] [6]),
    .sel(i_rs1idx),
    .o(n95[6]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b7 (
    .i0(1'b0),
    .i1(\rfxs[1] [7]),
    .i10(\rfxs[10] [7]),
    .i11(\rfxs[11] [7]),
    .i12(\rfxs[12] [7]),
    .i13(\rfxs[13] [7]),
    .i14(\rfxs[14] [7]),
    .i15(\rfxs[15] [7]),
    .i16(\rfxs[16] [7]),
    .i17(\rfxs[17] [7]),
    .i18(\rfxs[18] [7]),
    .i19(\rfxs[19] [7]),
    .i2(\rfxs[2] [7]),
    .i20(\rfxs[20] [7]),
    .i21(\rfxs[21] [7]),
    .i22(\rfxs[22] [7]),
    .i23(\rfxs[23] [7]),
    .i24(\rfxs[24] [7]),
    .i25(\rfxs[25] [7]),
    .i26(\rfxs[26] [7]),
    .i27(\rfxs[27] [7]),
    .i28(\rfxs[28] [7]),
    .i29(\rfxs[29] [7]),
    .i3(\rfxs[3] [7]),
    .i30(\rfxs[30] [7]),
    .i31(\rfxs[31] [7]),
    .i4(\rfxs[4] [7]),
    .i5(\rfxs[5] [7]),
    .i6(\rfxs[6] [7]),
    .i7(\rfxs[7] [7]),
    .i8(\rfxs[8] [7]),
    .i9(\rfxs[9] [7]),
    .sel(i_rs1idx),
    .o(n95[7]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b8 (
    .i0(1'b0),
    .i1(\rfxs[1] [8]),
    .i10(\rfxs[10] [8]),
    .i11(\rfxs[11] [8]),
    .i12(\rfxs[12] [8]),
    .i13(\rfxs[13] [8]),
    .i14(\rfxs[14] [8]),
    .i15(\rfxs[15] [8]),
    .i16(\rfxs[16] [8]),
    .i17(\rfxs[17] [8]),
    .i18(\rfxs[18] [8]),
    .i19(\rfxs[19] [8]),
    .i2(\rfxs[2] [8]),
    .i20(\rfxs[20] [8]),
    .i21(\rfxs[21] [8]),
    .i22(\rfxs[22] [8]),
    .i23(\rfxs[23] [8]),
    .i24(\rfxs[24] [8]),
    .i25(\rfxs[25] [8]),
    .i26(\rfxs[26] [8]),
    .i27(\rfxs[27] [8]),
    .i28(\rfxs[28] [8]),
    .i29(\rfxs[29] [8]),
    .i3(\rfxs[3] [8]),
    .i30(\rfxs[30] [8]),
    .i31(\rfxs[31] [8]),
    .i4(\rfxs[4] [8]),
    .i5(\rfxs[5] [8]),
    .i6(\rfxs[6] [8]),
    .i7(\rfxs[7] [8]),
    .i8(\rfxs[8] [8]),
    .i9(\rfxs[9] [8]),
    .sel(i_rs1idx),
    .o(n95[8]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux31_b9 (
    .i0(1'b0),
    .i1(\rfxs[1] [9]),
    .i10(\rfxs[10] [9]),
    .i11(\rfxs[11] [9]),
    .i12(\rfxs[12] [9]),
    .i13(\rfxs[13] [9]),
    .i14(\rfxs[14] [9]),
    .i15(\rfxs[15] [9]),
    .i16(\rfxs[16] [9]),
    .i17(\rfxs[17] [9]),
    .i18(\rfxs[18] [9]),
    .i19(\rfxs[19] [9]),
    .i2(\rfxs[2] [9]),
    .i20(\rfxs[20] [9]),
    .i21(\rfxs[21] [9]),
    .i22(\rfxs[22] [9]),
    .i23(\rfxs[23] [9]),
    .i24(\rfxs[24] [9]),
    .i25(\rfxs[25] [9]),
    .i26(\rfxs[26] [9]),
    .i27(\rfxs[27] [9]),
    .i28(\rfxs[28] [9]),
    .i29(\rfxs[29] [9]),
    .i3(\rfxs[3] [9]),
    .i30(\rfxs[30] [9]),
    .i31(\rfxs[31] [9]),
    .i4(\rfxs[4] [9]),
    .i5(\rfxs[5] [9]),
    .i6(\rfxs[6] [9]),
    .i7(\rfxs[7] [9]),
    .i8(\rfxs[8] [9]),
    .i9(\rfxs[9] [9]),
    .sel(i_rs1idx),
    .o(n95[9]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b0 (
    .i0(n95[0]),
    .i1(i_rd_wdata[0]),
    .sel(n94),
    .o(n96[0]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b1 (
    .i0(n95[1]),
    .i1(i_rd_wdata[1]),
    .sel(n94),
    .o(n96[1]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b10 (
    .i0(n95[10]),
    .i1(i_rd_wdata[10]),
    .sel(n94),
    .o(n96[10]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b11 (
    .i0(n95[11]),
    .i1(i_rd_wdata[11]),
    .sel(n94),
    .o(n96[11]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b12 (
    .i0(n95[12]),
    .i1(i_rd_wdata[12]),
    .sel(n94),
    .o(n96[12]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b13 (
    .i0(n95[13]),
    .i1(i_rd_wdata[13]),
    .sel(n94),
    .o(n96[13]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b14 (
    .i0(n95[14]),
    .i1(i_rd_wdata[14]),
    .sel(n94),
    .o(n96[14]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b15 (
    .i0(n95[15]),
    .i1(i_rd_wdata[15]),
    .sel(n94),
    .o(n96[15]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b16 (
    .i0(n95[16]),
    .i1(i_rd_wdata[16]),
    .sel(n94),
    .o(n96[16]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b17 (
    .i0(n95[17]),
    .i1(i_rd_wdata[17]),
    .sel(n94),
    .o(n96[17]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b18 (
    .i0(n95[18]),
    .i1(i_rd_wdata[18]),
    .sel(n94),
    .o(n96[18]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b19 (
    .i0(n95[19]),
    .i1(i_rd_wdata[19]),
    .sel(n94),
    .o(n96[19]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b2 (
    .i0(n95[2]),
    .i1(i_rd_wdata[2]),
    .sel(n94),
    .o(n96[2]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b20 (
    .i0(n95[20]),
    .i1(i_rd_wdata[20]),
    .sel(n94),
    .o(n96[20]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b21 (
    .i0(n95[21]),
    .i1(i_rd_wdata[21]),
    .sel(n94),
    .o(n96[21]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b22 (
    .i0(n95[22]),
    .i1(i_rd_wdata[22]),
    .sel(n94),
    .o(n96[22]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b23 (
    .i0(n95[23]),
    .i1(i_rd_wdata[23]),
    .sel(n94),
    .o(n96[23]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b24 (
    .i0(n95[24]),
    .i1(i_rd_wdata[24]),
    .sel(n94),
    .o(n96[24]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b25 (
    .i0(n95[25]),
    .i1(i_rd_wdata[25]),
    .sel(n94),
    .o(n96[25]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b26 (
    .i0(n95[26]),
    .i1(i_rd_wdata[26]),
    .sel(n94),
    .o(n96[26]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b27 (
    .i0(n95[27]),
    .i1(i_rd_wdata[27]),
    .sel(n94),
    .o(n96[27]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b28 (
    .i0(n95[28]),
    .i1(i_rd_wdata[28]),
    .sel(n94),
    .o(n96[28]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b29 (
    .i0(n95[29]),
    .i1(i_rd_wdata[29]),
    .sel(n94),
    .o(n96[29]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b3 (
    .i0(n95[3]),
    .i1(i_rd_wdata[3]),
    .sel(n94),
    .o(n96[3]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b30 (
    .i0(n95[30]),
    .i1(i_rd_wdata[30]),
    .sel(n94),
    .o(n96[30]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b31 (
    .i0(n95[31]),
    .i1(i_rd_wdata[31]),
    .sel(n94),
    .o(n96[31]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b4 (
    .i0(n95[4]),
    .i1(i_rd_wdata[4]),
    .sel(n94),
    .o(n96[4]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b5 (
    .i0(n95[5]),
    .i1(i_rd_wdata[5]),
    .sel(n94),
    .o(n96[5]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b6 (
    .i0(n95[6]),
    .i1(i_rd_wdata[6]),
    .sel(n94),
    .o(n96[6]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b7 (
    .i0(n95[7]),
    .i1(i_rd_wdata[7]),
    .sel(n94),
    .o(n96[7]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b8 (
    .i0(n95[8]),
    .i1(i_rd_wdata[8]),
    .sel(n94),
    .o(n96[8]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux32_b9 (
    .i0(n95[9]),
    .i1(i_rd_wdata[9]),
    .sel(n94),
    .o(n96[9]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b0 (
    .i0(1'b0),
    .i1(n96[0]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[0]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b1 (
    .i0(1'b0),
    .i1(n96[1]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[1]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b10 (
    .i0(1'b0),
    .i1(n96[10]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[10]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b11 (
    .i0(1'b0),
    .i1(n96[11]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[11]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b12 (
    .i0(1'b0),
    .i1(n96[12]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[12]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b13 (
    .i0(1'b0),
    .i1(n96[13]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[13]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b14 (
    .i0(1'b0),
    .i1(n96[14]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[14]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b15 (
    .i0(1'b0),
    .i1(n96[15]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[15]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b16 (
    .i0(1'b0),
    .i1(n96[16]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[16]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b17 (
    .i0(1'b0),
    .i1(n96[17]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[17]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b18 (
    .i0(1'b0),
    .i1(n96[18]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[18]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b19 (
    .i0(1'b0),
    .i1(n96[19]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[19]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b2 (
    .i0(1'b0),
    .i1(n96[2]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[2]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b20 (
    .i0(1'b0),
    .i1(n96[20]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[20]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b21 (
    .i0(1'b0),
    .i1(n96[21]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[21]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b22 (
    .i0(1'b0),
    .i1(n96[22]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[22]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b23 (
    .i0(1'b0),
    .i1(n96[23]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[23]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b24 (
    .i0(1'b0),
    .i1(n96[24]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[24]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b25 (
    .i0(1'b0),
    .i1(n96[25]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[25]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b26 (
    .i0(1'b0),
    .i1(n96[26]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[26]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b27 (
    .i0(1'b0),
    .i1(n96[27]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[27]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b28 (
    .i0(1'b0),
    .i1(n96[28]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[28]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b29 (
    .i0(1'b0),
    .i1(n96[29]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[29]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b3 (
    .i0(1'b0),
    .i1(n96[3]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[3]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b30 (
    .i0(1'b0),
    .i1(n96[30]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[30]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b31 (
    .i0(1'b0),
    .i1(n96[31]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[31]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b4 (
    .i0(1'b0),
    .i1(n96[4]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[4]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b5 (
    .i0(1'b0),
    .i1(n96[5]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[5]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b6 (
    .i0(1'b0),
    .i1(n96[6]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[6]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b7 (
    .i0(1'b0),
    .i1(n96[7]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[7]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b8 (
    .i0(1'b0),
    .i1(n96[8]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[8]));  // ../RTL/core/regfile.v(46)
  binary_mux_s1_w1 mux33_b9 (
    .i0(1'b0),
    .i1(n96[9]),
    .sel(i_rs1ren),
    .o(o_rs1_rdata[9]));  // ../RTL/core/regfile.v(46)
  binary_mux_s5_w1 mux34_b0 (
    .i0(1'b0),
    .i1(\rfxs[1] [0]),
    .i10(\rfxs[10] [0]),
    .i11(\rfxs[11] [0]),
    .i12(\rfxs[12] [0]),
    .i13(\rfxs[13] [0]),
    .i14(\rfxs[14] [0]),
    .i15(\rfxs[15] [0]),
    .i16(\rfxs[16] [0]),
    .i17(\rfxs[17] [0]),
    .i18(\rfxs[18] [0]),
    .i19(\rfxs[19] [0]),
    .i2(\rfxs[2] [0]),
    .i20(\rfxs[20] [0]),
    .i21(\rfxs[21] [0]),
    .i22(\rfxs[22] [0]),
    .i23(\rfxs[23] [0]),
    .i24(\rfxs[24] [0]),
    .i25(\rfxs[25] [0]),
    .i26(\rfxs[26] [0]),
    .i27(\rfxs[27] [0]),
    .i28(\rfxs[28] [0]),
    .i29(\rfxs[29] [0]),
    .i3(\rfxs[3] [0]),
    .i30(\rfxs[30] [0]),
    .i31(\rfxs[31] [0]),
    .i4(\rfxs[4] [0]),
    .i5(\rfxs[5] [0]),
    .i6(\rfxs[6] [0]),
    .i7(\rfxs[7] [0]),
    .i8(\rfxs[8] [0]),
    .i9(\rfxs[9] [0]),
    .sel(i_rs2idx),
    .o(n99[0]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b1 (
    .i0(1'b0),
    .i1(\rfxs[1] [1]),
    .i10(\rfxs[10] [1]),
    .i11(\rfxs[11] [1]),
    .i12(\rfxs[12] [1]),
    .i13(\rfxs[13] [1]),
    .i14(\rfxs[14] [1]),
    .i15(\rfxs[15] [1]),
    .i16(\rfxs[16] [1]),
    .i17(\rfxs[17] [1]),
    .i18(\rfxs[18] [1]),
    .i19(\rfxs[19] [1]),
    .i2(\rfxs[2] [1]),
    .i20(\rfxs[20] [1]),
    .i21(\rfxs[21] [1]),
    .i22(\rfxs[22] [1]),
    .i23(\rfxs[23] [1]),
    .i24(\rfxs[24] [1]),
    .i25(\rfxs[25] [1]),
    .i26(\rfxs[26] [1]),
    .i27(\rfxs[27] [1]),
    .i28(\rfxs[28] [1]),
    .i29(\rfxs[29] [1]),
    .i3(\rfxs[3] [1]),
    .i30(\rfxs[30] [1]),
    .i31(\rfxs[31] [1]),
    .i4(\rfxs[4] [1]),
    .i5(\rfxs[5] [1]),
    .i6(\rfxs[6] [1]),
    .i7(\rfxs[7] [1]),
    .i8(\rfxs[8] [1]),
    .i9(\rfxs[9] [1]),
    .sel(i_rs2idx),
    .o(n99[1]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b10 (
    .i0(1'b0),
    .i1(\rfxs[1] [10]),
    .i10(\rfxs[10] [10]),
    .i11(\rfxs[11] [10]),
    .i12(\rfxs[12] [10]),
    .i13(\rfxs[13] [10]),
    .i14(\rfxs[14] [10]),
    .i15(\rfxs[15] [10]),
    .i16(\rfxs[16] [10]),
    .i17(\rfxs[17] [10]),
    .i18(\rfxs[18] [10]),
    .i19(\rfxs[19] [10]),
    .i2(\rfxs[2] [10]),
    .i20(\rfxs[20] [10]),
    .i21(\rfxs[21] [10]),
    .i22(\rfxs[22] [10]),
    .i23(\rfxs[23] [10]),
    .i24(\rfxs[24] [10]),
    .i25(\rfxs[25] [10]),
    .i26(\rfxs[26] [10]),
    .i27(\rfxs[27] [10]),
    .i28(\rfxs[28] [10]),
    .i29(\rfxs[29] [10]),
    .i3(\rfxs[3] [10]),
    .i30(\rfxs[30] [10]),
    .i31(\rfxs[31] [10]),
    .i4(\rfxs[4] [10]),
    .i5(\rfxs[5] [10]),
    .i6(\rfxs[6] [10]),
    .i7(\rfxs[7] [10]),
    .i8(\rfxs[8] [10]),
    .i9(\rfxs[9] [10]),
    .sel(i_rs2idx),
    .o(n99[10]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b11 (
    .i0(1'b0),
    .i1(\rfxs[1] [11]),
    .i10(\rfxs[10] [11]),
    .i11(\rfxs[11] [11]),
    .i12(\rfxs[12] [11]),
    .i13(\rfxs[13] [11]),
    .i14(\rfxs[14] [11]),
    .i15(\rfxs[15] [11]),
    .i16(\rfxs[16] [11]),
    .i17(\rfxs[17] [11]),
    .i18(\rfxs[18] [11]),
    .i19(\rfxs[19] [11]),
    .i2(\rfxs[2] [11]),
    .i20(\rfxs[20] [11]),
    .i21(\rfxs[21] [11]),
    .i22(\rfxs[22] [11]),
    .i23(\rfxs[23] [11]),
    .i24(\rfxs[24] [11]),
    .i25(\rfxs[25] [11]),
    .i26(\rfxs[26] [11]),
    .i27(\rfxs[27] [11]),
    .i28(\rfxs[28] [11]),
    .i29(\rfxs[29] [11]),
    .i3(\rfxs[3] [11]),
    .i30(\rfxs[30] [11]),
    .i31(\rfxs[31] [11]),
    .i4(\rfxs[4] [11]),
    .i5(\rfxs[5] [11]),
    .i6(\rfxs[6] [11]),
    .i7(\rfxs[7] [11]),
    .i8(\rfxs[8] [11]),
    .i9(\rfxs[9] [11]),
    .sel(i_rs2idx),
    .o(n99[11]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b12 (
    .i0(1'b0),
    .i1(\rfxs[1] [12]),
    .i10(\rfxs[10] [12]),
    .i11(\rfxs[11] [12]),
    .i12(\rfxs[12] [12]),
    .i13(\rfxs[13] [12]),
    .i14(\rfxs[14] [12]),
    .i15(\rfxs[15] [12]),
    .i16(\rfxs[16] [12]),
    .i17(\rfxs[17] [12]),
    .i18(\rfxs[18] [12]),
    .i19(\rfxs[19] [12]),
    .i2(\rfxs[2] [12]),
    .i20(\rfxs[20] [12]),
    .i21(\rfxs[21] [12]),
    .i22(\rfxs[22] [12]),
    .i23(\rfxs[23] [12]),
    .i24(\rfxs[24] [12]),
    .i25(\rfxs[25] [12]),
    .i26(\rfxs[26] [12]),
    .i27(\rfxs[27] [12]),
    .i28(\rfxs[28] [12]),
    .i29(\rfxs[29] [12]),
    .i3(\rfxs[3] [12]),
    .i30(\rfxs[30] [12]),
    .i31(\rfxs[31] [12]),
    .i4(\rfxs[4] [12]),
    .i5(\rfxs[5] [12]),
    .i6(\rfxs[6] [12]),
    .i7(\rfxs[7] [12]),
    .i8(\rfxs[8] [12]),
    .i9(\rfxs[9] [12]),
    .sel(i_rs2idx),
    .o(n99[12]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b13 (
    .i0(1'b0),
    .i1(\rfxs[1] [13]),
    .i10(\rfxs[10] [13]),
    .i11(\rfxs[11] [13]),
    .i12(\rfxs[12] [13]),
    .i13(\rfxs[13] [13]),
    .i14(\rfxs[14] [13]),
    .i15(\rfxs[15] [13]),
    .i16(\rfxs[16] [13]),
    .i17(\rfxs[17] [13]),
    .i18(\rfxs[18] [13]),
    .i19(\rfxs[19] [13]),
    .i2(\rfxs[2] [13]),
    .i20(\rfxs[20] [13]),
    .i21(\rfxs[21] [13]),
    .i22(\rfxs[22] [13]),
    .i23(\rfxs[23] [13]),
    .i24(\rfxs[24] [13]),
    .i25(\rfxs[25] [13]),
    .i26(\rfxs[26] [13]),
    .i27(\rfxs[27] [13]),
    .i28(\rfxs[28] [13]),
    .i29(\rfxs[29] [13]),
    .i3(\rfxs[3] [13]),
    .i30(\rfxs[30] [13]),
    .i31(\rfxs[31] [13]),
    .i4(\rfxs[4] [13]),
    .i5(\rfxs[5] [13]),
    .i6(\rfxs[6] [13]),
    .i7(\rfxs[7] [13]),
    .i8(\rfxs[8] [13]),
    .i9(\rfxs[9] [13]),
    .sel(i_rs2idx),
    .o(n99[13]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b14 (
    .i0(1'b0),
    .i1(\rfxs[1] [14]),
    .i10(\rfxs[10] [14]),
    .i11(\rfxs[11] [14]),
    .i12(\rfxs[12] [14]),
    .i13(\rfxs[13] [14]),
    .i14(\rfxs[14] [14]),
    .i15(\rfxs[15] [14]),
    .i16(\rfxs[16] [14]),
    .i17(\rfxs[17] [14]),
    .i18(\rfxs[18] [14]),
    .i19(\rfxs[19] [14]),
    .i2(\rfxs[2] [14]),
    .i20(\rfxs[20] [14]),
    .i21(\rfxs[21] [14]),
    .i22(\rfxs[22] [14]),
    .i23(\rfxs[23] [14]),
    .i24(\rfxs[24] [14]),
    .i25(\rfxs[25] [14]),
    .i26(\rfxs[26] [14]),
    .i27(\rfxs[27] [14]),
    .i28(\rfxs[28] [14]),
    .i29(\rfxs[29] [14]),
    .i3(\rfxs[3] [14]),
    .i30(\rfxs[30] [14]),
    .i31(\rfxs[31] [14]),
    .i4(\rfxs[4] [14]),
    .i5(\rfxs[5] [14]),
    .i6(\rfxs[6] [14]),
    .i7(\rfxs[7] [14]),
    .i8(\rfxs[8] [14]),
    .i9(\rfxs[9] [14]),
    .sel(i_rs2idx),
    .o(n99[14]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b15 (
    .i0(1'b0),
    .i1(\rfxs[1] [15]),
    .i10(\rfxs[10] [15]),
    .i11(\rfxs[11] [15]),
    .i12(\rfxs[12] [15]),
    .i13(\rfxs[13] [15]),
    .i14(\rfxs[14] [15]),
    .i15(\rfxs[15] [15]),
    .i16(\rfxs[16] [15]),
    .i17(\rfxs[17] [15]),
    .i18(\rfxs[18] [15]),
    .i19(\rfxs[19] [15]),
    .i2(\rfxs[2] [15]),
    .i20(\rfxs[20] [15]),
    .i21(\rfxs[21] [15]),
    .i22(\rfxs[22] [15]),
    .i23(\rfxs[23] [15]),
    .i24(\rfxs[24] [15]),
    .i25(\rfxs[25] [15]),
    .i26(\rfxs[26] [15]),
    .i27(\rfxs[27] [15]),
    .i28(\rfxs[28] [15]),
    .i29(\rfxs[29] [15]),
    .i3(\rfxs[3] [15]),
    .i30(\rfxs[30] [15]),
    .i31(\rfxs[31] [15]),
    .i4(\rfxs[4] [15]),
    .i5(\rfxs[5] [15]),
    .i6(\rfxs[6] [15]),
    .i7(\rfxs[7] [15]),
    .i8(\rfxs[8] [15]),
    .i9(\rfxs[9] [15]),
    .sel(i_rs2idx),
    .o(n99[15]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b16 (
    .i0(1'b0),
    .i1(\rfxs[1] [16]),
    .i10(\rfxs[10] [16]),
    .i11(\rfxs[11] [16]),
    .i12(\rfxs[12] [16]),
    .i13(\rfxs[13] [16]),
    .i14(\rfxs[14] [16]),
    .i15(\rfxs[15] [16]),
    .i16(\rfxs[16] [16]),
    .i17(\rfxs[17] [16]),
    .i18(\rfxs[18] [16]),
    .i19(\rfxs[19] [16]),
    .i2(\rfxs[2] [16]),
    .i20(\rfxs[20] [16]),
    .i21(\rfxs[21] [16]),
    .i22(\rfxs[22] [16]),
    .i23(\rfxs[23] [16]),
    .i24(\rfxs[24] [16]),
    .i25(\rfxs[25] [16]),
    .i26(\rfxs[26] [16]),
    .i27(\rfxs[27] [16]),
    .i28(\rfxs[28] [16]),
    .i29(\rfxs[29] [16]),
    .i3(\rfxs[3] [16]),
    .i30(\rfxs[30] [16]),
    .i31(\rfxs[31] [16]),
    .i4(\rfxs[4] [16]),
    .i5(\rfxs[5] [16]),
    .i6(\rfxs[6] [16]),
    .i7(\rfxs[7] [16]),
    .i8(\rfxs[8] [16]),
    .i9(\rfxs[9] [16]),
    .sel(i_rs2idx),
    .o(n99[16]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b17 (
    .i0(1'b0),
    .i1(\rfxs[1] [17]),
    .i10(\rfxs[10] [17]),
    .i11(\rfxs[11] [17]),
    .i12(\rfxs[12] [17]),
    .i13(\rfxs[13] [17]),
    .i14(\rfxs[14] [17]),
    .i15(\rfxs[15] [17]),
    .i16(\rfxs[16] [17]),
    .i17(\rfxs[17] [17]),
    .i18(\rfxs[18] [17]),
    .i19(\rfxs[19] [17]),
    .i2(\rfxs[2] [17]),
    .i20(\rfxs[20] [17]),
    .i21(\rfxs[21] [17]),
    .i22(\rfxs[22] [17]),
    .i23(\rfxs[23] [17]),
    .i24(\rfxs[24] [17]),
    .i25(\rfxs[25] [17]),
    .i26(\rfxs[26] [17]),
    .i27(\rfxs[27] [17]),
    .i28(\rfxs[28] [17]),
    .i29(\rfxs[29] [17]),
    .i3(\rfxs[3] [17]),
    .i30(\rfxs[30] [17]),
    .i31(\rfxs[31] [17]),
    .i4(\rfxs[4] [17]),
    .i5(\rfxs[5] [17]),
    .i6(\rfxs[6] [17]),
    .i7(\rfxs[7] [17]),
    .i8(\rfxs[8] [17]),
    .i9(\rfxs[9] [17]),
    .sel(i_rs2idx),
    .o(n99[17]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b18 (
    .i0(1'b0),
    .i1(\rfxs[1] [18]),
    .i10(\rfxs[10] [18]),
    .i11(\rfxs[11] [18]),
    .i12(\rfxs[12] [18]),
    .i13(\rfxs[13] [18]),
    .i14(\rfxs[14] [18]),
    .i15(\rfxs[15] [18]),
    .i16(\rfxs[16] [18]),
    .i17(\rfxs[17] [18]),
    .i18(\rfxs[18] [18]),
    .i19(\rfxs[19] [18]),
    .i2(\rfxs[2] [18]),
    .i20(\rfxs[20] [18]),
    .i21(\rfxs[21] [18]),
    .i22(\rfxs[22] [18]),
    .i23(\rfxs[23] [18]),
    .i24(\rfxs[24] [18]),
    .i25(\rfxs[25] [18]),
    .i26(\rfxs[26] [18]),
    .i27(\rfxs[27] [18]),
    .i28(\rfxs[28] [18]),
    .i29(\rfxs[29] [18]),
    .i3(\rfxs[3] [18]),
    .i30(\rfxs[30] [18]),
    .i31(\rfxs[31] [18]),
    .i4(\rfxs[4] [18]),
    .i5(\rfxs[5] [18]),
    .i6(\rfxs[6] [18]),
    .i7(\rfxs[7] [18]),
    .i8(\rfxs[8] [18]),
    .i9(\rfxs[9] [18]),
    .sel(i_rs2idx),
    .o(n99[18]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b19 (
    .i0(1'b0),
    .i1(\rfxs[1] [19]),
    .i10(\rfxs[10] [19]),
    .i11(\rfxs[11] [19]),
    .i12(\rfxs[12] [19]),
    .i13(\rfxs[13] [19]),
    .i14(\rfxs[14] [19]),
    .i15(\rfxs[15] [19]),
    .i16(\rfxs[16] [19]),
    .i17(\rfxs[17] [19]),
    .i18(\rfxs[18] [19]),
    .i19(\rfxs[19] [19]),
    .i2(\rfxs[2] [19]),
    .i20(\rfxs[20] [19]),
    .i21(\rfxs[21] [19]),
    .i22(\rfxs[22] [19]),
    .i23(\rfxs[23] [19]),
    .i24(\rfxs[24] [19]),
    .i25(\rfxs[25] [19]),
    .i26(\rfxs[26] [19]),
    .i27(\rfxs[27] [19]),
    .i28(\rfxs[28] [19]),
    .i29(\rfxs[29] [19]),
    .i3(\rfxs[3] [19]),
    .i30(\rfxs[30] [19]),
    .i31(\rfxs[31] [19]),
    .i4(\rfxs[4] [19]),
    .i5(\rfxs[5] [19]),
    .i6(\rfxs[6] [19]),
    .i7(\rfxs[7] [19]),
    .i8(\rfxs[8] [19]),
    .i9(\rfxs[9] [19]),
    .sel(i_rs2idx),
    .o(n99[19]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b2 (
    .i0(1'b0),
    .i1(\rfxs[1] [2]),
    .i10(\rfxs[10] [2]),
    .i11(\rfxs[11] [2]),
    .i12(\rfxs[12] [2]),
    .i13(\rfxs[13] [2]),
    .i14(\rfxs[14] [2]),
    .i15(\rfxs[15] [2]),
    .i16(\rfxs[16] [2]),
    .i17(\rfxs[17] [2]),
    .i18(\rfxs[18] [2]),
    .i19(\rfxs[19] [2]),
    .i2(\rfxs[2] [2]),
    .i20(\rfxs[20] [2]),
    .i21(\rfxs[21] [2]),
    .i22(\rfxs[22] [2]),
    .i23(\rfxs[23] [2]),
    .i24(\rfxs[24] [2]),
    .i25(\rfxs[25] [2]),
    .i26(\rfxs[26] [2]),
    .i27(\rfxs[27] [2]),
    .i28(\rfxs[28] [2]),
    .i29(\rfxs[29] [2]),
    .i3(\rfxs[3] [2]),
    .i30(\rfxs[30] [2]),
    .i31(\rfxs[31] [2]),
    .i4(\rfxs[4] [2]),
    .i5(\rfxs[5] [2]),
    .i6(\rfxs[6] [2]),
    .i7(\rfxs[7] [2]),
    .i8(\rfxs[8] [2]),
    .i9(\rfxs[9] [2]),
    .sel(i_rs2idx),
    .o(n99[2]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b20 (
    .i0(1'b0),
    .i1(\rfxs[1] [20]),
    .i10(\rfxs[10] [20]),
    .i11(\rfxs[11] [20]),
    .i12(\rfxs[12] [20]),
    .i13(\rfxs[13] [20]),
    .i14(\rfxs[14] [20]),
    .i15(\rfxs[15] [20]),
    .i16(\rfxs[16] [20]),
    .i17(\rfxs[17] [20]),
    .i18(\rfxs[18] [20]),
    .i19(\rfxs[19] [20]),
    .i2(\rfxs[2] [20]),
    .i20(\rfxs[20] [20]),
    .i21(\rfxs[21] [20]),
    .i22(\rfxs[22] [20]),
    .i23(\rfxs[23] [20]),
    .i24(\rfxs[24] [20]),
    .i25(\rfxs[25] [20]),
    .i26(\rfxs[26] [20]),
    .i27(\rfxs[27] [20]),
    .i28(\rfxs[28] [20]),
    .i29(\rfxs[29] [20]),
    .i3(\rfxs[3] [20]),
    .i30(\rfxs[30] [20]),
    .i31(\rfxs[31] [20]),
    .i4(\rfxs[4] [20]),
    .i5(\rfxs[5] [20]),
    .i6(\rfxs[6] [20]),
    .i7(\rfxs[7] [20]),
    .i8(\rfxs[8] [20]),
    .i9(\rfxs[9] [20]),
    .sel(i_rs2idx),
    .o(n99[20]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b21 (
    .i0(1'b0),
    .i1(\rfxs[1] [21]),
    .i10(\rfxs[10] [21]),
    .i11(\rfxs[11] [21]),
    .i12(\rfxs[12] [21]),
    .i13(\rfxs[13] [21]),
    .i14(\rfxs[14] [21]),
    .i15(\rfxs[15] [21]),
    .i16(\rfxs[16] [21]),
    .i17(\rfxs[17] [21]),
    .i18(\rfxs[18] [21]),
    .i19(\rfxs[19] [21]),
    .i2(\rfxs[2] [21]),
    .i20(\rfxs[20] [21]),
    .i21(\rfxs[21] [21]),
    .i22(\rfxs[22] [21]),
    .i23(\rfxs[23] [21]),
    .i24(\rfxs[24] [21]),
    .i25(\rfxs[25] [21]),
    .i26(\rfxs[26] [21]),
    .i27(\rfxs[27] [21]),
    .i28(\rfxs[28] [21]),
    .i29(\rfxs[29] [21]),
    .i3(\rfxs[3] [21]),
    .i30(\rfxs[30] [21]),
    .i31(\rfxs[31] [21]),
    .i4(\rfxs[4] [21]),
    .i5(\rfxs[5] [21]),
    .i6(\rfxs[6] [21]),
    .i7(\rfxs[7] [21]),
    .i8(\rfxs[8] [21]),
    .i9(\rfxs[9] [21]),
    .sel(i_rs2idx),
    .o(n99[21]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b22 (
    .i0(1'b0),
    .i1(\rfxs[1] [22]),
    .i10(\rfxs[10] [22]),
    .i11(\rfxs[11] [22]),
    .i12(\rfxs[12] [22]),
    .i13(\rfxs[13] [22]),
    .i14(\rfxs[14] [22]),
    .i15(\rfxs[15] [22]),
    .i16(\rfxs[16] [22]),
    .i17(\rfxs[17] [22]),
    .i18(\rfxs[18] [22]),
    .i19(\rfxs[19] [22]),
    .i2(\rfxs[2] [22]),
    .i20(\rfxs[20] [22]),
    .i21(\rfxs[21] [22]),
    .i22(\rfxs[22] [22]),
    .i23(\rfxs[23] [22]),
    .i24(\rfxs[24] [22]),
    .i25(\rfxs[25] [22]),
    .i26(\rfxs[26] [22]),
    .i27(\rfxs[27] [22]),
    .i28(\rfxs[28] [22]),
    .i29(\rfxs[29] [22]),
    .i3(\rfxs[3] [22]),
    .i30(\rfxs[30] [22]),
    .i31(\rfxs[31] [22]),
    .i4(\rfxs[4] [22]),
    .i5(\rfxs[5] [22]),
    .i6(\rfxs[6] [22]),
    .i7(\rfxs[7] [22]),
    .i8(\rfxs[8] [22]),
    .i9(\rfxs[9] [22]),
    .sel(i_rs2idx),
    .o(n99[22]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b23 (
    .i0(1'b0),
    .i1(\rfxs[1] [23]),
    .i10(\rfxs[10] [23]),
    .i11(\rfxs[11] [23]),
    .i12(\rfxs[12] [23]),
    .i13(\rfxs[13] [23]),
    .i14(\rfxs[14] [23]),
    .i15(\rfxs[15] [23]),
    .i16(\rfxs[16] [23]),
    .i17(\rfxs[17] [23]),
    .i18(\rfxs[18] [23]),
    .i19(\rfxs[19] [23]),
    .i2(\rfxs[2] [23]),
    .i20(\rfxs[20] [23]),
    .i21(\rfxs[21] [23]),
    .i22(\rfxs[22] [23]),
    .i23(\rfxs[23] [23]),
    .i24(\rfxs[24] [23]),
    .i25(\rfxs[25] [23]),
    .i26(\rfxs[26] [23]),
    .i27(\rfxs[27] [23]),
    .i28(\rfxs[28] [23]),
    .i29(\rfxs[29] [23]),
    .i3(\rfxs[3] [23]),
    .i30(\rfxs[30] [23]),
    .i31(\rfxs[31] [23]),
    .i4(\rfxs[4] [23]),
    .i5(\rfxs[5] [23]),
    .i6(\rfxs[6] [23]),
    .i7(\rfxs[7] [23]),
    .i8(\rfxs[8] [23]),
    .i9(\rfxs[9] [23]),
    .sel(i_rs2idx),
    .o(n99[23]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b24 (
    .i0(1'b0),
    .i1(\rfxs[1] [24]),
    .i10(\rfxs[10] [24]),
    .i11(\rfxs[11] [24]),
    .i12(\rfxs[12] [24]),
    .i13(\rfxs[13] [24]),
    .i14(\rfxs[14] [24]),
    .i15(\rfxs[15] [24]),
    .i16(\rfxs[16] [24]),
    .i17(\rfxs[17] [24]),
    .i18(\rfxs[18] [24]),
    .i19(\rfxs[19] [24]),
    .i2(\rfxs[2] [24]),
    .i20(\rfxs[20] [24]),
    .i21(\rfxs[21] [24]),
    .i22(\rfxs[22] [24]),
    .i23(\rfxs[23] [24]),
    .i24(\rfxs[24] [24]),
    .i25(\rfxs[25] [24]),
    .i26(\rfxs[26] [24]),
    .i27(\rfxs[27] [24]),
    .i28(\rfxs[28] [24]),
    .i29(\rfxs[29] [24]),
    .i3(\rfxs[3] [24]),
    .i30(\rfxs[30] [24]),
    .i31(\rfxs[31] [24]),
    .i4(\rfxs[4] [24]),
    .i5(\rfxs[5] [24]),
    .i6(\rfxs[6] [24]),
    .i7(\rfxs[7] [24]),
    .i8(\rfxs[8] [24]),
    .i9(\rfxs[9] [24]),
    .sel(i_rs2idx),
    .o(n99[24]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b25 (
    .i0(1'b0),
    .i1(\rfxs[1] [25]),
    .i10(\rfxs[10] [25]),
    .i11(\rfxs[11] [25]),
    .i12(\rfxs[12] [25]),
    .i13(\rfxs[13] [25]),
    .i14(\rfxs[14] [25]),
    .i15(\rfxs[15] [25]),
    .i16(\rfxs[16] [25]),
    .i17(\rfxs[17] [25]),
    .i18(\rfxs[18] [25]),
    .i19(\rfxs[19] [25]),
    .i2(\rfxs[2] [25]),
    .i20(\rfxs[20] [25]),
    .i21(\rfxs[21] [25]),
    .i22(\rfxs[22] [25]),
    .i23(\rfxs[23] [25]),
    .i24(\rfxs[24] [25]),
    .i25(\rfxs[25] [25]),
    .i26(\rfxs[26] [25]),
    .i27(\rfxs[27] [25]),
    .i28(\rfxs[28] [25]),
    .i29(\rfxs[29] [25]),
    .i3(\rfxs[3] [25]),
    .i30(\rfxs[30] [25]),
    .i31(\rfxs[31] [25]),
    .i4(\rfxs[4] [25]),
    .i5(\rfxs[5] [25]),
    .i6(\rfxs[6] [25]),
    .i7(\rfxs[7] [25]),
    .i8(\rfxs[8] [25]),
    .i9(\rfxs[9] [25]),
    .sel(i_rs2idx),
    .o(n99[25]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b26 (
    .i0(1'b0),
    .i1(\rfxs[1] [26]),
    .i10(\rfxs[10] [26]),
    .i11(\rfxs[11] [26]),
    .i12(\rfxs[12] [26]),
    .i13(\rfxs[13] [26]),
    .i14(\rfxs[14] [26]),
    .i15(\rfxs[15] [26]),
    .i16(\rfxs[16] [26]),
    .i17(\rfxs[17] [26]),
    .i18(\rfxs[18] [26]),
    .i19(\rfxs[19] [26]),
    .i2(\rfxs[2] [26]),
    .i20(\rfxs[20] [26]),
    .i21(\rfxs[21] [26]),
    .i22(\rfxs[22] [26]),
    .i23(\rfxs[23] [26]),
    .i24(\rfxs[24] [26]),
    .i25(\rfxs[25] [26]),
    .i26(\rfxs[26] [26]),
    .i27(\rfxs[27] [26]),
    .i28(\rfxs[28] [26]),
    .i29(\rfxs[29] [26]),
    .i3(\rfxs[3] [26]),
    .i30(\rfxs[30] [26]),
    .i31(\rfxs[31] [26]),
    .i4(\rfxs[4] [26]),
    .i5(\rfxs[5] [26]),
    .i6(\rfxs[6] [26]),
    .i7(\rfxs[7] [26]),
    .i8(\rfxs[8] [26]),
    .i9(\rfxs[9] [26]),
    .sel(i_rs2idx),
    .o(n99[26]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b27 (
    .i0(1'b0),
    .i1(\rfxs[1] [27]),
    .i10(\rfxs[10] [27]),
    .i11(\rfxs[11] [27]),
    .i12(\rfxs[12] [27]),
    .i13(\rfxs[13] [27]),
    .i14(\rfxs[14] [27]),
    .i15(\rfxs[15] [27]),
    .i16(\rfxs[16] [27]),
    .i17(\rfxs[17] [27]),
    .i18(\rfxs[18] [27]),
    .i19(\rfxs[19] [27]),
    .i2(\rfxs[2] [27]),
    .i20(\rfxs[20] [27]),
    .i21(\rfxs[21] [27]),
    .i22(\rfxs[22] [27]),
    .i23(\rfxs[23] [27]),
    .i24(\rfxs[24] [27]),
    .i25(\rfxs[25] [27]),
    .i26(\rfxs[26] [27]),
    .i27(\rfxs[27] [27]),
    .i28(\rfxs[28] [27]),
    .i29(\rfxs[29] [27]),
    .i3(\rfxs[3] [27]),
    .i30(\rfxs[30] [27]),
    .i31(\rfxs[31] [27]),
    .i4(\rfxs[4] [27]),
    .i5(\rfxs[5] [27]),
    .i6(\rfxs[6] [27]),
    .i7(\rfxs[7] [27]),
    .i8(\rfxs[8] [27]),
    .i9(\rfxs[9] [27]),
    .sel(i_rs2idx),
    .o(n99[27]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b28 (
    .i0(1'b0),
    .i1(\rfxs[1] [28]),
    .i10(\rfxs[10] [28]),
    .i11(\rfxs[11] [28]),
    .i12(\rfxs[12] [28]),
    .i13(\rfxs[13] [28]),
    .i14(\rfxs[14] [28]),
    .i15(\rfxs[15] [28]),
    .i16(\rfxs[16] [28]),
    .i17(\rfxs[17] [28]),
    .i18(\rfxs[18] [28]),
    .i19(\rfxs[19] [28]),
    .i2(\rfxs[2] [28]),
    .i20(\rfxs[20] [28]),
    .i21(\rfxs[21] [28]),
    .i22(\rfxs[22] [28]),
    .i23(\rfxs[23] [28]),
    .i24(\rfxs[24] [28]),
    .i25(\rfxs[25] [28]),
    .i26(\rfxs[26] [28]),
    .i27(\rfxs[27] [28]),
    .i28(\rfxs[28] [28]),
    .i29(\rfxs[29] [28]),
    .i3(\rfxs[3] [28]),
    .i30(\rfxs[30] [28]),
    .i31(\rfxs[31] [28]),
    .i4(\rfxs[4] [28]),
    .i5(\rfxs[5] [28]),
    .i6(\rfxs[6] [28]),
    .i7(\rfxs[7] [28]),
    .i8(\rfxs[8] [28]),
    .i9(\rfxs[9] [28]),
    .sel(i_rs2idx),
    .o(n99[28]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b29 (
    .i0(1'b0),
    .i1(\rfxs[1] [29]),
    .i10(\rfxs[10] [29]),
    .i11(\rfxs[11] [29]),
    .i12(\rfxs[12] [29]),
    .i13(\rfxs[13] [29]),
    .i14(\rfxs[14] [29]),
    .i15(\rfxs[15] [29]),
    .i16(\rfxs[16] [29]),
    .i17(\rfxs[17] [29]),
    .i18(\rfxs[18] [29]),
    .i19(\rfxs[19] [29]),
    .i2(\rfxs[2] [29]),
    .i20(\rfxs[20] [29]),
    .i21(\rfxs[21] [29]),
    .i22(\rfxs[22] [29]),
    .i23(\rfxs[23] [29]),
    .i24(\rfxs[24] [29]),
    .i25(\rfxs[25] [29]),
    .i26(\rfxs[26] [29]),
    .i27(\rfxs[27] [29]),
    .i28(\rfxs[28] [29]),
    .i29(\rfxs[29] [29]),
    .i3(\rfxs[3] [29]),
    .i30(\rfxs[30] [29]),
    .i31(\rfxs[31] [29]),
    .i4(\rfxs[4] [29]),
    .i5(\rfxs[5] [29]),
    .i6(\rfxs[6] [29]),
    .i7(\rfxs[7] [29]),
    .i8(\rfxs[8] [29]),
    .i9(\rfxs[9] [29]),
    .sel(i_rs2idx),
    .o(n99[29]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b3 (
    .i0(1'b0),
    .i1(\rfxs[1] [3]),
    .i10(\rfxs[10] [3]),
    .i11(\rfxs[11] [3]),
    .i12(\rfxs[12] [3]),
    .i13(\rfxs[13] [3]),
    .i14(\rfxs[14] [3]),
    .i15(\rfxs[15] [3]),
    .i16(\rfxs[16] [3]),
    .i17(\rfxs[17] [3]),
    .i18(\rfxs[18] [3]),
    .i19(\rfxs[19] [3]),
    .i2(\rfxs[2] [3]),
    .i20(\rfxs[20] [3]),
    .i21(\rfxs[21] [3]),
    .i22(\rfxs[22] [3]),
    .i23(\rfxs[23] [3]),
    .i24(\rfxs[24] [3]),
    .i25(\rfxs[25] [3]),
    .i26(\rfxs[26] [3]),
    .i27(\rfxs[27] [3]),
    .i28(\rfxs[28] [3]),
    .i29(\rfxs[29] [3]),
    .i3(\rfxs[3] [3]),
    .i30(\rfxs[30] [3]),
    .i31(\rfxs[31] [3]),
    .i4(\rfxs[4] [3]),
    .i5(\rfxs[5] [3]),
    .i6(\rfxs[6] [3]),
    .i7(\rfxs[7] [3]),
    .i8(\rfxs[8] [3]),
    .i9(\rfxs[9] [3]),
    .sel(i_rs2idx),
    .o(n99[3]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b30 (
    .i0(1'b0),
    .i1(\rfxs[1] [30]),
    .i10(\rfxs[10] [30]),
    .i11(\rfxs[11] [30]),
    .i12(\rfxs[12] [30]),
    .i13(\rfxs[13] [30]),
    .i14(\rfxs[14] [30]),
    .i15(\rfxs[15] [30]),
    .i16(\rfxs[16] [30]),
    .i17(\rfxs[17] [30]),
    .i18(\rfxs[18] [30]),
    .i19(\rfxs[19] [30]),
    .i2(\rfxs[2] [30]),
    .i20(\rfxs[20] [30]),
    .i21(\rfxs[21] [30]),
    .i22(\rfxs[22] [30]),
    .i23(\rfxs[23] [30]),
    .i24(\rfxs[24] [30]),
    .i25(\rfxs[25] [30]),
    .i26(\rfxs[26] [30]),
    .i27(\rfxs[27] [30]),
    .i28(\rfxs[28] [30]),
    .i29(\rfxs[29] [30]),
    .i3(\rfxs[3] [30]),
    .i30(\rfxs[30] [30]),
    .i31(\rfxs[31] [30]),
    .i4(\rfxs[4] [30]),
    .i5(\rfxs[5] [30]),
    .i6(\rfxs[6] [30]),
    .i7(\rfxs[7] [30]),
    .i8(\rfxs[8] [30]),
    .i9(\rfxs[9] [30]),
    .sel(i_rs2idx),
    .o(n99[30]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b31 (
    .i0(1'b0),
    .i1(\rfxs[1] [31]),
    .i10(\rfxs[10] [31]),
    .i11(\rfxs[11] [31]),
    .i12(\rfxs[12] [31]),
    .i13(\rfxs[13] [31]),
    .i14(\rfxs[14] [31]),
    .i15(\rfxs[15] [31]),
    .i16(\rfxs[16] [31]),
    .i17(\rfxs[17] [31]),
    .i18(\rfxs[18] [31]),
    .i19(\rfxs[19] [31]),
    .i2(\rfxs[2] [31]),
    .i20(\rfxs[20] [31]),
    .i21(\rfxs[21] [31]),
    .i22(\rfxs[22] [31]),
    .i23(\rfxs[23] [31]),
    .i24(\rfxs[24] [31]),
    .i25(\rfxs[25] [31]),
    .i26(\rfxs[26] [31]),
    .i27(\rfxs[27] [31]),
    .i28(\rfxs[28] [31]),
    .i29(\rfxs[29] [31]),
    .i3(\rfxs[3] [31]),
    .i30(\rfxs[30] [31]),
    .i31(\rfxs[31] [31]),
    .i4(\rfxs[4] [31]),
    .i5(\rfxs[5] [31]),
    .i6(\rfxs[6] [31]),
    .i7(\rfxs[7] [31]),
    .i8(\rfxs[8] [31]),
    .i9(\rfxs[9] [31]),
    .sel(i_rs2idx),
    .o(n99[31]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b4 (
    .i0(1'b0),
    .i1(\rfxs[1] [4]),
    .i10(\rfxs[10] [4]),
    .i11(\rfxs[11] [4]),
    .i12(\rfxs[12] [4]),
    .i13(\rfxs[13] [4]),
    .i14(\rfxs[14] [4]),
    .i15(\rfxs[15] [4]),
    .i16(\rfxs[16] [4]),
    .i17(\rfxs[17] [4]),
    .i18(\rfxs[18] [4]),
    .i19(\rfxs[19] [4]),
    .i2(\rfxs[2] [4]),
    .i20(\rfxs[20] [4]),
    .i21(\rfxs[21] [4]),
    .i22(\rfxs[22] [4]),
    .i23(\rfxs[23] [4]),
    .i24(\rfxs[24] [4]),
    .i25(\rfxs[25] [4]),
    .i26(\rfxs[26] [4]),
    .i27(\rfxs[27] [4]),
    .i28(\rfxs[28] [4]),
    .i29(\rfxs[29] [4]),
    .i3(\rfxs[3] [4]),
    .i30(\rfxs[30] [4]),
    .i31(\rfxs[31] [4]),
    .i4(\rfxs[4] [4]),
    .i5(\rfxs[5] [4]),
    .i6(\rfxs[6] [4]),
    .i7(\rfxs[7] [4]),
    .i8(\rfxs[8] [4]),
    .i9(\rfxs[9] [4]),
    .sel(i_rs2idx),
    .o(n99[4]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b5 (
    .i0(1'b0),
    .i1(\rfxs[1] [5]),
    .i10(\rfxs[10] [5]),
    .i11(\rfxs[11] [5]),
    .i12(\rfxs[12] [5]),
    .i13(\rfxs[13] [5]),
    .i14(\rfxs[14] [5]),
    .i15(\rfxs[15] [5]),
    .i16(\rfxs[16] [5]),
    .i17(\rfxs[17] [5]),
    .i18(\rfxs[18] [5]),
    .i19(\rfxs[19] [5]),
    .i2(\rfxs[2] [5]),
    .i20(\rfxs[20] [5]),
    .i21(\rfxs[21] [5]),
    .i22(\rfxs[22] [5]),
    .i23(\rfxs[23] [5]),
    .i24(\rfxs[24] [5]),
    .i25(\rfxs[25] [5]),
    .i26(\rfxs[26] [5]),
    .i27(\rfxs[27] [5]),
    .i28(\rfxs[28] [5]),
    .i29(\rfxs[29] [5]),
    .i3(\rfxs[3] [5]),
    .i30(\rfxs[30] [5]),
    .i31(\rfxs[31] [5]),
    .i4(\rfxs[4] [5]),
    .i5(\rfxs[5] [5]),
    .i6(\rfxs[6] [5]),
    .i7(\rfxs[7] [5]),
    .i8(\rfxs[8] [5]),
    .i9(\rfxs[9] [5]),
    .sel(i_rs2idx),
    .o(n99[5]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b6 (
    .i0(1'b0),
    .i1(\rfxs[1] [6]),
    .i10(\rfxs[10] [6]),
    .i11(\rfxs[11] [6]),
    .i12(\rfxs[12] [6]),
    .i13(\rfxs[13] [6]),
    .i14(\rfxs[14] [6]),
    .i15(\rfxs[15] [6]),
    .i16(\rfxs[16] [6]),
    .i17(\rfxs[17] [6]),
    .i18(\rfxs[18] [6]),
    .i19(\rfxs[19] [6]),
    .i2(\rfxs[2] [6]),
    .i20(\rfxs[20] [6]),
    .i21(\rfxs[21] [6]),
    .i22(\rfxs[22] [6]),
    .i23(\rfxs[23] [6]),
    .i24(\rfxs[24] [6]),
    .i25(\rfxs[25] [6]),
    .i26(\rfxs[26] [6]),
    .i27(\rfxs[27] [6]),
    .i28(\rfxs[28] [6]),
    .i29(\rfxs[29] [6]),
    .i3(\rfxs[3] [6]),
    .i30(\rfxs[30] [6]),
    .i31(\rfxs[31] [6]),
    .i4(\rfxs[4] [6]),
    .i5(\rfxs[5] [6]),
    .i6(\rfxs[6] [6]),
    .i7(\rfxs[7] [6]),
    .i8(\rfxs[8] [6]),
    .i9(\rfxs[9] [6]),
    .sel(i_rs2idx),
    .o(n99[6]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b7 (
    .i0(1'b0),
    .i1(\rfxs[1] [7]),
    .i10(\rfxs[10] [7]),
    .i11(\rfxs[11] [7]),
    .i12(\rfxs[12] [7]),
    .i13(\rfxs[13] [7]),
    .i14(\rfxs[14] [7]),
    .i15(\rfxs[15] [7]),
    .i16(\rfxs[16] [7]),
    .i17(\rfxs[17] [7]),
    .i18(\rfxs[18] [7]),
    .i19(\rfxs[19] [7]),
    .i2(\rfxs[2] [7]),
    .i20(\rfxs[20] [7]),
    .i21(\rfxs[21] [7]),
    .i22(\rfxs[22] [7]),
    .i23(\rfxs[23] [7]),
    .i24(\rfxs[24] [7]),
    .i25(\rfxs[25] [7]),
    .i26(\rfxs[26] [7]),
    .i27(\rfxs[27] [7]),
    .i28(\rfxs[28] [7]),
    .i29(\rfxs[29] [7]),
    .i3(\rfxs[3] [7]),
    .i30(\rfxs[30] [7]),
    .i31(\rfxs[31] [7]),
    .i4(\rfxs[4] [7]),
    .i5(\rfxs[5] [7]),
    .i6(\rfxs[6] [7]),
    .i7(\rfxs[7] [7]),
    .i8(\rfxs[8] [7]),
    .i9(\rfxs[9] [7]),
    .sel(i_rs2idx),
    .o(n99[7]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b8 (
    .i0(1'b0),
    .i1(\rfxs[1] [8]),
    .i10(\rfxs[10] [8]),
    .i11(\rfxs[11] [8]),
    .i12(\rfxs[12] [8]),
    .i13(\rfxs[13] [8]),
    .i14(\rfxs[14] [8]),
    .i15(\rfxs[15] [8]),
    .i16(\rfxs[16] [8]),
    .i17(\rfxs[17] [8]),
    .i18(\rfxs[18] [8]),
    .i19(\rfxs[19] [8]),
    .i2(\rfxs[2] [8]),
    .i20(\rfxs[20] [8]),
    .i21(\rfxs[21] [8]),
    .i22(\rfxs[22] [8]),
    .i23(\rfxs[23] [8]),
    .i24(\rfxs[24] [8]),
    .i25(\rfxs[25] [8]),
    .i26(\rfxs[26] [8]),
    .i27(\rfxs[27] [8]),
    .i28(\rfxs[28] [8]),
    .i29(\rfxs[29] [8]),
    .i3(\rfxs[3] [8]),
    .i30(\rfxs[30] [8]),
    .i31(\rfxs[31] [8]),
    .i4(\rfxs[4] [8]),
    .i5(\rfxs[5] [8]),
    .i6(\rfxs[6] [8]),
    .i7(\rfxs[7] [8]),
    .i8(\rfxs[8] [8]),
    .i9(\rfxs[9] [8]),
    .sel(i_rs2idx),
    .o(n99[8]));  // ../RTL/core/regfile.v(47)
  binary_mux_s5_w1 mux34_b9 (
    .i0(1'b0),
    .i1(\rfxs[1] [9]),
    .i10(\rfxs[10] [9]),
    .i11(\rfxs[11] [9]),
    .i12(\rfxs[12] [9]),
    .i13(\rfxs[13] [9]),
    .i14(\rfxs[14] [9]),
    .i15(\rfxs[15] [9]),
    .i16(\rfxs[16] [9]),
    .i17(\rfxs[17] [9]),
    .i18(\rfxs[18] [9]),
    .i19(\rfxs[19] [9]),
    .i2(\rfxs[2] [9]),
    .i20(\rfxs[20] [9]),
    .i21(\rfxs[21] [9]),
    .i22(\rfxs[22] [9]),
    .i23(\rfxs[23] [9]),
    .i24(\rfxs[24] [9]),
    .i25(\rfxs[25] [9]),
    .i26(\rfxs[26] [9]),
    .i27(\rfxs[27] [9]),
    .i28(\rfxs[28] [9]),
    .i29(\rfxs[29] [9]),
    .i3(\rfxs[3] [9]),
    .i30(\rfxs[30] [9]),
    .i31(\rfxs[31] [9]),
    .i4(\rfxs[4] [9]),
    .i5(\rfxs[5] [9]),
    .i6(\rfxs[6] [9]),
    .i7(\rfxs[7] [9]),
    .i8(\rfxs[8] [9]),
    .i9(\rfxs[9] [9]),
    .sel(i_rs2idx),
    .o(n99[9]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b0 (
    .i0(n99[0]),
    .i1(i_rd_wdata[0]),
    .sel(n98),
    .o(n100[0]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b1 (
    .i0(n99[1]),
    .i1(i_rd_wdata[1]),
    .sel(n98),
    .o(n100[1]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b10 (
    .i0(n99[10]),
    .i1(i_rd_wdata[10]),
    .sel(n98),
    .o(n100[10]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b11 (
    .i0(n99[11]),
    .i1(i_rd_wdata[11]),
    .sel(n98),
    .o(n100[11]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b12 (
    .i0(n99[12]),
    .i1(i_rd_wdata[12]),
    .sel(n98),
    .o(n100[12]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b13 (
    .i0(n99[13]),
    .i1(i_rd_wdata[13]),
    .sel(n98),
    .o(n100[13]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b14 (
    .i0(n99[14]),
    .i1(i_rd_wdata[14]),
    .sel(n98),
    .o(n100[14]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b15 (
    .i0(n99[15]),
    .i1(i_rd_wdata[15]),
    .sel(n98),
    .o(n100[15]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b16 (
    .i0(n99[16]),
    .i1(i_rd_wdata[16]),
    .sel(n98),
    .o(n100[16]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b17 (
    .i0(n99[17]),
    .i1(i_rd_wdata[17]),
    .sel(n98),
    .o(n100[17]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b18 (
    .i0(n99[18]),
    .i1(i_rd_wdata[18]),
    .sel(n98),
    .o(n100[18]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b19 (
    .i0(n99[19]),
    .i1(i_rd_wdata[19]),
    .sel(n98),
    .o(n100[19]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b2 (
    .i0(n99[2]),
    .i1(i_rd_wdata[2]),
    .sel(n98),
    .o(n100[2]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b20 (
    .i0(n99[20]),
    .i1(i_rd_wdata[20]),
    .sel(n98),
    .o(n100[20]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b21 (
    .i0(n99[21]),
    .i1(i_rd_wdata[21]),
    .sel(n98),
    .o(n100[21]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b22 (
    .i0(n99[22]),
    .i1(i_rd_wdata[22]),
    .sel(n98),
    .o(n100[22]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b23 (
    .i0(n99[23]),
    .i1(i_rd_wdata[23]),
    .sel(n98),
    .o(n100[23]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b24 (
    .i0(n99[24]),
    .i1(i_rd_wdata[24]),
    .sel(n98),
    .o(n100[24]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b25 (
    .i0(n99[25]),
    .i1(i_rd_wdata[25]),
    .sel(n98),
    .o(n100[25]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b26 (
    .i0(n99[26]),
    .i1(i_rd_wdata[26]),
    .sel(n98),
    .o(n100[26]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b27 (
    .i0(n99[27]),
    .i1(i_rd_wdata[27]),
    .sel(n98),
    .o(n100[27]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b28 (
    .i0(n99[28]),
    .i1(i_rd_wdata[28]),
    .sel(n98),
    .o(n100[28]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b29 (
    .i0(n99[29]),
    .i1(i_rd_wdata[29]),
    .sel(n98),
    .o(n100[29]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b3 (
    .i0(n99[3]),
    .i1(i_rd_wdata[3]),
    .sel(n98),
    .o(n100[3]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b30 (
    .i0(n99[30]),
    .i1(i_rd_wdata[30]),
    .sel(n98),
    .o(n100[30]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b31 (
    .i0(n99[31]),
    .i1(i_rd_wdata[31]),
    .sel(n98),
    .o(n100[31]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b4 (
    .i0(n99[4]),
    .i1(i_rd_wdata[4]),
    .sel(n98),
    .o(n100[4]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b5 (
    .i0(n99[5]),
    .i1(i_rd_wdata[5]),
    .sel(n98),
    .o(n100[5]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b6 (
    .i0(n99[6]),
    .i1(i_rd_wdata[6]),
    .sel(n98),
    .o(n100[6]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b7 (
    .i0(n99[7]),
    .i1(i_rd_wdata[7]),
    .sel(n98),
    .o(n100[7]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b8 (
    .i0(n99[8]),
    .i1(i_rd_wdata[8]),
    .sel(n98),
    .o(n100[8]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux35_b9 (
    .i0(n99[9]),
    .i1(i_rd_wdata[9]),
    .sel(n98),
    .o(n100[9]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b0 (
    .i0(1'b0),
    .i1(n100[0]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[0]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b1 (
    .i0(1'b0),
    .i1(n100[1]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[1]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b10 (
    .i0(1'b0),
    .i1(n100[10]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[10]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b11 (
    .i0(1'b0),
    .i1(n100[11]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[11]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b12 (
    .i0(1'b0),
    .i1(n100[12]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[12]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b13 (
    .i0(1'b0),
    .i1(n100[13]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[13]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b14 (
    .i0(1'b0),
    .i1(n100[14]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[14]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b15 (
    .i0(1'b0),
    .i1(n100[15]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[15]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b16 (
    .i0(1'b0),
    .i1(n100[16]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[16]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b17 (
    .i0(1'b0),
    .i1(n100[17]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[17]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b18 (
    .i0(1'b0),
    .i1(n100[18]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[18]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b19 (
    .i0(1'b0),
    .i1(n100[19]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[19]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b2 (
    .i0(1'b0),
    .i1(n100[2]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[2]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b20 (
    .i0(1'b0),
    .i1(n100[20]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[20]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b21 (
    .i0(1'b0),
    .i1(n100[21]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[21]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b22 (
    .i0(1'b0),
    .i1(n100[22]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[22]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b23 (
    .i0(1'b0),
    .i1(n100[23]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[23]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b24 (
    .i0(1'b0),
    .i1(n100[24]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[24]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b25 (
    .i0(1'b0),
    .i1(n100[25]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[25]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b26 (
    .i0(1'b0),
    .i1(n100[26]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[26]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b27 (
    .i0(1'b0),
    .i1(n100[27]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[27]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b28 (
    .i0(1'b0),
    .i1(n100[28]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[28]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b29 (
    .i0(1'b0),
    .i1(n100[29]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[29]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b3 (
    .i0(1'b0),
    .i1(n100[3]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[3]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b30 (
    .i0(1'b0),
    .i1(n100[30]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[30]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b31 (
    .i0(1'b0),
    .i1(n100[31]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[31]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b4 (
    .i0(1'b0),
    .i1(n100[4]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[4]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b5 (
    .i0(1'b0),
    .i1(n100[5]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[5]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b6 (
    .i0(1'b0),
    .i1(n100[6]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[6]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b7 (
    .i0(1'b0),
    .i1(n100[7]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[7]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b8 (
    .i0(1'b0),
    .i1(n100[8]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[8]));  // ../RTL/core/regfile.v(47)
  binary_mux_s1_w1 mux36_b9 (
    .i0(1'b0),
    .i1(n100[9]),
    .sel(i_rs2ren),
    .o(o_rs2_rdata[9]));  // ../RTL/core/regfile.v(47)
  AL_DFF_X reg0_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg0_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[1] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg10_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n31),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[11] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg11_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n34),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[12] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg12_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n37),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[13] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg13_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n40),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[14] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg14_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n43),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[15] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg15_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n46),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[16] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg16_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n49),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[17] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg17_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n52),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[18] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg18_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n55),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[19] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg19_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n58),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[20] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg1_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n4),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[2] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg20_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n61),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[21] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg21_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n64),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[22] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg22_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n67),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[23] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg23_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n70),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[24] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg24_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n73),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[25] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg25_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n76),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[26] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg26_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n79),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[27] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg27_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n82),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[28] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg28_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n85),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[29] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg29_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n88),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[30] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg2_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n7),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[3] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg30_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n91),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[31] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg3_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n10),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[4] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg4_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n13),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[5] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg5_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n16),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[6] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg6_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n19),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[7] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg7_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n22),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[8] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg8_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n25),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[9] [9]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [0]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [1]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [10]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [11]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [12]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [13]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [14]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [15]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [16]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [17]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [18]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [19]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [2]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [20]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [21]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [22]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [23]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [24]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [25]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [26]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [27]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [28]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [29]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [3]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [30]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [31]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [4]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [5]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [6]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [7]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [8]));  // ../RTL/core/regfile.v(36)
  AL_DFF_X reg9_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .en(n28),
    .sr(1'b0),
    .ss(1'b0),
    .q(\rfxs[10] [9]));  // ../RTL/core/regfile.v(36)
  and u133 (n7, i_rdwen, n6);  // ../RTL/core/regfile.v(37)
  and u197 (n10, i_rdwen, n9);  // ../RTL/core/regfile.v(37)
  and u261 (n13, i_rdwen, n12);  // ../RTL/core/regfile.v(37)
  and u325 (n16, i_rdwen, n15);  // ../RTL/core/regfile.v(37)
  and u389 (n19, i_rdwen, n18);  // ../RTL/core/regfile.v(37)
  and u453 (n22, i_rdwen, n21);  // ../RTL/core/regfile.v(37)
  and u5 (n1, i_rdwen, n0);  // ../RTL/core/regfile.v(37)
  and u517 (n25, i_rdwen, n24);  // ../RTL/core/regfile.v(37)
  and u581 (n28, i_rdwen, n27);  // ../RTL/core/regfile.v(37)
  and u645 (n31, i_rdwen, n30);  // ../RTL/core/regfile.v(37)
  and u69 (n4, i_rdwen, n3);  // ../RTL/core/regfile.v(37)
  and u709 (n34, i_rdwen, n33);  // ../RTL/core/regfile.v(37)
  and u773 (n37, i_rdwen, n36);  // ../RTL/core/regfile.v(37)
  and u837 (n40, i_rdwen, n39);  // ../RTL/core/regfile.v(37)
  and u901 (n43, i_rdwen, n42);  // ../RTL/core/regfile.v(37)
  and u963 (n46, i_rdwen, n45);  // ../RTL/core/regfile.v(37)
  and u965 (n49, i_rdwen, n48);  // ../RTL/core/regfile.v(37)
  and u967 (n52, i_rdwen, n51);  // ../RTL/core/regfile.v(37)
  and u969 (n55, i_rdwen, n54);  // ../RTL/core/regfile.v(37)
  and u971 (n58, i_rdwen, n57);  // ../RTL/core/regfile.v(37)
  and u973 (n61, i_rdwen, n60);  // ../RTL/core/regfile.v(37)
  and u975 (n64, i_rdwen, n63);  // ../RTL/core/regfile.v(37)
  and u977 (n67, i_rdwen, n66);  // ../RTL/core/regfile.v(37)
  and u979 (n70, i_rdwen, n69);  // ../RTL/core/regfile.v(37)
  and u981 (n73, i_rdwen, n72);  // ../RTL/core/regfile.v(37)
  and u983 (n76, i_rdwen, n75);  // ../RTL/core/regfile.v(37)
  and u985 (n79, i_rdwen, n78);  // ../RTL/core/regfile.v(37)
  and u987 (n82, i_rdwen, n81);  // ../RTL/core/regfile.v(37)
  and u989 (n85, i_rdwen, n84);  // ../RTL/core/regfile.v(37)
  and u991 (n88, i_rdwen, n87);  // ../RTL/core/regfile.v(37)
  and u993 (n91, i_rdwen, n90);  // ../RTL/core/regfile.v(37)
  and u994 (n94, n93, i_rdwen);  // ../RTL/core/regfile.v(46)
  and u995 (n98, n97, i_rdwen);  // ../RTL/core/regfile.v(47)

endmodule 

module FPU32  // ../RTL/core/fpu.v(7)
  (
  i_clk,
  i_op1,
  i_op2,
  i_rsn,
  o_addres,
  o_divres,
  o_mulres,
  o_subres
  );

  input i_clk;  // ../RTL/core/fpu.v(8)
  input [31:0] i_op1;  // ../RTL/core/fpu.v(11)
  input [31:0] i_op2;  // ../RTL/core/fpu.v(12)
  input i_rsn;  // ../RTL/core/fpu.v(9)
  output [31:0] o_addres;  // ../RTL/core/fpu.v(15)
  output [31:0] o_divres;  // ../RTL/core/fpu.v(18)
  output [31:0] o_mulres;  // ../RTL/core/fpu.v(17)
  output [31:0] o_subres;  // ../RTL/core/fpu.v(16)

  wire [47:0] \u_mul/M_mul_result ;  // ../RTL/core/fpu.v(253)
  wire [23:0] \u_mul/normalized_M_mul_result ;  // ../RTL/core/fpu.v(254)
  wire [8:0] \u_mul/sum_E ;  // ../RTL/core/fpu.v(252)
  wire \u_mul/ADD01/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD01/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD01/n1 ;
  wire \u_mul/ADD01/ADD01/n12 ;
  wire \u_mul/ADD01/ADD01/n13 ;
  wire \u_mul/ADD01/ADD01/n14 ;
  wire \u_mul/ADD01/ADD01/n15 ;
  wire \u_mul/ADD01/ADD01/n16 ;
  wire \u_mul/ADD01/ADD01/n17 ;
  wire \u_mul/ADD01/ADD01/n18 ;
  wire \u_mul/ADD01/ADD01/n19 ;
  wire \u_mul/ADD01/ADD01/n2 ;
  wire \u_mul/ADD01/ADD01/n5 ;
  wire \u_mul/ADD01/ADD01/n6 ;
  wire \u_mul/ADD01/ADD01/n7 ;
  wire \u_mul/ADD01/ADD01/n8 ;
  wire \u_mul/ADD01/ADD01/n9 ;
  wire \u_mul/ADD01/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD01/p0_neg ;
  wire \u_mul/ADD01/ADD01/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD01/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD01/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD02/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD02/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD02/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD02/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD02/n0 ;
  wire \u_mul/ADD01/ADD02/n1 ;
  wire \u_mul/ADD01/ADD02/n10 ;
  wire \u_mul/ADD01/ADD02/n11 ;
  wire \u_mul/ADD01/ADD02/n2 ;
  wire \u_mul/ADD01/ADD02/n3 ;
  wire \u_mul/ADD01/ADD02/n4 ;
  wire \u_mul/ADD01/ADD02/n5 ;
  wire \u_mul/ADD01/ADD02/n6 ;
  wire \u_mul/ADD01/ADD02/n7 ;
  wire \u_mul/ADD01/ADD02/n8 ;
  wire \u_mul/ADD01/ADD02/n9 ;
  wire \u_mul/ADD01/ADD02/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD02/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD02/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD01/ADD02/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD02/ADD01/ADD01/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD02/ADD01/ADD01/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD02/ADD01/ADD01/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD02/ADD01/ADD01/n0 ;
  wire \u_mul/ADD02/ADD01/ADD01/n1 ;
  wire \u_mul/ADD02/ADD01/ADD01/n10 ;
  wire \u_mul/ADD02/ADD01/ADD01/n11 ;
  wire \u_mul/ADD02/ADD01/ADD01/n14 ;
  wire \u_mul/ADD02/ADD01/ADD01/n17 ;
  wire \u_mul/ADD02/ADD01/ADD01/n18 ;
  wire \u_mul/ADD02/ADD01/ADD01/n20 ;
  wire \u_mul/ADD02/ADD01/ADD01/n21 ;
  wire \u_mul/ADD02/ADD01/ADD01/n3 ;
  wire \u_mul/ADD02/ADD01/ADD01/n4 ;
  wire \u_mul/ADD02/ADD01/ADD01/n7 ;
  wire \u_mul/ADD02/ADD01/ADD01/n8 ;
  wire \u_mul/ADD02/ADD01/ADD02/n0 ;
  wire \u_mul/ADD02/ADD01/ADD02/n10 ;
  wire \u_mul/ADD02/ADD01/ADD02/n11 ;
  wire \u_mul/ADD02/ADD01/ADD02/n3 ;
  wire \u_mul/ADD02/ADD01/ADD02/n4 ;
  wire \u_mul/ADD02/ADD01/ADD02/n7 ;
  wire \u_mul/ADD02/ADD01/ctemp ;  // ../RTL/core/fpu_utils.v(76)
  wire \u_mul/ADD23/ADD01/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD23/ADD01/ADD01/n1 ;
  wire \u_mul/ADD23/ADD01/ADD01/n14 ;
  wire \u_mul/ADD23/ADD01/ADD01/n17 ;
  wire \u_mul/ADD23/ADD01/ADD01/n18 ;
  wire \u_mul/ADD23/ADD01/ADD01/n7 ;
  wire \u_mul/ADD23/ADD01/ADD01/n8 ;
  wire \u_mul/ADD23/ADD01/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD23/ADD01/ADD02/n0 ;
  wire \u_mul/ADD23/ADD01/ADD02/n10 ;
  wire \u_mul/ADD23/ADD01/ADD02/n11 ;
  wire \u_mul/ADD23/ADD01/ADD02/n14 ;
  wire \u_mul/ADD23/ADD01/ADD02/n17 ;
  wire \u_mul/ADD23/ADD01/ADD02/n20 ;
  wire \u_mul/ADD23/ADD01/ADD02/n21 ;
  wire \u_mul/ADD23/ADD01/ADD02/n3 ;
  wire \u_mul/ADD23/ADD01/ADD02/n4 ;
  wire \u_mul/ADD23/ADD01/ADD02/n7 ;
  wire \u_mul/ADD23/ADD02/ADD01/n0 ;
  wire \u_mul/ADD23/ADD02/ADD01/n10 ;
  wire \u_mul/ADD23/ADD02/ADD01/n11 ;
  wire \u_mul/ADD23/ADD02/ADD01/n14 ;
  wire \u_mul/ADD23/ADD02/ADD01/n17 ;
  wire \u_mul/ADD23/ADD02/ADD01/n20 ;
  wire \u_mul/ADD23/ADD02/ADD01/n21 ;
  wire \u_mul/ADD23/ADD02/ADD01/n3 ;
  wire \u_mul/ADD23/ADD02/ADD01/n4 ;
  wire \u_mul/ADD23/ADD02/ADD01/n7 ;
  wire \u_mul/ADD23/ADD02/ADD02/n0 ;
  wire \u_mul/ADD23/ADD02/ADD02/n10 ;
  wire \u_mul/ADD23/ADD02/ADD02/n11 ;
  wire \u_mul/ADD23/ADD02/ADD02/n14 ;
  wire \u_mul/ADD23/ADD02/ADD02/n17 ;
  wire \u_mul/ADD23/ADD02/ADD02/n20 ;
  wire \u_mul/ADD23/ADD02/ADD02/n21 ;
  wire \u_mul/ADD23/ADD02/ADD02/n3 ;
  wire \u_mul/ADD23/ADD02/ADD02/n4 ;
  wire \u_mul/ADD23/ADD02/ADD02/n7 ;
  wire \u_mul/ADD23/ADD03/ADD01/n0 ;
  wire \u_mul/ADD23/ADD03/ADD01/n10 ;
  wire \u_mul/ADD23/ADD03/ADD01/n11 ;
  wire \u_mul/ADD23/ADD03/ADD01/n14 ;
  wire \u_mul/ADD23/ADD03/ADD01/n17 ;
  wire \u_mul/ADD23/ADD03/ADD01/n20 ;
  wire \u_mul/ADD23/ADD03/ADD01/n21 ;
  wire \u_mul/ADD23/ADD03/ADD01/n3 ;
  wire \u_mul/ADD23/ADD03/ADD01/n4 ;
  wire \u_mul/ADD23/ADD03/ADD01/n7 ;
  wire \u_mul/ADD23/ADD03/ADD02/n0 ;
  wire \u_mul/ADD23/ADD03/ADD02/n3 ;
  wire \u_mul/ADD23/ADD03/ADD02/n4 ;
  wire \u_mul/RO01/w1 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO01/w2 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO01/w3 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO01/w4 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO01/w5 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO01/w6 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO01/w1 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO01/w2 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO01/w3 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO01/w4 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO01/w5 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO01/w6 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO02/w1 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO02/w2 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO02/w3 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO02/w4 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO02/w5 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO02/w6 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO03/w1 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO03/w2 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO03/w3 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO03/w4 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO03/w5 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/RO03/w6 ;  // ../RTL/core/fpu_utils.v(13)
  wire \u_mul/RO03/n0 ;
  wire \u_mul/RO03/o1 ;  // ../RTL/core/fpu_utils.v(24)
  wire \u_mul/RO03/o2 ;  // ../RTL/core/fpu_utils.v(25)
  wire \u_mul/RO04/o3 ;  // ../RTL/core/fpu_utils.v(26)
  wire \u_mul/final_product_round ;  // ../RTL/core/fpu.v(280)
  wire \u_mul/mul_round1 ;  // ../RTL/core/fpu.v(278)
  wire \u_mul/mul_round2 ;  // ../RTL/core/fpu.v(279)
  wire \u_mul/reduced_or_E1 ;  // ../RTL/core/fpu.v(256)
  wire \u_mul/sum_E[7]_neg ;

  assign o_mulres[0] = \u_mul/ADD23/ADD01/ADD01/p0 ;
  add_sub_1 u_add (
    .n1(i_op1),
    .n2(i_op2),
    .sub(1'b0),
    .result(o_addres));  // ../RTL/core/fpu.v(23)
  not \u_mul/ADD01/ADD01/p0_inv  (\u_mul/ADD01/ADD01/p0_neg , \u_mul/ADD01/ADD01/p0 );
  and \u_mul/ADD01/ADD01/u0  (\u_mul/ADD01/ADD01/g0 , i_op1[23], i_op2[23]);  // ../RTL/core/fpu_utils.v(55)
  and \u_mul/ADD01/ADD01/u1  (\u_mul/ADD01/ADD01/g1 , i_op1[24], i_op2[24]);  // ../RTL/core/fpu_utils.v(56)
  and \u_mul/ADD01/ADD01/u10  (\u_mul/ADD01/ADD01/n1 , \u_mul/ADD01/ADD01/p1 , \u_mul/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \u_mul/ADD01/ADD01/u11  (\u_mul/ADD01/ADD01/n2 , \u_mul/ADD01/ADD01/g1 , \u_mul/ADD01/ADD01/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD01/ADD01/u15  (\u_mul/ADD01/ADD01/n5 , \u_mul/ADD01/ADD01/p2 , \u_mul/ADD01/ADD01/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \u_mul/ADD01/ADD01/u16  (\u_mul/ADD01/ADD01/n6 , \u_mul/ADD01/ADD01/g2 , \u_mul/ADD01/ADD01/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD01/ADD01/u17  (\u_mul/ADD01/ADD01/n7 , \u_mul/ADD01/ADD01/p2 , \u_mul/ADD01/ADD01/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD01/ADD01/u18  (\u_mul/ADD01/ADD01/n8 , \u_mul/ADD01/ADD01/n7 , \u_mul/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \u_mul/ADD01/ADD01/u19  (\u_mul/ADD01/ADD01/n9 , \u_mul/ADD01/ADD01/n6 , \u_mul/ADD01/ADD01/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD01/ADD01/u2  (\u_mul/ADD01/ADD01/g2 , i_op1[25], i_op2[25]);  // ../RTL/core/fpu_utils.v(57)
  xor \u_mul/ADD01/ADD01/u20  (\u_mul/sum_E [3], \u_mul/ADD01/ADD01/p3 , \u_mul/ADD01/ADD01/n9 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD01/ADD01/u24  (\u_mul/ADD01/ADD01/n12 , \u_mul/ADD01/ADD01/p3 , \u_mul/ADD01/ADD01/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \u_mul/ADD01/ADD01/u25  (\u_mul/ADD01/ADD01/n13 , \u_mul/ADD01/ADD01/g3 , \u_mul/ADD01/ADD01/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD01/ADD01/u26  (\u_mul/ADD01/ADD01/n14 , \u_mul/ADD01/ADD01/p3 , \u_mul/ADD01/ADD01/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD01/ADD01/u27  (\u_mul/ADD01/ADD01/n15 , \u_mul/ADD01/ADD01/n14 , \u_mul/ADD01/ADD01/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \u_mul/ADD01/ADD01/u28  (\u_mul/ADD01/ADD01/n16 , \u_mul/ADD01/ADD01/n13 , \u_mul/ADD01/ADD01/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD01/ADD01/u29  (\u_mul/sum_E [2], \u_mul/ADD01/ADD01/p2 , \u_mul/ADD01/ADD01/n2 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD01/ADD01/u3  (\u_mul/ADD01/ADD01/g3 , i_op1[26], i_op2[26]);  // ../RTL/core/fpu_utils.v(58)
  and \u_mul/ADD01/ADD01/u30  (\u_mul/ADD01/ADD01/n17 , \u_mul/ADD01/ADD01/n14 , \u_mul/ADD01/ADD01/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD01/ADD01/u31  (\u_mul/ADD01/ADD01/n18 , \u_mul/ADD01/ADD01/n17 , \u_mul/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \u_mul/ADD01/ADD01/u32  (\u_mul/ADD01/ADD01/n19 , \u_mul/ADD01/ADD01/n16 , \u_mul/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD01/ADD01/u33  (\u_mul/sum_E [1], \u_mul/ADD01/ADD01/p1 , \u_mul/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD01/ADD01/u4  (\u_mul/ADD01/ADD01/p0 , i_op1[23], i_op2[23]);  // ../RTL/core/fpu_utils.v(59)
  xor \u_mul/ADD01/ADD01/u5  (\u_mul/ADD01/ADD01/p1 , i_op1[24], i_op2[24]);  // ../RTL/core/fpu_utils.v(60)
  xor \u_mul/ADD01/ADD01/u6  (\u_mul/ADD01/ADD01/p2 , i_op1[25], i_op2[25]);  // ../RTL/core/fpu_utils.v(61)
  xor \u_mul/ADD01/ADD01/u7  (\u_mul/ADD01/ADD01/p3 , i_op1[26], i_op2[26]);  // ../RTL/core/fpu_utils.v(62)
  and \u_mul/ADD01/ADD02/u0  (\u_mul/ADD01/ADD02/g0 , i_op1[27], i_op2[27]);  // ../RTL/core/fpu_utils.v(55)
  and \u_mul/ADD01/ADD02/u1  (\u_mul/ADD01/ADD02/g1 , i_op1[28], i_op2[28]);  // ../RTL/core/fpu_utils.v(56)
  and \u_mul/ADD01/ADD02/u10  (\u_mul/ADD01/ADD02/n1 , \u_mul/ADD01/ADD02/p1 , \u_mul/ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \u_mul/ADD01/ADD02/u11  (\u_mul/ADD01/ADD02/n2 , \u_mul/ADD01/ADD02/g1 , \u_mul/ADD01/ADD02/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD01/ADD02/u12  (\u_mul/ADD01/ADD02/n3 , \u_mul/ADD01/ADD02/p1 , \u_mul/ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD01/ADD02/u13  (\u_mul/ADD01/ADD02/n4 , \u_mul/ADD01/ADD02/n3 , \u_mul/ADD01/ADD01/n19 );  // ../RTL/core/fpu_utils.v(64)
  or \u_mul/ADD01/ADD02/u14  (\u_mul/ADD01/ADD02/c1 , \u_mul/ADD01/ADD02/n2 , \u_mul/ADD01/ADD02/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD01/ADD02/u15  (\u_mul/ADD01/ADD02/n5 , \u_mul/ADD01/ADD02/p2 , \u_mul/ADD01/ADD02/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \u_mul/ADD01/ADD02/u16  (\u_mul/ADD01/ADD02/n6 , \u_mul/ADD01/ADD02/g2 , \u_mul/ADD01/ADD02/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD01/ADD02/u17  (\u_mul/ADD01/ADD02/n7 , \u_mul/ADD01/ADD02/p2 , \u_mul/ADD01/ADD02/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD01/ADD02/u18  (\u_mul/ADD01/ADD02/n8 , \u_mul/ADD01/ADD02/n7 , \u_mul/ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \u_mul/ADD01/ADD02/u19  (\u_mul/ADD01/ADD02/n9 , \u_mul/ADD01/ADD02/n6 , \u_mul/ADD01/ADD02/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD01/ADD02/u2  (\u_mul/ADD01/ADD02/g2 , i_op1[29], i_op2[29]);  // ../RTL/core/fpu_utils.v(57)
  xor \u_mul/ADD01/ADD02/u20  (\u_mul/sum_E [7], \u_mul/ADD01/ADD02/p3 , \u_mul/ADD01/ADD02/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD01/ADD02/u21  (\u_mul/ADD01/ADD02/n10 , \u_mul/ADD01/ADD02/n7 , \u_mul/ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD01/ADD02/u22  (\u_mul/ADD01/ADD02/n11 , \u_mul/ADD01/ADD02/n10 , \u_mul/ADD01/ADD01/n19 );  // ../RTL/core/fpu_utils.v(65)
  or \u_mul/ADD01/ADD02/u23  (\u_mul/ADD01/ADD02/c2 , \u_mul/ADD01/ADD02/n9 , \u_mul/ADD01/ADD02/n11 );  // ../RTL/core/fpu_utils.v(65)
  xor \u_mul/ADD01/ADD02/u29  (\u_mul/sum_E [6], \u_mul/ADD01/ADD02/p2 , \u_mul/ADD01/ADD02/c1 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD01/ADD02/u33  (\u_mul/sum_E [5], \u_mul/ADD01/ADD02/p1 , \u_mul/ADD01/ADD02/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD01/ADD02/u34  (\u_mul/sum_E [4], \u_mul/ADD01/ADD02/p0 , \u_mul/ADD01/ADD01/n19 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD01/ADD02/u4  (\u_mul/ADD01/ADD02/p0 , i_op1[27], i_op2[27]);  // ../RTL/core/fpu_utils.v(59)
  xor \u_mul/ADD01/ADD02/u5  (\u_mul/ADD01/ADD02/p1 , i_op1[28], i_op2[28]);  // ../RTL/core/fpu_utils.v(60)
  xor \u_mul/ADD01/ADD02/u6  (\u_mul/ADD01/ADD02/p2 , i_op1[29], i_op2[29]);  // ../RTL/core/fpu_utils.v(61)
  xor \u_mul/ADD01/ADD02/u7  (\u_mul/ADD01/ADD02/p3 , i_op1[30], i_op2[30]);  // ../RTL/core/fpu_utils.v(62)
  and \u_mul/ADD01/ADD02/u8  (\u_mul/ADD01/ADD02/n0 , \u_mul/ADD01/ADD02/p0 , \u_mul/ADD01/ADD01/n19 );  // ../RTL/core/fpu_utils.v(63)
  or \u_mul/ADD01/ADD02/u9  (\u_mul/ADD01/ADD02/c0 , \u_mul/ADD01/ADD02/g0 , \u_mul/ADD01/ADD02/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \u_mul/ADD02/ADD01/ADD01/u10  (\u_mul/ADD02/ADD01/ADD01/n1 , \u_mul/sum_E [1], \u_mul/ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD02/ADD01/ADD01/u12  (\u_mul/ADD02/ADD01/ADD01/n3 , \u_mul/sum_E [1], \u_mul/ADD01/ADD01/p0_neg );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD02/ADD01/ADD01/u13  (\u_mul/ADD02/ADD01/ADD01/n4 , \u_mul/ADD02/ADD01/ADD01/n3 , \u_mul/M_mul_result [47]);  // ../RTL/core/fpu_utils.v(64)
  or \u_mul/ADD02/ADD01/ADD01/u14  (\u_mul/ADD02/ADD01/ADD01/c1 , \u_mul/ADD02/ADD01/ADD01/n1 , \u_mul/ADD02/ADD01/ADD01/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD02/ADD01/ADD01/u17  (\u_mul/ADD02/ADD01/ADD01/n7 , \u_mul/sum_E [2], \u_mul/sum_E [1]);  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD02/ADD01/ADD01/u18  (\u_mul/ADD02/ADD01/ADD01/n8 , \u_mul/ADD02/ADD01/ADD01/n7 , \u_mul/ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  xor \u_mul/ADD02/ADD01/ADD01/u20  (o_mulres[26], \u_mul/sum_E [3], \u_mul/ADD02/ADD01/ADD01/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD02/ADD01/ADD01/u21  (\u_mul/ADD02/ADD01/ADD01/n10 , \u_mul/ADD02/ADD01/ADD01/n7 , \u_mul/ADD01/ADD01/p0_neg );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD02/ADD01/ADD01/u22  (\u_mul/ADD02/ADD01/ADD01/n11 , \u_mul/ADD02/ADD01/ADD01/n10 , \u_mul/M_mul_result [47]);  // ../RTL/core/fpu_utils.v(65)
  or \u_mul/ADD02/ADD01/ADD01/u23  (\u_mul/ADD02/ADD01/ADD01/c2 , \u_mul/ADD02/ADD01/ADD01/n8 , \u_mul/ADD02/ADD01/ADD01/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD02/ADD01/ADD01/u26  (\u_mul/ADD02/ADD01/ADD01/n14 , \u_mul/sum_E [3], \u_mul/sum_E [2]);  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD02/ADD01/ADD01/u29  (o_mulres[25], \u_mul/sum_E [2], \u_mul/ADD02/ADD01/ADD01/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD02/ADD01/ADD01/u30  (\u_mul/ADD02/ADD01/ADD01/n17 , \u_mul/ADD02/ADD01/ADD01/n14 , \u_mul/sum_E [1]);  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD02/ADD01/ADD01/u31  (\u_mul/ADD02/ADD01/ADD01/n18 , \u_mul/ADD02/ADD01/ADD01/n17 , \u_mul/ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD02/ADD01/ADD01/u33  (o_mulres[24], \u_mul/sum_E [1], \u_mul/ADD02/ADD01/ADD01/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD02/ADD01/ADD01/u34  (o_mulres[23], \u_mul/ADD01/ADD01/p0_neg , \u_mul/M_mul_result [47]);  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD02/ADD01/ADD01/u35  (\u_mul/ADD02/ADD01/ADD01/n20 , \u_mul/ADD02/ADD01/ADD01/n17 , \u_mul/ADD01/ADD01/p0_neg );  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD02/ADD01/ADD01/u36  (\u_mul/ADD02/ADD01/ADD01/n21 , \u_mul/ADD02/ADD01/ADD01/n20 , \u_mul/M_mul_result [47]);  // ../RTL/core/fpu_utils.v(66)
  or \u_mul/ADD02/ADD01/ADD01/u37  (\u_mul/ADD02/ADD01/ctemp , \u_mul/ADD02/ADD01/ADD01/n18 , \u_mul/ADD02/ADD01/ADD01/n21 );  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD02/ADD01/ADD01/u8  (\u_mul/ADD02/ADD01/ADD01/n0 , \u_mul/ADD01/ADD01/p0_neg , \u_mul/M_mul_result [47]);  // ../RTL/core/fpu_utils.v(63)
  or \u_mul/ADD02/ADD01/ADD01/u9  (\u_mul/ADD02/ADD01/ADD01/c0 , \u_mul/ADD01/ADD01/p0 , \u_mul/ADD02/ADD01/ADD01/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \u_mul/ADD02/ADD01/ADD02/u12  (\u_mul/ADD02/ADD01/ADD02/n3 , \u_mul/sum_E [5], \u_mul/sum_E [4]);  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD02/ADD01/ADD02/u13  (\u_mul/ADD02/ADD01/ADD02/n4 , \u_mul/ADD02/ADD01/ADD02/n3 , \u_mul/ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD02/ADD01/ADD02/u17  (\u_mul/ADD02/ADD01/ADD02/n7 , \u_mul/sum_E [6], \u_mul/sum_E [5]);  // ../RTL/core/fpu_utils.v(65)
  xor \u_mul/ADD02/ADD01/ADD02/u20  (o_mulres[30], \u_mul/sum_E[7]_neg , \u_mul/ADD02/ADD01/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD02/ADD01/ADD02/u21  (\u_mul/ADD02/ADD01/ADD02/n10 , \u_mul/ADD02/ADD01/ADD02/n7 , \u_mul/sum_E [4]);  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD02/ADD01/ADD02/u22  (\u_mul/ADD02/ADD01/ADD02/n11 , \u_mul/ADD02/ADD01/ADD02/n10 , \u_mul/ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(65)
  xor \u_mul/ADD02/ADD01/ADD02/u29  (o_mulres[29], \u_mul/sum_E [6], \u_mul/ADD02/ADD01/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD02/ADD01/ADD02/u33  (o_mulres[28], \u_mul/sum_E [5], \u_mul/ADD02/ADD01/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD02/ADD01/ADD02/u34  (o_mulres[27], \u_mul/sum_E [4], \u_mul/ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD02/ADD01/ADD02/u8  (\u_mul/ADD02/ADD01/ADD02/n0 , \u_mul/sum_E [4], \u_mul/ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(63)
  and \u_mul/ADD23/ADD01/ADD01/u0  (\u_mul/ADD23/ADD01/ADD01/g0 , \u_mul/normalized_M_mul_result [0], \u_mul/final_product_round );  // ../RTL/core/fpu_utils.v(55)
  and \u_mul/ADD23/ADD01/ADD01/u10  (\u_mul/ADD23/ADD01/ADD01/n1 , \u_mul/normalized_M_mul_result [1], \u_mul/ADD23/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD23/ADD01/ADD01/u17  (\u_mul/ADD23/ADD01/ADD01/n7 , \u_mul/normalized_M_mul_result [2], \u_mul/normalized_M_mul_result [1]);  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD23/ADD01/ADD01/u18  (\u_mul/ADD23/ADD01/ADD01/n8 , \u_mul/ADD23/ADD01/ADD01/n7 , \u_mul/ADD23/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(65)
  xor \u_mul/ADD23/ADD01/ADD01/u20  (o_mulres[3], \u_mul/normalized_M_mul_result [3], \u_mul/ADD23/ADD01/ADD01/n8 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD01/ADD01/u26  (\u_mul/ADD23/ADD01/ADD01/n14 , \u_mul/normalized_M_mul_result [3], \u_mul/normalized_M_mul_result [2]);  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD23/ADD01/ADD01/u29  (o_mulres[2], \u_mul/normalized_M_mul_result [2], \u_mul/ADD23/ADD01/ADD01/n1 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD01/ADD01/u30  (\u_mul/ADD23/ADD01/ADD01/n17 , \u_mul/ADD23/ADD01/ADD01/n14 , \u_mul/normalized_M_mul_result [1]);  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD23/ADD01/ADD01/u31  (\u_mul/ADD23/ADD01/ADD01/n18 , \u_mul/ADD23/ADD01/ADD01/n17 , \u_mul/ADD23/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD23/ADD01/ADD01/u33  (o_mulres[1], \u_mul/normalized_M_mul_result [1], \u_mul/ADD23/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD23/ADD01/ADD01/u4  (\u_mul/ADD23/ADD01/ADD01/p0 , \u_mul/normalized_M_mul_result [0], \u_mul/final_product_round );  // ../RTL/core/fpu_utils.v(59)
  and \u_mul/ADD23/ADD01/ADD02/u12  (\u_mul/ADD23/ADD01/ADD02/n3 , \u_mul/normalized_M_mul_result [5], \u_mul/normalized_M_mul_result [4]);  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD23/ADD01/ADD02/u13  (\u_mul/ADD23/ADD01/ADD02/n4 , \u_mul/ADD23/ADD01/ADD02/n3 , \u_mul/ADD23/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD23/ADD01/ADD02/u17  (\u_mul/ADD23/ADD01/ADD02/n7 , \u_mul/normalized_M_mul_result [6], \u_mul/normalized_M_mul_result [5]);  // ../RTL/core/fpu_utils.v(65)
  xor \u_mul/ADD23/ADD01/ADD02/u20  (o_mulres[7], \u_mul/normalized_M_mul_result [7], \u_mul/ADD23/ADD01/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD01/ADD02/u21  (\u_mul/ADD23/ADD01/ADD02/n10 , \u_mul/ADD23/ADD01/ADD02/n7 , \u_mul/normalized_M_mul_result [4]);  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD23/ADD01/ADD02/u22  (\u_mul/ADD23/ADD01/ADD02/n11 , \u_mul/ADD23/ADD01/ADD02/n10 , \u_mul/ADD23/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD23/ADD01/ADD02/u26  (\u_mul/ADD23/ADD01/ADD02/n14 , \u_mul/normalized_M_mul_result [7], \u_mul/normalized_M_mul_result [6]);  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD23/ADD01/ADD02/u29  (o_mulres[6], \u_mul/normalized_M_mul_result [6], \u_mul/ADD23/ADD01/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD01/ADD02/u30  (\u_mul/ADD23/ADD01/ADD02/n17 , \u_mul/ADD23/ADD01/ADD02/n14 , \u_mul/normalized_M_mul_result [5]);  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD23/ADD01/ADD02/u33  (o_mulres[5], \u_mul/normalized_M_mul_result [5], \u_mul/ADD23/ADD01/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD23/ADD01/ADD02/u34  (o_mulres[4], \u_mul/normalized_M_mul_result [4], \u_mul/ADD23/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD01/ADD02/u35  (\u_mul/ADD23/ADD01/ADD02/n20 , \u_mul/ADD23/ADD01/ADD02/n17 , \u_mul/normalized_M_mul_result [4]);  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD23/ADD01/ADD02/u36  (\u_mul/ADD23/ADD01/ADD02/n21 , \u_mul/ADD23/ADD01/ADD02/n20 , \u_mul/ADD23/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD23/ADD01/ADD02/u8  (\u_mul/ADD23/ADD01/ADD02/n0 , \u_mul/normalized_M_mul_result [4], \u_mul/ADD23/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(63)
  and \u_mul/ADD23/ADD02/ADD01/u12  (\u_mul/ADD23/ADD02/ADD01/n3 , \u_mul/normalized_M_mul_result [9], \u_mul/normalized_M_mul_result [8]);  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD23/ADD02/ADD01/u13  (\u_mul/ADD23/ADD02/ADD01/n4 , \u_mul/ADD23/ADD02/ADD01/n3 , \u_mul/ADD23/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD23/ADD02/ADD01/u17  (\u_mul/ADD23/ADD02/ADD01/n7 , \u_mul/normalized_M_mul_result [10], \u_mul/normalized_M_mul_result [9]);  // ../RTL/core/fpu_utils.v(65)
  xor \u_mul/ADD23/ADD02/ADD01/u20  (o_mulres[11], \u_mul/normalized_M_mul_result [11], \u_mul/ADD23/ADD02/ADD01/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD02/ADD01/u21  (\u_mul/ADD23/ADD02/ADD01/n10 , \u_mul/ADD23/ADD02/ADD01/n7 , \u_mul/normalized_M_mul_result [8]);  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD23/ADD02/ADD01/u22  (\u_mul/ADD23/ADD02/ADD01/n11 , \u_mul/ADD23/ADD02/ADD01/n10 , \u_mul/ADD23/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD23/ADD02/ADD01/u26  (\u_mul/ADD23/ADD02/ADD01/n14 , \u_mul/normalized_M_mul_result [11], \u_mul/normalized_M_mul_result [10]);  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD23/ADD02/ADD01/u29  (o_mulres[10], \u_mul/normalized_M_mul_result [10], \u_mul/ADD23/ADD02/ADD01/n4 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD02/ADD01/u30  (\u_mul/ADD23/ADD02/ADD01/n17 , \u_mul/ADD23/ADD02/ADD01/n14 , \u_mul/normalized_M_mul_result [9]);  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD23/ADD02/ADD01/u33  (o_mulres[9], \u_mul/normalized_M_mul_result [9], \u_mul/ADD23/ADD02/ADD01/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD23/ADD02/ADD01/u34  (o_mulres[8], \u_mul/normalized_M_mul_result [8], \u_mul/ADD23/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD02/ADD01/u35  (\u_mul/ADD23/ADD02/ADD01/n20 , \u_mul/ADD23/ADD02/ADD01/n17 , \u_mul/normalized_M_mul_result [8]);  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD23/ADD02/ADD01/u36  (\u_mul/ADD23/ADD02/ADD01/n21 , \u_mul/ADD23/ADD02/ADD01/n20 , \u_mul/ADD23/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD23/ADD02/ADD01/u8  (\u_mul/ADD23/ADD02/ADD01/n0 , \u_mul/normalized_M_mul_result [8], \u_mul/ADD23/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(63)
  and \u_mul/ADD23/ADD02/ADD02/u12  (\u_mul/ADD23/ADD02/ADD02/n3 , \u_mul/normalized_M_mul_result [13], \u_mul/normalized_M_mul_result [12]);  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD23/ADD02/ADD02/u13  (\u_mul/ADD23/ADD02/ADD02/n4 , \u_mul/ADD23/ADD02/ADD02/n3 , \u_mul/ADD23/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD23/ADD02/ADD02/u17  (\u_mul/ADD23/ADD02/ADD02/n7 , \u_mul/normalized_M_mul_result [14], \u_mul/normalized_M_mul_result [13]);  // ../RTL/core/fpu_utils.v(65)
  xor \u_mul/ADD23/ADD02/ADD02/u20  (o_mulres[15], \u_mul/normalized_M_mul_result [15], \u_mul/ADD23/ADD02/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD02/ADD02/u21  (\u_mul/ADD23/ADD02/ADD02/n10 , \u_mul/ADD23/ADD02/ADD02/n7 , \u_mul/normalized_M_mul_result [12]);  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD23/ADD02/ADD02/u22  (\u_mul/ADD23/ADD02/ADD02/n11 , \u_mul/ADD23/ADD02/ADD02/n10 , \u_mul/ADD23/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD23/ADD02/ADD02/u26  (\u_mul/ADD23/ADD02/ADD02/n14 , \u_mul/normalized_M_mul_result [15], \u_mul/normalized_M_mul_result [14]);  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD23/ADD02/ADD02/u29  (o_mulres[14], \u_mul/normalized_M_mul_result [14], \u_mul/ADD23/ADD02/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD02/ADD02/u30  (\u_mul/ADD23/ADD02/ADD02/n17 , \u_mul/ADD23/ADD02/ADD02/n14 , \u_mul/normalized_M_mul_result [13]);  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD23/ADD02/ADD02/u33  (o_mulres[13], \u_mul/normalized_M_mul_result [13], \u_mul/ADD23/ADD02/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD23/ADD02/ADD02/u34  (o_mulres[12], \u_mul/normalized_M_mul_result [12], \u_mul/ADD23/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD02/ADD02/u35  (\u_mul/ADD23/ADD02/ADD02/n20 , \u_mul/ADD23/ADD02/ADD02/n17 , \u_mul/normalized_M_mul_result [12]);  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD23/ADD02/ADD02/u36  (\u_mul/ADD23/ADD02/ADD02/n21 , \u_mul/ADD23/ADD02/ADD02/n20 , \u_mul/ADD23/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD23/ADD02/ADD02/u8  (\u_mul/ADD23/ADD02/ADD02/n0 , \u_mul/normalized_M_mul_result [12], \u_mul/ADD23/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(63)
  and \u_mul/ADD23/ADD03/ADD01/u12  (\u_mul/ADD23/ADD03/ADD01/n3 , \u_mul/normalized_M_mul_result [17], \u_mul/normalized_M_mul_result [16]);  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD23/ADD03/ADD01/u13  (\u_mul/ADD23/ADD03/ADD01/n4 , \u_mul/ADD23/ADD03/ADD01/n3 , \u_mul/ADD23/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD23/ADD03/ADD01/u17  (\u_mul/ADD23/ADD03/ADD01/n7 , \u_mul/normalized_M_mul_result [18], \u_mul/normalized_M_mul_result [17]);  // ../RTL/core/fpu_utils.v(65)
  xor \u_mul/ADD23/ADD03/ADD01/u20  (o_mulres[19], \u_mul/normalized_M_mul_result [19], \u_mul/ADD23/ADD03/ADD01/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD03/ADD01/u21  (\u_mul/ADD23/ADD03/ADD01/n10 , \u_mul/ADD23/ADD03/ADD01/n7 , \u_mul/normalized_M_mul_result [16]);  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD23/ADD03/ADD01/u22  (\u_mul/ADD23/ADD03/ADD01/n11 , \u_mul/ADD23/ADD03/ADD01/n10 , \u_mul/ADD23/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(65)
  and \u_mul/ADD23/ADD03/ADD01/u26  (\u_mul/ADD23/ADD03/ADD01/n14 , \u_mul/normalized_M_mul_result [19], \u_mul/normalized_M_mul_result [18]);  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD23/ADD03/ADD01/u29  (o_mulres[18], \u_mul/normalized_M_mul_result [18], \u_mul/ADD23/ADD03/ADD01/n4 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD03/ADD01/u30  (\u_mul/ADD23/ADD03/ADD01/n17 , \u_mul/ADD23/ADD03/ADD01/n14 , \u_mul/normalized_M_mul_result [17]);  // ../RTL/core/fpu_utils.v(66)
  xor \u_mul/ADD23/ADD03/ADD01/u33  (o_mulres[17], \u_mul/normalized_M_mul_result [17], \u_mul/ADD23/ADD03/ADD01/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD23/ADD03/ADD01/u34  (o_mulres[16], \u_mul/normalized_M_mul_result [16], \u_mul/ADD23/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD03/ADD01/u35  (\u_mul/ADD23/ADD03/ADD01/n20 , \u_mul/ADD23/ADD03/ADD01/n17 , \u_mul/normalized_M_mul_result [16]);  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD23/ADD03/ADD01/u36  (\u_mul/ADD23/ADD03/ADD01/n21 , \u_mul/ADD23/ADD03/ADD01/n20 , \u_mul/ADD23/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  and \u_mul/ADD23/ADD03/ADD01/u8  (\u_mul/ADD23/ADD03/ADD01/n0 , \u_mul/normalized_M_mul_result [16], \u_mul/ADD23/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(63)
  and \u_mul/ADD23/ADD03/ADD02/u12  (\u_mul/ADD23/ADD03/ADD02/n3 , \u_mul/normalized_M_mul_result [21], \u_mul/normalized_M_mul_result [20]);  // ../RTL/core/fpu_utils.v(64)
  and \u_mul/ADD23/ADD03/ADD02/u13  (\u_mul/ADD23/ADD03/ADD02/n4 , \u_mul/ADD23/ADD03/ADD02/n3 , \u_mul/ADD23/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(64)
  xor \u_mul/ADD23/ADD03/ADD02/u29  (o_mulres[22], \u_mul/normalized_M_mul_result [22], \u_mul/ADD23/ADD03/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD23/ADD03/ADD02/u33  (o_mulres[21], \u_mul/normalized_M_mul_result [21], \u_mul/ADD23/ADD03/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \u_mul/ADD23/ADD03/ADD02/u34  (o_mulres[20], \u_mul/normalized_M_mul_result [20], \u_mul/ADD23/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(71)
  and \u_mul/ADD23/ADD03/ADD02/u8  (\u_mul/ADD23/ADD03/ADD02/n0 , \u_mul/normalized_M_mul_result [20], \u_mul/ADD23/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(63)
  AL_MUX \u_mul/M01/u3  (
    .i0(\u_mul/mul_round1 ),
    .i1(\u_mul/mul_round2 ),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/final_product_round ));
  AL_MUX \u_mul/M02/M01/M01/u3  (
    .i0(\u_mul/M_mul_result [23]),
    .i1(\u_mul/M_mul_result [24]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [0]));
  AL_MUX \u_mul/M02/M01/M02/u3  (
    .i0(\u_mul/M_mul_result [24]),
    .i1(\u_mul/M_mul_result [25]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [1]));
  AL_MUX \u_mul/M02/M01/M03/u3  (
    .i0(\u_mul/M_mul_result [25]),
    .i1(\u_mul/M_mul_result [26]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [2]));
  AL_MUX \u_mul/M02/M01/M04/u3  (
    .i0(\u_mul/M_mul_result [26]),
    .i1(\u_mul/M_mul_result [27]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [3]));
  AL_MUX \u_mul/M02/M01/M05/u3  (
    .i0(\u_mul/M_mul_result [27]),
    .i1(\u_mul/M_mul_result [28]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [4]));
  AL_MUX \u_mul/M02/M01/M06/u3  (
    .i0(\u_mul/M_mul_result [28]),
    .i1(\u_mul/M_mul_result [29]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [5]));
  AL_MUX \u_mul/M02/M01/M07/u3  (
    .i0(\u_mul/M_mul_result [29]),
    .i1(\u_mul/M_mul_result [30]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [6]));
  AL_MUX \u_mul/M02/M01/M08/u3  (
    .i0(\u_mul/M_mul_result [30]),
    .i1(\u_mul/M_mul_result [31]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [7]));
  AL_MUX \u_mul/M02/M02/M01/u3  (
    .i0(\u_mul/M_mul_result [31]),
    .i1(\u_mul/M_mul_result [32]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [8]));
  AL_MUX \u_mul/M02/M02/M02/u3  (
    .i0(\u_mul/M_mul_result [32]),
    .i1(\u_mul/M_mul_result [33]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [9]));
  AL_MUX \u_mul/M02/M02/M03/u3  (
    .i0(\u_mul/M_mul_result [33]),
    .i1(\u_mul/M_mul_result [34]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [10]));
  AL_MUX \u_mul/M02/M02/M04/u3  (
    .i0(\u_mul/M_mul_result [34]),
    .i1(\u_mul/M_mul_result [35]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [11]));
  AL_MUX \u_mul/M02/M02/M05/u3  (
    .i0(\u_mul/M_mul_result [35]),
    .i1(\u_mul/M_mul_result [36]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [12]));
  AL_MUX \u_mul/M02/M02/M06/u3  (
    .i0(\u_mul/M_mul_result [36]),
    .i1(\u_mul/M_mul_result [37]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [13]));
  AL_MUX \u_mul/M02/M02/M07/u3  (
    .i0(\u_mul/M_mul_result [37]),
    .i1(\u_mul/M_mul_result [38]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [14]));
  AL_MUX \u_mul/M02/M02/M08/u3  (
    .i0(\u_mul/M_mul_result [38]),
    .i1(\u_mul/M_mul_result [39]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [15]));
  AL_MUX \u_mul/M02/M03/M01/u3  (
    .i0(\u_mul/M_mul_result [39]),
    .i1(\u_mul/M_mul_result [40]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [16]));
  AL_MUX \u_mul/M02/M03/M02/u3  (
    .i0(\u_mul/M_mul_result [40]),
    .i1(\u_mul/M_mul_result [41]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [17]));
  AL_MUX \u_mul/M02/M03/M03/u3  (
    .i0(\u_mul/M_mul_result [41]),
    .i1(\u_mul/M_mul_result [42]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [18]));
  AL_MUX \u_mul/M02/M03/M04/u3  (
    .i0(\u_mul/M_mul_result [42]),
    .i1(\u_mul/M_mul_result [43]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [19]));
  AL_MUX \u_mul/M02/M03/M05/u3  (
    .i0(\u_mul/M_mul_result [43]),
    .i1(\u_mul/M_mul_result [44]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [20]));
  AL_MUX \u_mul/M02/M03/M06/u3  (
    .i0(\u_mul/M_mul_result [44]),
    .i1(\u_mul/M_mul_result [45]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [21]));
  AL_MUX \u_mul/M02/M03/M07/u3  (
    .i0(\u_mul/M_mul_result [45]),
    .i1(\u_mul/M_mul_result [46]),
    .sel(\u_mul/M_mul_result [47]),
    .o(\u_mul/normalized_M_mul_result [22]));
  mult_u24_u24_o48 \u_mul/MUL01/mult0  (
    .i0({\u_mul/reduced_or_E1 ,i_op1[22:0]}),
    .i1({\u_mul/reduced_or_E1 ,i_op2[22:0]}),
    .o(\u_mul/M_mul_result ));  // ../RTL/core/fpu_utils.v(135)
  or \u_mul/RO01/u0  (\u_mul/RO01/w1 , i_op1[24], i_op1[23]);  // ../RTL/core/fpu_utils.v(14)
  or \u_mul/RO01/u1  (\u_mul/RO01/w2 , i_op1[25], \u_mul/RO01/w1 );  // ../RTL/core/fpu_utils.v(15)
  or \u_mul/RO01/u2  (\u_mul/RO01/w3 , i_op1[26], \u_mul/RO01/w2 );  // ../RTL/core/fpu_utils.v(16)
  or \u_mul/RO01/u3  (\u_mul/RO01/w4 , i_op1[27], \u_mul/RO01/w3 );  // ../RTL/core/fpu_utils.v(17)
  or \u_mul/RO01/u4  (\u_mul/RO01/w5 , i_op1[28], \u_mul/RO01/w4 );  // ../RTL/core/fpu_utils.v(18)
  or \u_mul/RO01/u5  (\u_mul/RO01/w6 , i_op1[29], \u_mul/RO01/w5 );  // ../RTL/core/fpu_utils.v(19)
  or \u_mul/RO01/u6  (\u_mul/reduced_or_E1 , i_op1[30], \u_mul/RO01/w6 );  // ../RTL/core/fpu_utils.v(20)
  or \u_mul/RO03/RO01/u0  (\u_mul/RO03/RO01/w1 , \u_mul/M_mul_result [1], \u_mul/M_mul_result [0]);  // ../RTL/core/fpu_utils.v(14)
  or \u_mul/RO03/RO01/u1  (\u_mul/RO03/RO01/w2 , \u_mul/M_mul_result [2], \u_mul/RO03/RO01/w1 );  // ../RTL/core/fpu_utils.v(15)
  or \u_mul/RO03/RO01/u2  (\u_mul/RO03/RO01/w3 , \u_mul/M_mul_result [3], \u_mul/RO03/RO01/w2 );  // ../RTL/core/fpu_utils.v(16)
  or \u_mul/RO03/RO01/u3  (\u_mul/RO03/RO01/w4 , \u_mul/M_mul_result [4], \u_mul/RO03/RO01/w3 );  // ../RTL/core/fpu_utils.v(17)
  or \u_mul/RO03/RO01/u4  (\u_mul/RO03/RO01/w5 , \u_mul/M_mul_result [5], \u_mul/RO03/RO01/w4 );  // ../RTL/core/fpu_utils.v(18)
  or \u_mul/RO03/RO01/u5  (\u_mul/RO03/RO01/w6 , \u_mul/M_mul_result [6], \u_mul/RO03/RO01/w5 );  // ../RTL/core/fpu_utils.v(19)
  or \u_mul/RO03/RO01/u6  (\u_mul/RO03/o1 , \u_mul/M_mul_result [7], \u_mul/RO03/RO01/w6 );  // ../RTL/core/fpu_utils.v(20)
  or \u_mul/RO03/RO02/u0  (\u_mul/RO03/RO02/w1 , \u_mul/M_mul_result [9], \u_mul/M_mul_result [8]);  // ../RTL/core/fpu_utils.v(14)
  or \u_mul/RO03/RO02/u1  (\u_mul/RO03/RO02/w2 , \u_mul/M_mul_result [10], \u_mul/RO03/RO02/w1 );  // ../RTL/core/fpu_utils.v(15)
  or \u_mul/RO03/RO02/u2  (\u_mul/RO03/RO02/w3 , \u_mul/M_mul_result [11], \u_mul/RO03/RO02/w2 );  // ../RTL/core/fpu_utils.v(16)
  or \u_mul/RO03/RO02/u3  (\u_mul/RO03/RO02/w4 , \u_mul/M_mul_result [12], \u_mul/RO03/RO02/w3 );  // ../RTL/core/fpu_utils.v(17)
  or \u_mul/RO03/RO02/u4  (\u_mul/RO03/RO02/w5 , \u_mul/M_mul_result [13], \u_mul/RO03/RO02/w4 );  // ../RTL/core/fpu_utils.v(18)
  or \u_mul/RO03/RO02/u5  (\u_mul/RO03/RO02/w6 , \u_mul/M_mul_result [14], \u_mul/RO03/RO02/w5 );  // ../RTL/core/fpu_utils.v(19)
  or \u_mul/RO03/RO02/u6  (\u_mul/RO03/o2 , \u_mul/M_mul_result [15], \u_mul/RO03/RO02/w6 );  // ../RTL/core/fpu_utils.v(20)
  or \u_mul/RO03/RO03/u0  (\u_mul/RO03/RO03/w1 , \u_mul/M_mul_result [17], \u_mul/M_mul_result [16]);  // ../RTL/core/fpu_utils.v(14)
  or \u_mul/RO03/RO03/u1  (\u_mul/RO03/RO03/w2 , \u_mul/M_mul_result [18], \u_mul/RO03/RO03/w1 );  // ../RTL/core/fpu_utils.v(15)
  or \u_mul/RO03/RO03/u2  (\u_mul/RO03/RO03/w3 , \u_mul/M_mul_result [19], \u_mul/RO03/RO03/w2 );  // ../RTL/core/fpu_utils.v(16)
  or \u_mul/RO03/RO03/u3  (\u_mul/RO03/RO03/w4 , \u_mul/M_mul_result [20], \u_mul/RO03/RO03/w3 );  // ../RTL/core/fpu_utils.v(17)
  or \u_mul/RO03/RO03/u4  (\u_mul/RO03/RO03/w5 , \u_mul/M_mul_result [21], \u_mul/RO03/RO03/w4 );  // ../RTL/core/fpu_utils.v(18)
  or \u_mul/RO03/RO03/u5  (\u_mul/RO03/RO03/w6 , \u_mul/M_mul_result [22], \u_mul/RO03/RO03/w5 );  // ../RTL/core/fpu_utils.v(19)
  or \u_mul/RO03/u0  (\u_mul/mul_round1 , \u_mul/RO03/RO03/w6 , \u_mul/RO03/n0 );  // ../RTL/core/fpu_utils.v(27)
  or \u_mul/RO03/u1  (\u_mul/RO03/n0 , \u_mul/RO03/o2 , \u_mul/RO03/o1 );  // ../RTL/core/fpu_utils.v(27)
  or \u_mul/RO04/RO03/u6  (\u_mul/RO04/o3 , \u_mul/M_mul_result [23], \u_mul/RO03/RO03/w6 );  // ../RTL/core/fpu_utils.v(20)
  or \u_mul/RO04/u0  (\u_mul/mul_round2 , \u_mul/RO04/o3 , \u_mul/RO03/n0 );  // ../RTL/core/fpu_utils.v(27)
  not \u_mul/sum_E[7]_inv  (\u_mul/sum_E[7]_neg , \u_mul/sum_E [7]);
  xor \u_mul/u5  (o_mulres[31], i_op1[31], i_op2[31]);  // ../RTL/core/fpu.v(266)
  add_sub u_sub (
    .n1(i_op1),
    .n2(i_op2),
    .sub(1'b1),
    .result(o_subres));  // ../RTL/core/fpu.v(33)

endmodule 

module lt_u32_u32
  (
  ci,
  i0,
  i1,
  o
  );

  input ci;
  input [31:0] i0;
  input [31:0] i1;
  output o;

  wire [31:0] diff;
  wire diff_12_18;
  wire diff_19_26;
  wire diff_27_31;
  wire diff_6_11;
  wire less_12_18;
  wire \less_12_18_inst/diff_0 ;
  wire \less_12_18_inst/diff_1 ;
  wire \less_12_18_inst/diff_2 ;
  wire \less_12_18_inst/diff_3 ;
  wire \less_12_18_inst/diff_4 ;
  wire \less_12_18_inst/diff_5 ;
  wire \less_12_18_inst/diff_6 ;
  wire \less_12_18_inst/o_0 ;
  wire \less_12_18_inst/o_1 ;
  wire \less_12_18_inst/o_2 ;
  wire \less_12_18_inst/o_3 ;
  wire \less_12_18_inst/o_4 ;
  wire \less_12_18_inst/o_5 ;
  wire less_19_26;
  wire \less_19_26_inst/diff_0 ;
  wire \less_19_26_inst/diff_1 ;
  wire \less_19_26_inst/diff_2 ;
  wire \less_19_26_inst/diff_3 ;
  wire \less_19_26_inst/diff_4 ;
  wire \less_19_26_inst/diff_5 ;
  wire \less_19_26_inst/diff_6 ;
  wire \less_19_26_inst/diff_7 ;
  wire \less_19_26_inst/o_0 ;
  wire \less_19_26_inst/o_1 ;
  wire \less_19_26_inst/o_2 ;
  wire \less_19_26_inst/o_3 ;
  wire \less_19_26_inst/o_4 ;
  wire \less_19_26_inst/o_5 ;
  wire \less_19_26_inst/o_6 ;
  wire less_27_31;
  wire \less_27_31_inst/diff_0 ;
  wire \less_27_31_inst/diff_1 ;
  wire \less_27_31_inst/diff_2 ;
  wire \less_27_31_inst/diff_3 ;
  wire \less_27_31_inst/diff_4 ;
  wire \less_27_31_inst/o_0 ;
  wire \less_27_31_inst/o_1 ;
  wire \less_27_31_inst/o_2 ;
  wire \less_27_31_inst/o_3 ;
  wire less_6_11;
  wire \less_6_11_inst/diff_0 ;
  wire \less_6_11_inst/diff_1 ;
  wire \less_6_11_inst/diff_2 ;
  wire \less_6_11_inst/diff_3 ;
  wire \less_6_11_inst/diff_4 ;
  wire \less_6_11_inst/diff_5 ;
  wire \less_6_11_inst/o_0 ;
  wire \less_6_11_inst/o_1 ;
  wire \less_6_11_inst/o_2 ;
  wire \less_6_11_inst/o_3 ;
  wire \less_6_11_inst/o_4 ;
  wire o_0;
  wire o_1;
  wire o_2;
  wire o_3;
  wire o_4;
  wire o_5;
  wire o_6;
  wire o_7;
  wire o_8;

  or any_diff_12_18 (diff_12_18, diff[12], diff[13], diff[14], diff[15], diff[16], diff[17], diff[18]);
  or any_diff_19_26 (diff_19_26, diff[19], diff[20], diff[21], diff[22], diff[23], diff[24], diff[25], diff[26]);
  or any_diff_27_31 (diff_27_31, diff[27], diff[28], diff[29], diff[30], diff[31]);
  or any_diff_6_11 (diff_6_11, diff[6], diff[7], diff[8], diff[9], diff[10], diff[11]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_12 (diff[12], i0[12], i1[12]);
  xor diff_13 (diff[13], i0[13], i1[13]);
  xor diff_14 (diff[14], i0[14], i1[14]);
  xor diff_15 (diff[15], i0[15], i1[15]);
  xor diff_16 (diff[16], i0[16], i1[16]);
  xor diff_17 (diff[17], i0[17], i1[17]);
  xor diff_18 (diff[18], i0[18], i1[18]);
  xor diff_19 (diff[19], i0[19], i1[19]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_20 (diff[20], i0[20], i1[20]);
  xor diff_21 (diff[21], i0[21], i1[21]);
  xor diff_22 (diff[22], i0[22], i1[22]);
  xor diff_23 (diff[23], i0[23], i1[23]);
  xor diff_24 (diff[24], i0[24], i1[24]);
  xor diff_25 (diff[25], i0[25], i1[25]);
  xor diff_26 (diff[26], i0[26], i1[26]);
  xor diff_27 (diff[27], i0[27], i1[27]);
  xor diff_28 (diff[28], i0[28], i1[28]);
  xor diff_29 (diff[29], i0[29], i1[29]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_30 (diff[30], i0[30], i1[30]);
  xor diff_31 (diff[31], i0[31], i1[31]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);
  AL_MUX \less_12_18_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[12]),
    .sel(\less_12_18_inst/diff_0 ),
    .o(\less_12_18_inst/o_0 ));
  AL_MUX \less_12_18_inst/mux_1  (
    .i0(\less_12_18_inst/o_0 ),
    .i1(i1[13]),
    .sel(\less_12_18_inst/diff_1 ),
    .o(\less_12_18_inst/o_1 ));
  AL_MUX \less_12_18_inst/mux_2  (
    .i0(\less_12_18_inst/o_1 ),
    .i1(i1[14]),
    .sel(\less_12_18_inst/diff_2 ),
    .o(\less_12_18_inst/o_2 ));
  AL_MUX \less_12_18_inst/mux_3  (
    .i0(\less_12_18_inst/o_2 ),
    .i1(i1[15]),
    .sel(\less_12_18_inst/diff_3 ),
    .o(\less_12_18_inst/o_3 ));
  AL_MUX \less_12_18_inst/mux_4  (
    .i0(\less_12_18_inst/o_3 ),
    .i1(i1[16]),
    .sel(\less_12_18_inst/diff_4 ),
    .o(\less_12_18_inst/o_4 ));
  AL_MUX \less_12_18_inst/mux_5  (
    .i0(\less_12_18_inst/o_4 ),
    .i1(i1[17]),
    .sel(\less_12_18_inst/diff_5 ),
    .o(\less_12_18_inst/o_5 ));
  AL_MUX \less_12_18_inst/mux_6  (
    .i0(\less_12_18_inst/o_5 ),
    .i1(i1[18]),
    .sel(\less_12_18_inst/diff_6 ),
    .o(less_12_18));
  xor \less_12_18_inst/xor_0  (\less_12_18_inst/diff_0 , i0[12], i1[12]);
  xor \less_12_18_inst/xor_1  (\less_12_18_inst/diff_1 , i0[13], i1[13]);
  xor \less_12_18_inst/xor_2  (\less_12_18_inst/diff_2 , i0[14], i1[14]);
  xor \less_12_18_inst/xor_3  (\less_12_18_inst/diff_3 , i0[15], i1[15]);
  xor \less_12_18_inst/xor_4  (\less_12_18_inst/diff_4 , i0[16], i1[16]);
  xor \less_12_18_inst/xor_5  (\less_12_18_inst/diff_5 , i0[17], i1[17]);
  xor \less_12_18_inst/xor_6  (\less_12_18_inst/diff_6 , i0[18], i1[18]);
  AL_MUX \less_19_26_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[19]),
    .sel(\less_19_26_inst/diff_0 ),
    .o(\less_19_26_inst/o_0 ));
  AL_MUX \less_19_26_inst/mux_1  (
    .i0(\less_19_26_inst/o_0 ),
    .i1(i1[20]),
    .sel(\less_19_26_inst/diff_1 ),
    .o(\less_19_26_inst/o_1 ));
  AL_MUX \less_19_26_inst/mux_2  (
    .i0(\less_19_26_inst/o_1 ),
    .i1(i1[21]),
    .sel(\less_19_26_inst/diff_2 ),
    .o(\less_19_26_inst/o_2 ));
  AL_MUX \less_19_26_inst/mux_3  (
    .i0(\less_19_26_inst/o_2 ),
    .i1(i1[22]),
    .sel(\less_19_26_inst/diff_3 ),
    .o(\less_19_26_inst/o_3 ));
  AL_MUX \less_19_26_inst/mux_4  (
    .i0(\less_19_26_inst/o_3 ),
    .i1(i1[23]),
    .sel(\less_19_26_inst/diff_4 ),
    .o(\less_19_26_inst/o_4 ));
  AL_MUX \less_19_26_inst/mux_5  (
    .i0(\less_19_26_inst/o_4 ),
    .i1(i1[24]),
    .sel(\less_19_26_inst/diff_5 ),
    .o(\less_19_26_inst/o_5 ));
  AL_MUX \less_19_26_inst/mux_6  (
    .i0(\less_19_26_inst/o_5 ),
    .i1(i1[25]),
    .sel(\less_19_26_inst/diff_6 ),
    .o(\less_19_26_inst/o_6 ));
  AL_MUX \less_19_26_inst/mux_7  (
    .i0(\less_19_26_inst/o_6 ),
    .i1(i1[26]),
    .sel(\less_19_26_inst/diff_7 ),
    .o(less_19_26));
  xor \less_19_26_inst/xor_0  (\less_19_26_inst/diff_0 , i0[19], i1[19]);
  xor \less_19_26_inst/xor_1  (\less_19_26_inst/diff_1 , i0[20], i1[20]);
  xor \less_19_26_inst/xor_2  (\less_19_26_inst/diff_2 , i0[21], i1[21]);
  xor \less_19_26_inst/xor_3  (\less_19_26_inst/diff_3 , i0[22], i1[22]);
  xor \less_19_26_inst/xor_4  (\less_19_26_inst/diff_4 , i0[23], i1[23]);
  xor \less_19_26_inst/xor_5  (\less_19_26_inst/diff_5 , i0[24], i1[24]);
  xor \less_19_26_inst/xor_6  (\less_19_26_inst/diff_6 , i0[25], i1[25]);
  xor \less_19_26_inst/xor_7  (\less_19_26_inst/diff_7 , i0[26], i1[26]);
  AL_MUX \less_27_31_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[27]),
    .sel(\less_27_31_inst/diff_0 ),
    .o(\less_27_31_inst/o_0 ));
  AL_MUX \less_27_31_inst/mux_1  (
    .i0(\less_27_31_inst/o_0 ),
    .i1(i1[28]),
    .sel(\less_27_31_inst/diff_1 ),
    .o(\less_27_31_inst/o_1 ));
  AL_MUX \less_27_31_inst/mux_2  (
    .i0(\less_27_31_inst/o_1 ),
    .i1(i1[29]),
    .sel(\less_27_31_inst/diff_2 ),
    .o(\less_27_31_inst/o_2 ));
  AL_MUX \less_27_31_inst/mux_3  (
    .i0(\less_27_31_inst/o_2 ),
    .i1(i1[30]),
    .sel(\less_27_31_inst/diff_3 ),
    .o(\less_27_31_inst/o_3 ));
  AL_MUX \less_27_31_inst/mux_4  (
    .i0(\less_27_31_inst/o_3 ),
    .i1(i1[31]),
    .sel(\less_27_31_inst/diff_4 ),
    .o(less_27_31));
  xor \less_27_31_inst/xor_0  (\less_27_31_inst/diff_0 , i0[27], i1[27]);
  xor \less_27_31_inst/xor_1  (\less_27_31_inst/diff_1 , i0[28], i1[28]);
  xor \less_27_31_inst/xor_2  (\less_27_31_inst/diff_2 , i0[29], i1[29]);
  xor \less_27_31_inst/xor_3  (\less_27_31_inst/diff_3 , i0[30], i1[30]);
  xor \less_27_31_inst/xor_4  (\less_27_31_inst/diff_4 , i0[31], i1[31]);
  AL_MUX \less_6_11_inst/mux_0  (
    .i0(1'b0),
    .i1(i1[6]),
    .sel(\less_6_11_inst/diff_0 ),
    .o(\less_6_11_inst/o_0 ));
  AL_MUX \less_6_11_inst/mux_1  (
    .i0(\less_6_11_inst/o_0 ),
    .i1(i1[7]),
    .sel(\less_6_11_inst/diff_1 ),
    .o(\less_6_11_inst/o_1 ));
  AL_MUX \less_6_11_inst/mux_2  (
    .i0(\less_6_11_inst/o_1 ),
    .i1(i1[8]),
    .sel(\less_6_11_inst/diff_2 ),
    .o(\less_6_11_inst/o_2 ));
  AL_MUX \less_6_11_inst/mux_3  (
    .i0(\less_6_11_inst/o_2 ),
    .i1(i1[9]),
    .sel(\less_6_11_inst/diff_3 ),
    .o(\less_6_11_inst/o_3 ));
  AL_MUX \less_6_11_inst/mux_4  (
    .i0(\less_6_11_inst/o_3 ),
    .i1(i1[10]),
    .sel(\less_6_11_inst/diff_4 ),
    .o(\less_6_11_inst/o_4 ));
  AL_MUX \less_6_11_inst/mux_5  (
    .i0(\less_6_11_inst/o_4 ),
    .i1(i1[11]),
    .sel(\less_6_11_inst/diff_5 ),
    .o(less_6_11));
  xor \less_6_11_inst/xor_0  (\less_6_11_inst/diff_0 , i0[6], i1[6]);
  xor \less_6_11_inst/xor_1  (\less_6_11_inst/diff_1 , i0[7], i1[7]);
  xor \less_6_11_inst/xor_2  (\less_6_11_inst/diff_2 , i0[8], i1[8]);
  xor \less_6_11_inst/xor_3  (\less_6_11_inst/diff_3 , i0[9], i1[9]);
  xor \less_6_11_inst/xor_4  (\less_6_11_inst/diff_4 , i0[10], i1[10]);
  xor \less_6_11_inst/xor_5  (\less_6_11_inst/diff_5 , i0[11], i1[11]);
  AL_MUX mux_0 (
    .i0(ci),
    .i1(i1[0]),
    .sel(diff[0]),
    .o(o_0));
  AL_MUX mux_1 (
    .i0(o_0),
    .i1(i1[1]),
    .sel(diff[1]),
    .o(o_1));
  AL_MUX mux_2 (
    .i0(o_1),
    .i1(i1[2]),
    .sel(diff[2]),
    .o(o_2));
  AL_MUX mux_3 (
    .i0(o_2),
    .i1(i1[3]),
    .sel(diff[3]),
    .o(o_3));
  AL_MUX mux_4 (
    .i0(o_3),
    .i1(i1[4]),
    .sel(diff[4]),
    .o(o_4));
  AL_MUX mux_5 (
    .i0(o_4),
    .i1(i1[5]),
    .sel(diff[5]),
    .o(o_5));
  AL_MUX mux_6 (
    .i0(o_5),
    .i1(less_6_11),
    .sel(diff_6_11),
    .o(o_6));
  AL_MUX mux_7 (
    .i0(o_6),
    .i1(less_12_18),
    .sel(diff_12_18),
    .o(o_7));
  AL_MUX mux_8 (
    .i0(o_7),
    .i1(less_19_26),
    .sel(diff_19_26),
    .o(o_8));
  AL_MUX mux_9 (
    .i0(o_8),
    .i1(less_27_31),
    .sel(diff_27_31),
    .o(o));

endmodule 

module add_pu32_mu32_o32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output [31:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a23;
  wire net_a24;
  wire net_a25;
  wire net_a26;
  wire net_a27;
  wire net_a28;
  wire net_a29;
  wire net_a3;
  wire net_a30;
  wire net_a31;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb10;
  wire net_nb11;
  wire net_nb12;
  wire net_nb13;
  wire net_nb14;
  wire net_nb15;
  wire net_nb16;
  wire net_nb17;
  wire net_nb18;
  wire net_nb19;
  wire net_nb2;
  wire net_nb20;
  wire net_nb21;
  wire net_nb22;
  wire net_nb23;
  wire net_nb24;
  wire net_nb25;
  wire net_nb26;
  wire net_nb27;
  wire net_nb28;
  wire net_nb29;
  wire net_nb3;
  wire net_nb30;
  wire net_nb31;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a31 = i0[31];
  assign net_a30 = i0[30];
  assign net_a29 = i0[29];
  assign net_a28 = i0[28];
  assign net_a27 = i0[27];
  assign net_a26 = i0[26];
  assign net_a25 = i0[25];
  assign net_a24 = i0[24];
  assign net_a23 = i0[23];
  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b31 = i1[31];
  assign net_b30 = i1[30];
  assign net_b29 = i1[29];
  assign net_b28 = i1[28];
  assign net_b27 = i1[27];
  assign net_b26 = i1[26];
  assign net_b25 = i1[25];
  assign net_b24 = i1[24];
  assign net_b23 = i1[23];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_nb10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_nb11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_nb12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_nb13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_nb14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_nb15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_nb16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_nb17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_nb18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_nb19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_nb20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_nb21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_nb22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(net_a23),
    .b(net_nb23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(net_a24),
    .b(net_nb24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(net_a25),
    .b(net_nb25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(net_a26),
    .b(net_nb26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(net_a27),
    .b(net_nb27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(net_a28),
    .b(net_nb28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(net_a29),
    .b(net_nb29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(net_a30),
    .b(net_nb30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(net_a31),
    .b(net_nb31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b10 (net_nb10, net_b10);
  not inv_b11 (net_nb11, net_b11);
  not inv_b12 (net_nb12, net_b12);
  not inv_b13 (net_nb13, net_b13);
  not inv_b14 (net_nb14, net_b14);
  not inv_b15 (net_nb15, net_b15);
  not inv_b16 (net_nb16, net_b16);
  not inv_b17 (net_nb17, net_b17);
  not inv_b18 (net_nb18, net_b18);
  not inv_b19 (net_nb19, net_b19);
  not inv_b2 (net_nb2, net_b2);
  not inv_b20 (net_nb20, net_b20);
  not inv_b21 (net_nb21, net_b21);
  not inv_b22 (net_nb22, net_b22);
  not inv_b23 (net_nb23, net_b23);
  not inv_b24 (net_nb24, net_b24);
  not inv_b25 (net_nb25, net_b25);
  not inv_b26 (net_nb26, net_b26);
  not inv_b27 (net_nb27, net_b27);
  not inv_b28 (net_nb28, net_b28);
  not inv_b29 (net_nb29, net_b29);
  not inv_b3 (net_nb3, net_b3);
  not inv_b30 (net_nb30, net_b30);
  not inv_b31 (net_nb31, net_b31);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);

endmodule 

module eq_w32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output o;

  wire or_or_or_or_or_xor_i_o;
  wire \or_or_or_or_xor_i0[0_o ;
  wire \or_or_or_or_xor_i0[1_o ;
  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_or_xor_i0[16]__o ;
  wire \or_or_or_xor_i0[24]__o ;
  wire \or_or_or_xor_i0[8]_i_o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[12]_i1[_o ;
  wire \or_or_xor_i0[16]_i1[_o ;
  wire \or_or_xor_i0[20]_i1[_o ;
  wire \or_or_xor_i0[24]_i1[_o ;
  wire \or_or_xor_i0[28]_i1[_o ;
  wire \or_or_xor_i0[4]_i1[4_o ;
  wire \or_or_xor_i0[8]_i1[8_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[10]_i1[10]_o ;
  wire \or_xor_i0[12]_i1[12]_o ;
  wire \or_xor_i0[14]_i1[14]_o ;
  wire \or_xor_i0[16]_i1[16]_o ;
  wire \or_xor_i0[18]_i1[18]_o ;
  wire \or_xor_i0[20]_i1[20]_o ;
  wire \or_xor_i0[22]_i1[22]_o ;
  wire \or_xor_i0[24]_i1[24]_o ;
  wire \or_xor_i0[26]_i1[26]_o ;
  wire \or_xor_i0[28]_i1[28]_o ;
  wire \or_xor_i0[2]_i1[2]_o_o ;
  wire \or_xor_i0[30]_i1[30]_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[8]_i1[8]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[12]_i1[12]_o ;
  wire \xor_i0[13]_i1[13]_o ;
  wire \xor_i0[14]_i1[14]_o ;
  wire \xor_i0[15]_i1[15]_o ;
  wire \xor_i0[16]_i1[16]_o ;
  wire \xor_i0[17]_i1[17]_o ;
  wire \xor_i0[18]_i1[18]_o ;
  wire \xor_i0[19]_i1[19]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[20]_i1[20]_o ;
  wire \xor_i0[21]_i1[21]_o ;
  wire \xor_i0[22]_i1[22]_o ;
  wire \xor_i0[23]_i1[23]_o ;
  wire \xor_i0[24]_i1[24]_o ;
  wire \xor_i0[25]_i1[25]_o ;
  wire \xor_i0[26]_i1[26]_o ;
  wire \xor_i0[27]_i1[27]_o ;
  wire \xor_i0[28]_i1[28]_o ;
  wire \xor_i0[29]_i1[29]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[30]_i1[30]_o ;
  wire \xor_i0[31]_i1[31]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, or_or_or_or_or_xor_i_o);
  or or_or_or_or_or_xor_i (or_or_or_or_or_xor_i_o, \or_or_or_or_xor_i0[0_o , \or_or_or_or_xor_i0[1_o );
  or \or_or_or_or_xor_i0[0  (\or_or_or_or_xor_i0[0_o , \or_or_or_xor_i0[0]_i_o , \or_or_or_xor_i0[8]_i_o );
  or \or_or_or_or_xor_i0[1  (\or_or_or_or_xor_i0[1_o , \or_or_or_xor_i0[16]__o , \or_or_or_xor_i0[24]__o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[4]_i1[4_o );
  or \or_or_or_xor_i0[16]_  (\or_or_or_xor_i0[16]__o , \or_or_xor_i0[16]_i1[_o , \or_or_xor_i0[20]_i1[_o );
  or \or_or_or_xor_i0[24]_  (\or_or_or_xor_i0[24]__o , \or_or_xor_i0[24]_i1[_o , \or_or_xor_i0[28]_i1[_o );
  or \or_or_or_xor_i0[8]_i  (\or_or_or_xor_i0[8]_i_o , \or_or_xor_i0[8]_i1[8_o , \or_or_xor_i0[12]_i1[_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[2]_i1[2]_o_o );
  or \or_or_xor_i0[12]_i1[  (\or_or_xor_i0[12]_i1[_o , \or_xor_i0[12]_i1[12]_o , \or_xor_i0[14]_i1[14]_o );
  or \or_or_xor_i0[16]_i1[  (\or_or_xor_i0[16]_i1[_o , \or_xor_i0[16]_i1[16]_o , \or_xor_i0[18]_i1[18]_o );
  or \or_or_xor_i0[20]_i1[  (\or_or_xor_i0[20]_i1[_o , \or_xor_i0[20]_i1[20]_o , \or_xor_i0[22]_i1[22]_o );
  or \or_or_xor_i0[24]_i1[  (\or_or_xor_i0[24]_i1[_o , \or_xor_i0[24]_i1[24]_o , \or_xor_i0[26]_i1[26]_o );
  or \or_or_xor_i0[28]_i1[  (\or_or_xor_i0[28]_i1[_o , \or_xor_i0[28]_i1[28]_o , \or_xor_i0[30]_i1[30]_o );
  or \or_or_xor_i0[4]_i1[4  (\or_or_xor_i0[4]_i1[4_o , \or_xor_i0[4]_i1[4]_o_o , \or_xor_i0[6]_i1[6]_o_o );
  or \or_or_xor_i0[8]_i1[8  (\or_or_xor_i0[8]_i1[8_o , \or_xor_i0[8]_i1[8]_o_o , \or_xor_i0[10]_i1[10]_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  or \or_xor_i0[10]_i1[10]  (\or_xor_i0[10]_i1[10]_o , \xor_i0[10]_i1[10]_o , \xor_i0[11]_i1[11]_o );
  or \or_xor_i0[12]_i1[12]  (\or_xor_i0[12]_i1[12]_o , \xor_i0[12]_i1[12]_o , \xor_i0[13]_i1[13]_o );
  or \or_xor_i0[14]_i1[14]  (\or_xor_i0[14]_i1[14]_o , \xor_i0[14]_i1[14]_o , \xor_i0[15]_i1[15]_o );
  or \or_xor_i0[16]_i1[16]  (\or_xor_i0[16]_i1[16]_o , \xor_i0[16]_i1[16]_o , \xor_i0[17]_i1[17]_o );
  or \or_xor_i0[18]_i1[18]  (\or_xor_i0[18]_i1[18]_o , \xor_i0[18]_i1[18]_o , \xor_i0[19]_i1[19]_o );
  or \or_xor_i0[20]_i1[20]  (\or_xor_i0[20]_i1[20]_o , \xor_i0[20]_i1[20]_o , \xor_i0[21]_i1[21]_o );
  or \or_xor_i0[22]_i1[22]  (\or_xor_i0[22]_i1[22]_o , \xor_i0[22]_i1[22]_o , \xor_i0[23]_i1[23]_o );
  or \or_xor_i0[24]_i1[24]  (\or_xor_i0[24]_i1[24]_o , \xor_i0[24]_i1[24]_o , \xor_i0[25]_i1[25]_o );
  or \or_xor_i0[26]_i1[26]  (\or_xor_i0[26]_i1[26]_o , \xor_i0[26]_i1[26]_o , \xor_i0[27]_i1[27]_o );
  or \or_xor_i0[28]_i1[28]  (\or_xor_i0[28]_i1[28]_o , \xor_i0[28]_i1[28]_o , \xor_i0[29]_i1[29]_o );
  or \or_xor_i0[2]_i1[2]_o  (\or_xor_i0[2]_i1[2]_o_o , \xor_i0[2]_i1[2]_o , \xor_i0[3]_i1[3]_o );
  or \or_xor_i0[30]_i1[30]  (\or_xor_i0[30]_i1[30]_o , \xor_i0[30]_i1[30]_o , \xor_i0[31]_i1[31]_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \xor_i0[7]_i1[7]_o );
  or \or_xor_i0[8]_i1[8]_o  (\or_xor_i0[8]_i1[8]_o_o , \xor_i0[8]_i1[8]_o , \xor_i0[9]_i1[9]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (\xor_i0[12]_i1[12]_o , i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (\xor_i0[13]_i1[13]_o , i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (\xor_i0[14]_i1[14]_o , i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (\xor_i0[15]_i1[15]_o , i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (\xor_i0[16]_i1[16]_o , i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (\xor_i0[17]_i1[17]_o , i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (\xor_i0[18]_i1[18]_o , i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (\xor_i0[19]_i1[19]_o , i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (\xor_i0[20]_i1[20]_o , i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (\xor_i0[21]_i1[21]_o , i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (\xor_i0[22]_i1[22]_o , i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (\xor_i0[23]_i1[23]_o , i0[23], i1[23]);
  xor \xor_i0[24]_i1[24]  (\xor_i0[24]_i1[24]_o , i0[24], i1[24]);
  xor \xor_i0[25]_i1[25]  (\xor_i0[25]_i1[25]_o , i0[25], i1[25]);
  xor \xor_i0[26]_i1[26]  (\xor_i0[26]_i1[26]_o , i0[26], i1[26]);
  xor \xor_i0[27]_i1[27]  (\xor_i0[27]_i1[27]_o , i0[27], i1[27]);
  xor \xor_i0[28]_i1[28]  (\xor_i0[28]_i1[28]_o , i0[28], i1[28]);
  xor \xor_i0[29]_i1[29]  (\xor_i0[29]_i1[29]_o , i0[29], i1[29]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[30]_i1[30]  (\xor_i0[30]_i1[30]_o , i0[30], i1[30]);
  xor \xor_i0[31]_i1[31]  (\xor_i0[31]_i1[31]_o , i0[31], i1[31]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module ne_w32
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output o;

  wire [31:0] diff;

  or any_diff (o, diff[0], diff[1], diff[2], diff[3], diff[4], diff[5], diff[6], diff[7], diff[8], diff[9], diff[10], diff[11], diff[12], diff[13], diff[14], diff[15], diff[16], diff[17], diff[18], diff[19], diff[20], diff[21], diff[22], diff[23], diff[24], diff[25], diff[26], diff[27], diff[28], diff[29], diff[30], diff[31]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);
  xor diff_10 (diff[10], i0[10], i1[10]);
  xor diff_11 (diff[11], i0[11], i1[11]);
  xor diff_12 (diff[12], i0[12], i1[12]);
  xor diff_13 (diff[13], i0[13], i1[13]);
  xor diff_14 (diff[14], i0[14], i1[14]);
  xor diff_15 (diff[15], i0[15], i1[15]);
  xor diff_16 (diff[16], i0[16], i1[16]);
  xor diff_17 (diff[17], i0[17], i1[17]);
  xor diff_18 (diff[18], i0[18], i1[18]);
  xor diff_19 (diff[19], i0[19], i1[19]);
  xor diff_2 (diff[2], i0[2], i1[2]);
  xor diff_20 (diff[20], i0[20], i1[20]);
  xor diff_21 (diff[21], i0[21], i1[21]);
  xor diff_22 (diff[22], i0[22], i1[22]);
  xor diff_23 (diff[23], i0[23], i1[23]);
  xor diff_24 (diff[24], i0[24], i1[24]);
  xor diff_25 (diff[25], i0[25], i1[25]);
  xor diff_26 (diff[26], i0[26], i1[26]);
  xor diff_27 (diff[27], i0[27], i1[27]);
  xor diff_28 (diff[28], i0[28], i1[28]);
  xor diff_29 (diff[29], i0[29], i1[29]);
  xor diff_3 (diff[3], i0[3], i1[3]);
  xor diff_30 (diff[30], i0[30], i1[30]);
  xor diff_31 (diff[31], i0[31], i1[31]);
  xor diff_4 (diff[4], i0[4], i1[4]);
  xor diff_5 (diff[5], i0[5], i1[5]);
  xor diff_6 (diff[6], i0[6], i1[6]);
  xor diff_7 (diff[7], i0[7], i1[7]);
  xor diff_8 (diff[8], i0[8], i1[8]);
  xor diff_9 (diff[9], i0[9], i1[9]);

endmodule 

module eq_w2
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output o;

  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[1]_i1[1]_o ;

  not none_diff (o, \or_xor_i0[0]_i1[0]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \xor_i0[1]_i1[1]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);

endmodule 

module ne_w2
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output o;

  wire [1:0] diff;

  or any_diff (o, diff[0], diff[1]);
  xor diff_0 (diff[0], i0[0], i1[0]);
  xor diff_1 (diff[1], i0[1], i1[1]);

endmodule 

module add_pu2_mu2_o3
  (
  i0,
  i1,
  o
  );

  input [1:0] i0;
  input [1:0] i1;
  output [2:0] o;

  wire net_a0;
  wire net_a1;
  wire net_b0;
  wire net_b1;
  wire net_cout0;
  wire net_cout1;
  wire net_nb0;
  wire net_nb1;
  wire net_ncout;
  wire net_sum0;
  wire net_sum1;

  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[2] = net_ncout;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_cout (net_ncout, net_cout1);

endmodule 

module EXU_MDU  // ../RTL/core/exu_mdu.v(14)
  (
  i_clk,
  i_decinfo_grp,
  i_flush,
  i_mdu_op1,
  i_mdu_op2,
  i_mdu_rdidx,
  i_mdu_rdwen,
  i_mduinfo,
  i_rstn,
  i_vld,
  o_mdu_rdidx,
  o_mdu_rdwdata,
  o_mdu_rdwen,
  o_will_rdidx,
  o_will_rdwen,
  o_working
  );

  input i_clk;  // ../RTL/core/exu_mdu.v(15)
  input [5:0] i_decinfo_grp;  // ../RTL/core/exu_mdu.v(21)
  input i_flush;  // ../RTL/core/exu_mdu.v(19)
  input [31:0] i_mdu_op1;  // ../RTL/core/exu_mdu.v(25)
  input [31:0] i_mdu_op2;  // ../RTL/core/exu_mdu.v(26)
  input [4:0] i_mdu_rdidx;  // ../RTL/core/exu_mdu.v(24)
  input i_mdu_rdwen;  // ../RTL/core/exu_mdu.v(23)
  input [9:0] i_mduinfo;  // ../RTL/core/exu_mdu.v(22)
  input i_rstn;  // ../RTL/core/exu_mdu.v(16)
  input i_vld;  // ../RTL/core/exu_mdu.v(18)
  output [4:0] o_mdu_rdidx;  // ../RTL/core/exu_mdu.v(36)
  output [31:0] o_mdu_rdwdata;  // ../RTL/core/exu_mdu.v(37)
  output o_mdu_rdwen;  // ../RTL/core/exu_mdu.v(35)
  output [4:0] o_will_rdidx;  // ../RTL/core/exu_mdu.v(32)
  output o_will_rdwen;  // ../RTL/core/exu_mdu.v(31)
  output o_working;  // ../RTL/core/exu_mdu.v(29)

  wire [7:0] cnt;  // ../RTL/core/exu_mdu.v(85)
  wire [31:0] div_signed_quo;  // ../RTL/core/exu_mdu.v(125)
  wire [31:0] div_signed_rem;  // ../RTL/core/exu_mdu.v(126)
  wire [31:0] div_unsigned_quo;  // ../RTL/core/exu_mdu.v(140)
  wire [31:0] div_unsigned_rem;  // ../RTL/core/exu_mdu.v(141)
  wire [9:0] mduinfo;  // ../RTL/core/exu_mdu.v(50)
  wire [63:0] mul_ss;  // ../RTL/core/exu_mdu.v(90)
  wire [63:0] mul_su;  // ../RTL/core/exu_mdu.v(92)
  wire [63:0] mul_uu;  // ../RTL/core/exu_mdu.v(91)
  wire [7:0] n19;
  wire [7:0] n22;
  wire [7:0] n25;
  wire [7:0] n29;
  wire [31:0] n34;
  wire [31:0] n35;
  wire [31:0] n37;
  wire [31:0] n38;
  wire [31:0] n39;
  wire [31:0] n40;
  wire [31:0] n41;
  wire [31:0] n42;
  wire [31:0] n43;
  wire [31:0] n44;
  wire [31:0] n45;
  wire [31:0] op1;  // ../RTL/core/exu_mdu.v(87)
  wire [31:0] op2;  // ../RTL/core/exu_mdu.v(88)
  wire [5:0] \u_DIV_SIGNED/al_00000256AA0CE7C0 ;  // al_ip/div_signed_gate.v(42)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA0CEB40 ;  // al_ip/div_signed_gate.v(58)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA0CF470 ;  // al_ip/div_signed_gate.v(57)
  wire [62:0] \u_DIV_SIGNED/al_00000256AA0D0BA0 ;  // al_ip/div_signed_gate.v(43)
  wire [5:0] \u_DIV_SIGNED/al_00000256AA0D29D0 ;  // al_ip/div_signed_gate.v(48)
  wire [5:0] \u_DIV_SIGNED/al_00000256AA0D38B0 ;  // al_ip/div_signed_gate.v(53)
  wire [62:0] \u_DIV_SIGNED/al_00000256AA0D5590 ;  // al_ip/div_signed_gate.v(54)
  wire [62:0] \u_DIV_SIGNED/al_00000256AA0D7970 ;  // al_ip/div_signed_gate.v(55)
  wire [62:0] \u_DIV_SIGNED/al_00000256AA0D80E0 ;  // al_ip/div_signed_gate.v(56)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA3FF0F0 ;  // al_ip/div_signed_gate.v(44)
  wire [62:0] \u_DIV_SIGNED/al_00000256AA400D60 ;  // al_ip/div_signed_gate.v(45)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA402C70 ;  // al_ip/div_signed_gate.v(47)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA403450 ;  // al_ip/div_signed_gate.v(46)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA4072E0 ;  // al_ip/div_signed_gate.v(49)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA4073C0 ;  // al_ip/div_signed_gate.v(50)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA4098F0 ;  // al_ip/div_signed_gate.v(52)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA40B170 ;  // al_ip/div_signed_gate.v(51)
  wire [5:0] \u_DIV_UNSIGNED/al_00000286E57DB3B0 ;  // al_ip/div_unsigned_gate.v(42)
  wire [31:0] \u_DIV_UNSIGNED/al_00000286E57DBF10 ;  // al_ip/div_unsigned_gate.v(50)
  wire [31:0] \u_DIV_UNSIGNED/al_00000286E57DC290 ;  // al_ip/div_unsigned_gate.v(49)
  wire [62:0] \u_DIV_UNSIGNED/al_00000286E57DE2F0 ;  // al_ip/div_unsigned_gate.v(43)
  wire [62:0] \u_DIV_UNSIGNED/al_00000286E57DEE50 ;  // al_ip/div_unsigned_gate.v(46)
  wire [5:0] \u_DIV_UNSIGNED/al_00000286E57E03C0 ;  // al_ip/div_unsigned_gate.v(44)
  wire [5:0] \u_DIV_UNSIGNED/al_00000286E57E04A0 ;  // al_ip/div_unsigned_gate.v(45)
  wire [62:0] \u_DIV_UNSIGNED/al_00000286E57E1690 ;  // al_ip/div_unsigned_gate.v(47)
  wire [31:0] \u_DIV_UNSIGNED/al_00000286E57E4870 ;  // al_ip/div_unsigned_gate.v(48)
  wire div_finish;  // ../RTL/core/exu_mdu.v(153)
  wire div_signed_finish;  // ../RTL/core/exu_mdu.v(124)
  wire div_signed_start;  // ../RTL/core/exu_mdu.v(127)
  wire div_unsigned_finish;  // ../RTL/core/exu_mdu.v(139)
  wire div_unsigned_start;  // ../RTL/core/exu_mdu.v(142)
  wire i_flush_neg;
  wire mdu_finish;  // ../RTL/core/exu_mdu.v(41)
  wire mdu_finish_neg;
  wire mdu_vld;  // ../RTL/core/exu_mdu.v(47)
  wire mul_finish;  // ../RTL/core/exu_mdu.v(89)
  wire mul_start;  // ../RTL/core/exu_mdu.v(93)
  wire mul_start_neg;
  wire mul_vld;  // ../RTL/core/exu_mdu.v(86)
  wire mux10_b0_sel_is_2_o;
  wire mux2_b0_sel_is_2_o;
  wire n0;
  wire n1;
  wire n10;
  wire n14;
  wire n15;
  wire n16;
  wire n18;
  wire n20;
  wire n24;
  wire n26;
  wire n3;
  wire n30;
  wire n33;
  wire n36;
  wire n4;
  wire n5;
  wire n6;
  wire n8;
  wire rem_op1_sym;  // ../RTL/core/exu_mdu.v(45)
  wire u28_sel_is_3_o;
  wire u30_sel_is_2_o;
  wire u9_sel_is_0_o;
  wire \u_DIV_SIGNED/al_00000256AA3DB060 ;  // al_ip/div_signed_gate.v(128)
  wire \u_DIV_SIGNED/al_00000256AA3DB110 ;  // al_ip/div_signed_gate.v(103)
  wire \u_DIV_SIGNED/al_00000256AA3DB320 ;  // al_ip/div_signed_gate.v(120)
  wire \u_DIV_SIGNED/al_00000256AA3DB3D0 ;  // al_ip/div_signed_gate.v(127)
  wire \u_DIV_SIGNED/al_00000256AA3DB480 ;  // al_ip/div_signed_gate.v(129)
  wire \u_DIV_SIGNED/al_00000256AA3DB5E0 ;  // al_ip/div_signed_gate.v(116)
  wire \u_DIV_SIGNED/al_00000256AA3DB7F0 ;  // al_ip/div_signed_gate.v(196)
  wire \u_DIV_SIGNED/al_00000256AA3DBC10 ;  // al_ip/div_signed_gate.v(106)
  wire \u_DIV_SIGNED/al_00000256AA3DBCC0 ;  // al_ip/div_signed_gate.v(117)
  wire \u_DIV_SIGNED/al_00000256AA3DBD70 ;  // al_ip/div_signed_gate.v(102)
  wire \u_DIV_SIGNED/al_00000256AA3DBF80 ;  // al_ip/div_signed_gate.v(113)
  wire \u_DIV_SIGNED/al_00000256AA3DC030 ;  // al_ip/div_signed_gate.v(263)
  wire \u_DIV_SIGNED/al_00000256AA3DC3A0 ;  // al_ip/div_signed_gate.v(104)
  wire \u_DIV_SIGNED/al_00000256AA3DC450 ;  // al_ip/div_signed_gate.v(107)
  wire \u_DIV_SIGNED/al_00000256AA3DC500 ;  // al_ip/div_signed_gate.v(115)
  wire \u_DIV_SIGNED/al_00000256AA3DC5B0 ;  // al_ip/div_signed_gate.v(264)
  wire \u_DIV_SIGNED/al_00000256AA3DC870 ;  // al_ip/div_signed_gate.v(105)
  wire \u_DIV_SIGNED/al_00000256AA3DC9D0 ;  // al_ip/div_signed_gate.v(122)
  wire \u_DIV_SIGNED/al_00000256AA3DCA80 ;  // al_ip/div_signed_gate.v(126)
  wire \u_DIV_SIGNED/al_00000256AA3DCB30 ;  // al_ip/div_signed_gate.v(108)
  wire \u_DIV_SIGNED/al_00000256AA3DCC90 ;  // al_ip/div_signed_gate.v(114)
  wire \u_DIV_SIGNED/al_00000256AA3DCD40 ;  // al_ip/div_signed_gate.v(121)
  wire \u_DIV_SIGNED/al_00000256AA3DD210 ;  // al_ip/div_signed_gate.v(100)
  wire \u_DIV_SIGNED/al_00000256AA3DD2C0 ;  // al_ip/div_signed_gate.v(101)
  wire \u_DIV_SIGNED/al_00000256AA3DD370 ;  // al_ip/div_signed_gate.v(110)
  wire \u_DIV_SIGNED/al_00000256AA3DD420 ;  // al_ip/div_signed_gate.v(111)
  wire \u_DIV_SIGNED/al_00000256AA3DD4D0 ;  // al_ip/div_signed_gate.v(112)
  wire \u_DIV_SIGNED/al_00000256AA3DD580 ;  // al_ip/div_signed_gate.v(118)
  wire \u_DIV_SIGNED/al_00000256AA3DD840 ;  // al_ip/div_signed_gate.v(123)
  wire \u_DIV_SIGNED/al_00000256AA3DD8F0 ;  // al_ip/div_signed_gate.v(124)
  wire \u_DIV_SIGNED/al_00000256AA3DD9A0 ;  // al_ip/div_signed_gate.v(261)
  wire \u_DIV_SIGNED/al_00000256AA3DDA50 ;  // al_ip/div_signed_gate.v(109)
  wire \u_DIV_SIGNED/al_00000256AA3DDB00 ;  // al_ip/div_signed_gate.v(125)
  wire \u_DIV_SIGNED/al_00000256AA3DDBB0 ;  // al_ip/div_signed_gate.v(119)
  wire \u_DIV_SIGNED/al_00000256AA3DEA20 ;  // al_ip/div_signed_gate.v(131)
  wire \u_DIV_SIGNED/al_00000256AA3DEB80 ;  // al_ip/div_signed_gate.v(130)
  wire \u_DIV_SIGNED/al_00000256AA3E0300 ;  // al_ip/div_signed_gate.v(163)
  wire \u_DIV_SIGNED/al_00000256AA421080 ;  // al_ip/div_signed_gate.v(77)
  wire \u_DIV_SIGNED/al_00000256AA421130 ;  // al_ip/div_signed_gate.v(79)
  wire \u_DIV_SIGNED/al_00000256AA421290 ;  // al_ip/div_signed_gate.v(89)
  wire \u_DIV_SIGNED/al_00000256AA421550 ;  // al_ip/div_signed_gate.v(82)
  wire \u_DIV_SIGNED/al_00000256AA421600 ;  // al_ip/div_signed_gate.v(93)
  wire \u_DIV_SIGNED/al_00000256AA4216B0 ;  // al_ip/div_signed_gate.v(90)
  wire \u_DIV_SIGNED/al_00000256AA421760 ;  // al_ip/div_signed_gate.v(72)
  wire \u_DIV_SIGNED/al_00000256AA421810 ;  // al_ip/div_signed_gate.v(81)
  wire \u_DIV_SIGNED/al_00000256AA4218C0 ;  // al_ip/div_signed_gate.v(91)
  wire \u_DIV_SIGNED/al_00000256AA421B80 ;  // al_ip/div_signed_gate.v(94)
  wire \u_DIV_SIGNED/al_00000256AA421C30 ;  // al_ip/div_signed_gate.v(95)
  wire \u_DIV_SIGNED/al_00000256AA421CE0 ;  // al_ip/div_signed_gate.v(88)
  wire \u_DIV_SIGNED/al_00000256AA421EF0 ;  // al_ip/div_signed_gate.v(78)
  wire \u_DIV_SIGNED/al_00000256AA4221B0 ;  // al_ip/div_signed_gate.v(83)
  wire \u_DIV_SIGNED/al_00000256AA422310 ;  // al_ip/div_signed_gate.v(86)
  wire \u_DIV_SIGNED/al_00000256AA4223C0 ;  // al_ip/div_signed_gate.v(96)
  wire \u_DIV_SIGNED/al_00000256AA422470 ;  // al_ip/div_signed_gate.v(97)
  wire \u_DIV_SIGNED/al_00000256AA422520 ;  // al_ip/div_signed_gate.v(85)
  wire \u_DIV_SIGNED/al_00000256AA4225D0 ;  // al_ip/div_signed_gate.v(98)
  wire \u_DIV_SIGNED/al_00000256AA422680 ;  // al_ip/div_signed_gate.v(262)
  wire \u_DIV_SIGNED/al_00000256AA422940 ;  // al_ip/div_signed_gate.v(75)
  wire \u_DIV_SIGNED/al_00000256AA422E10 ;  // al_ip/div_signed_gate.v(73)
  wire \u_DIV_SIGNED/al_00000256AA422EC0 ;  // al_ip/div_signed_gate.v(92)
  wire \u_DIV_SIGNED/al_00000256AA423020 ;  // al_ip/div_signed_gate.v(74)
  wire \u_DIV_SIGNED/al_00000256AA423230 ;  // al_ip/div_signed_gate.v(87)
  wire \u_DIV_SIGNED/al_00000256AA4232E0 ;  // al_ip/div_signed_gate.v(99)
  wire \u_DIV_SIGNED/al_00000256AA423390 ;  // al_ip/div_signed_gate.v(71)
  wire \u_DIV_SIGNED/al_00000256AA423650 ;  // al_ip/div_signed_gate.v(80)
  wire \u_DIV_SIGNED/al_00000256AA423700 ;  // al_ip/div_signed_gate.v(84)
  wire \u_DIV_SIGNED/al_00000256AA4237B0 ;  // al_ip/div_signed_gate.v(76)
  wire \u_DIV_SIGNED/al_00000256AA423910 ;  // al_ip/div_signed_gate.v(68)
  wire \u_DIV_SIGNED/al_00000256AA423B20 ;  // al_ip/div_signed_gate.v(69)
  wire \u_DIV_SIGNED/al_00000256AA423BD0 ;  // al_ip/div_signed_gate.v(70)
  wire \u_DIV_SIGNED/al_00000256AA443080 ;  // al_ip/div_signed_gate.v(140)
  wire \u_DIV_SIGNED/al_00000256AA443130 ;  // al_ip/div_signed_gate.v(150)
  wire \u_DIV_SIGNED/al_00000256AA4436B0 ;  // al_ip/div_signed_gate.v(135)
  wire \u_DIV_SIGNED/al_00000256AA443760 ;  // al_ip/div_signed_gate.v(141)
  wire \u_DIV_SIGNED/al_00000256AA443810 ;  // al_ip/div_signed_gate.v(143)
  wire \u_DIV_SIGNED/al_00000256AA443C30 ;  // al_ip/div_signed_gate.v(132)
  wire \u_DIV_SIGNED/al_00000256AA443CE0 ;  // al_ip/div_signed_gate.v(137)
  wire \u_DIV_SIGNED/al_00000256AA443E40 ;  // al_ip/div_signed_gate.v(139)
  wire \u_DIV_SIGNED/al_00000256AA443EF0 ;  // al_ip/div_signed_gate.v(142)
  wire \u_DIV_SIGNED/al_00000256AA444050 ;  // al_ip/div_signed_gate.v(144)
  wire \u_DIV_SIGNED/al_00000256AA444100 ;  // al_ip/div_signed_gate.v(148)
  wire \u_DIV_SIGNED/al_00000256AA444260 ;  // al_ip/div_signed_gate.v(154)
  wire \u_DIV_SIGNED/al_00000256AA444310 ;  // al_ip/div_signed_gate.v(156)
  wire \u_DIV_SIGNED/al_00000256AA444520 ;  // al_ip/div_signed_gate.v(136)
  wire \u_DIV_SIGNED/al_00000256AA4445D0 ;  // al_ip/div_signed_gate.v(157)
  wire \u_DIV_SIGNED/al_00000256AA444680 ;  // al_ip/div_signed_gate.v(146)
  wire \u_DIV_SIGNED/al_00000256AA444730 ;  // al_ip/div_signed_gate.v(158)
  wire \u_DIV_SIGNED/al_00000256AA444940 ;  // al_ip/div_signed_gate.v(159)
  wire \u_DIV_SIGNED/al_00000256AA444B50 ;  // al_ip/div_signed_gate.v(152)
  wire \u_DIV_SIGNED/al_00000256AA444CB0 ;  // al_ip/div_signed_gate.v(155)
  wire \u_DIV_SIGNED/al_00000256AA444D60 ;  // al_ip/div_signed_gate.v(160)
  wire \u_DIV_SIGNED/al_00000256AA444E10 ;  // al_ip/div_signed_gate.v(161)
  wire \u_DIV_SIGNED/al_00000256AA444EC0 ;  // al_ip/div_signed_gate.v(162)
  wire \u_DIV_SIGNED/al_00000256AA445020 ;  // al_ip/div_signed_gate.v(151)
  wire \u_DIV_SIGNED/al_00000256AA445230 ;  // al_ip/div_signed_gate.v(133)
  wire \u_DIV_SIGNED/al_00000256AA4452E0 ;  // al_ip/div_signed_gate.v(147)
  wire \u_DIV_SIGNED/al_00000256AA445390 ;  // al_ip/div_signed_gate.v(149)
  wire \u_DIV_SIGNED/al_00000256AA445860 ;  // al_ip/div_signed_gate.v(134)
  wire \u_DIV_SIGNED/al_00000256AA445910 ;  // al_ip/div_signed_gate.v(138)
  wire \u_DIV_SIGNED/al_00000256AA4459C0 ;  // al_ip/div_signed_gate.v(145)
  wire \u_DIV_SIGNED/al_00000256AA445B20 ;  // al_ip/div_signed_gate.v(153)
  wire \u_DIV_SIGNED/al_00000256AA653100 ;  // al_ip/div_signed_gate.v(64)
  wire \u_DIV_SIGNED/al_00000256AA6537E0 ;  // al_ip/div_signed_gate.v(62)
  wire \u_DIV_SIGNED/al_00000256AA653890 ;  // al_ip/div_signed_gate.v(65)
  wire \u_DIV_SIGNED/al_00000256AA6539F0 ;  // al_ip/div_signed_gate.v(66)
  wire \u_DIV_SIGNED/al_00000256AA653E10 ;  // al_ip/div_signed_gate.v(67)
  wire \u_DIV_SIGNED/al_00000256AA6547B0 ;  // al_ip/div_signed_gate.v(63)
  wire \u_DIV_SIGNED/al_00000256AA88A8D0 ;  // al_ip/div_signed_gate.v(202)
  wire \u_DIV_SIGNED/al_00000256AA88A980 ;  // al_ip/div_signed_gate.v(260)
  wire \u_DIV_SIGNED/al_00000256AA88AA30 ;  // al_ip/div_signed_gate.v(199)
  wire \u_DIV_SIGNED/al_00000256AA88AAE0 ;  // al_ip/div_signed_gate.v(259)
  wire \u_DIV_SIGNED/al_00000256AA88AB90 ;  // al_ip/div_signed_gate.v(205)
  wire \u_DIV_SIGNED/al_00000256AA88AC40 ;  // al_ip/div_signed_gate.v(187)
  wire \u_DIV_SIGNED/al_00000256AA88ACF0 ;  // al_ip/div_signed_gate.v(190)
  wire \u_DIV_SIGNED/al_00000256AA88ADA0 ;  // al_ip/div_signed_gate.v(242)
  wire \u_DIV_SIGNED/al_00000256AA88AE50 ;  // al_ip/div_signed_gate.v(253)
  wire \u_DIV_SIGNED/al_00000256AA88AF00 ;  // al_ip/div_signed_gate.v(195)
  wire \u_DIV_SIGNED/al_00000256AA88AFB0 ;  // al_ip/div_signed_gate.v(203)
  wire \u_DIV_SIGNED/al_00000256AA88B060 ;  // al_ip/div_signed_gate.v(186)
  wire \u_DIV_SIGNED/al_00000256AA88B110 ;  // al_ip/div_signed_gate.v(206)
  wire \u_DIV_SIGNED/al_00000256AA88B1C0 ;  // al_ip/div_signed_gate.v(176)
  wire \u_DIV_SIGNED/al_00000256AA88B270 ;  // al_ip/div_signed_gate.v(191)
  wire \u_DIV_SIGNED/al_00000256AA88B320 ;  // al_ip/div_signed_gate.v(179)
  wire \u_DIV_SIGNED/al_00000256AA88B3D0 ;  // al_ip/div_signed_gate.v(207)
  wire \u_DIV_SIGNED/al_00000256AA88B480 ;  // al_ip/div_signed_gate.v(208)
  wire \u_DIV_SIGNED/al_00000256AA88B530 ;  // al_ip/div_signed_gate.v(193)
  wire \u_DIV_SIGNED/al_00000256AA88B5E0 ;  // al_ip/div_signed_gate.v(177)
  wire \u_DIV_SIGNED/al_00000256AA88B690 ;  // al_ip/div_signed_gate.v(197)
  wire \u_DIV_SIGNED/al_00000256AA88B740 ;  // al_ip/div_signed_gate.v(210)
  wire \u_DIV_SIGNED/al_00000256AA88B7F0 ;  // al_ip/div_signed_gate.v(212)
  wire \u_DIV_SIGNED/al_00000256AA88B8A0 ;  // al_ip/div_signed_gate.v(172)
  wire \u_DIV_SIGNED/al_00000256AA88B950 ;  // al_ip/div_signed_gate.v(184)
  wire \u_DIV_SIGNED/al_00000256AA88BA00 ;  // al_ip/div_signed_gate.v(211)
  wire \u_DIV_SIGNED/al_00000256AA88BAB0 ;  // al_ip/div_signed_gate.v(213)
  wire \u_DIV_SIGNED/al_00000256AA88BB60 ;  // al_ip/div_signed_gate.v(214)
  wire \u_DIV_SIGNED/al_00000256AA88BC10 ;  // al_ip/div_signed_gate.v(215)
  wire \u_DIV_SIGNED/al_00000256AA88BCC0 ;  // al_ip/div_signed_gate.v(200)
  wire \u_DIV_SIGNED/al_00000256AA88BD70 ;  // al_ip/div_signed_gate.v(216)
  wire \u_DIV_SIGNED/al_00000256AA88BE20 ;  // al_ip/div_signed_gate.v(217)
  wire \u_DIV_SIGNED/al_00000256AA88BED0 ;  // al_ip/div_signed_gate.v(173)
  wire \u_DIV_SIGNED/al_00000256AA88BF80 ;  // al_ip/div_signed_gate.v(218)
  wire \u_DIV_SIGNED/al_00000256AA88C030 ;  // al_ip/div_signed_gate.v(219)
  wire \u_DIV_SIGNED/al_00000256AA88C0E0 ;  // al_ip/div_signed_gate.v(221)
  wire \u_DIV_SIGNED/al_00000256AA88C190 ;  // al_ip/div_signed_gate.v(165)
  wire \u_DIV_SIGNED/al_00000256AA88C240 ;  // al_ip/div_signed_gate.v(169)
  wire \u_DIV_SIGNED/al_00000256AA88C2F0 ;  // al_ip/div_signed_gate.v(174)
  wire \u_DIV_SIGNED/al_00000256AA88C3A0 ;  // al_ip/div_signed_gate.v(204)
  wire \u_DIV_SIGNED/al_00000256AA88C450 ;  // al_ip/div_signed_gate.v(220)
  wire \u_DIV_SIGNED/al_00000256AA88C500 ;  // al_ip/div_signed_gate.v(198)
  wire \u_DIV_SIGNED/al_00000256AA88C5B0 ;  // al_ip/div_signed_gate.v(180)
  wire \u_DIV_SIGNED/al_00000256AA88C660 ;  // al_ip/div_signed_gate.v(171)
  wire \u_DIV_SIGNED/al_00000256AA88C710 ;  // al_ip/div_signed_gate.v(189)
  wire \u_DIV_SIGNED/al_00000256AA88C870 ;  // al_ip/div_signed_gate.v(168)
  wire \u_DIV_SIGNED/al_00000256AA88C920 ;  // al_ip/div_signed_gate.v(166)
  wire \u_DIV_SIGNED/al_00000256AA88C9D0 ;  // al_ip/div_signed_gate.v(170)
  wire \u_DIV_SIGNED/al_00000256AA88CA80 ;  // al_ip/div_signed_gate.v(182)
  wire \u_DIV_SIGNED/al_00000256AA88CB30 ;  // al_ip/div_signed_gate.v(188)
  wire \u_DIV_SIGNED/al_00000256AA88CBE0 ;  // al_ip/div_signed_gate.v(178)
  wire \u_DIV_SIGNED/al_00000256AA88CC90 ;  // al_ip/div_signed_gate.v(192)
  wire \u_DIV_SIGNED/al_00000256AA88CD40 ;  // al_ip/div_signed_gate.v(194)
  wire \u_DIV_SIGNED/al_00000256AA88CDF0 ;  // al_ip/div_signed_gate.v(209)
  wire \u_DIV_SIGNED/al_00000256AA88CEA0 ;  // al_ip/div_signed_gate.v(175)
  wire \u_DIV_SIGNED/al_00000256AA88CF50 ;  // al_ip/div_signed_gate.v(185)
  wire \u_DIV_SIGNED/al_00000256AA88D000 ;  // al_ip/div_signed_gate.v(231)
  wire \u_DIV_SIGNED/al_00000256AA88D0B0 ;  // al_ip/div_signed_gate.v(258)
  wire \u_DIV_SIGNED/al_00000256AA88D160 ;  // al_ip/div_signed_gate.v(201)
  wire \u_DIV_SIGNED/al_00000256AA88D210 ;  // al_ip/div_signed_gate.v(164)
  wire \u_DIV_SIGNED/al_00000256AA88D2C0 ;  // al_ip/div_signed_gate.v(183)
  wire \u_DIV_SIGNED/al_00000256AA88D370 ;  // al_ip/div_signed_gate.v(181)
  wire \u_DIV_SIGNED/al_00000256AA88D420 ;  // al_ip/div_signed_gate.v(167)
  wire \u_DIV_SIGNED/al_00000256AA88D630 ;  // al_ip/div_signed_gate.v(257)
  wire \u_DIV_SIGNED/al_00000256AA88DA50 ;  // al_ip/div_signed_gate.v(254)
  wire \u_DIV_SIGNED/al_00000256AA88DB00 ;  // al_ip/div_signed_gate.v(224)
  wire \u_DIV_SIGNED/al_00000256AA88DD10 ;  // al_ip/div_signed_gate.v(227)
  wire \u_DIV_SIGNED/al_00000256AA88DE70 ;  // al_ip/div_signed_gate.v(237)
  wire \u_DIV_SIGNED/al_00000256AA88DF20 ;  // al_ip/div_signed_gate.v(241)
  wire \u_DIV_SIGNED/al_00000256AA88DFD0 ;  // al_ip/div_signed_gate.v(248)
  wire \u_DIV_SIGNED/al_00000256AA88E130 ;  // al_ip/div_signed_gate.v(235)
  wire \u_DIV_SIGNED/al_00000256AA88E1E0 ;  // al_ip/div_signed_gate.v(239)
  wire \u_DIV_SIGNED/al_00000256AA88E290 ;  // al_ip/div_signed_gate.v(247)
  wire \u_DIV_SIGNED/al_00000256AA88E340 ;  // al_ip/div_signed_gate.v(252)
  wire \u_DIV_SIGNED/al_00000256AA88E810 ;  // al_ip/div_signed_gate.v(251)
  wire \u_DIV_SIGNED/al_00000256AA88E970 ;  // al_ip/div_signed_gate.v(229)
  wire \u_DIV_SIGNED/al_00000256AA88EA20 ;  // al_ip/div_signed_gate.v(256)
  wire \u_DIV_SIGNED/al_00000256AA88EC30 ;  // al_ip/div_signed_gate.v(225)
  wire \u_DIV_SIGNED/al_00000256AA88ECE0 ;  // al_ip/div_signed_gate.v(245)
  wire \u_DIV_SIGNED/al_00000256AA88EE40 ;  // al_ip/div_signed_gate.v(226)
  wire \u_DIV_SIGNED/al_00000256AA88F260 ;  // al_ip/div_signed_gate.v(236)
  wire \u_DIV_SIGNED/al_00000256AA88F310 ;  // al_ip/div_signed_gate.v(240)
  wire \u_DIV_SIGNED/al_00000256AA88F3C0 ;  // al_ip/div_signed_gate.v(230)
  wire \u_DIV_SIGNED/al_00000256AA88F470 ;  // al_ip/div_signed_gate.v(228)
  wire \u_DIV_SIGNED/al_00000256AA88F520 ;  // al_ip/div_signed_gate.v(244)
  wire \u_DIV_SIGNED/al_00000256AA88F5D0 ;  // al_ip/div_signed_gate.v(223)
  wire \u_DIV_SIGNED/al_00000256AA88F680 ;  // al_ip/div_signed_gate.v(250)
  wire \u_DIV_SIGNED/al_00000256AA88F730 ;  // al_ip/div_signed_gate.v(255)
  wire \u_DIV_SIGNED/al_00000256AA88F890 ;  // al_ip/div_signed_gate.v(233)
  wire \u_DIV_SIGNED/al_00000256AA88F940 ;  // al_ip/div_signed_gate.v(243)
  wire \u_DIV_SIGNED/al_00000256AA88F9F0 ;  // al_ip/div_signed_gate.v(246)
  wire \u_DIV_SIGNED/al_00000256AA88FAA0 ;  // al_ip/div_signed_gate.v(234)
  wire \u_DIV_SIGNED/al_00000256AA88FB50 ;  // al_ip/div_signed_gate.v(238)
  wire \u_DIV_SIGNED/al_00000256AA88FC00 ;  // al_ip/div_signed_gate.v(222)
  wire \u_DIV_SIGNED/al_00000256AA88FCB0 ;  // al_ip/div_signed_gate.v(249)
  wire \u_DIV_SIGNED/al_00000256AA88FD60 ;  // al_ip/div_signed_gate.v(232)
  wire \u_DIV_SIGNED/al_00000256AA893670 ;  // al_ip/div_signed_gate.v(59)
  wire \u_DIV_SIGNED/al_00000256AA8940C0 ;  // al_ip/div_signed_gate.v(61)
  wire \u_DIV_SIGNED/al_00000256AA895350 ;  // al_ip/div_signed_gate.v(60)
  wire \u_DIV_SIGNED/al_00000256AA898580 ;  // al_ip/div_signed_gate.v(265)
  wire \u_DIV_SIGNED/al_00000256AA898630 ;  // al_ip/div_signed_gate.v(285)
  wire \u_DIV_SIGNED/al_00000256AA8986E0 ;  // al_ip/div_signed_gate.v(287)
  wire \u_DIV_SIGNED/al_00000256AA8988F0 ;  // al_ip/div_signed_gate.v(274)
  wire \u_DIV_SIGNED/al_00000256AA898D10 ;  // al_ip/div_signed_gate.v(283)
  wire \u_DIV_SIGNED/al_00000256AA898DC0 ;  // al_ip/div_signed_gate.v(276)
  wire \u_DIV_SIGNED/al_00000256AA898E70 ;  // al_ip/div_signed_gate.v(281)
  wire \u_DIV_SIGNED/al_00000256AA898F20 ;  // al_ip/div_signed_gate.v(284)
  wire \u_DIV_SIGNED/al_00000256AA898FD0 ;  // al_ip/div_signed_gate.v(288)
  wire \u_DIV_SIGNED/al_00000256AA899080 ;  // al_ip/div_signed_gate.v(296)
  wire \u_DIV_SIGNED/al_00000256AA899130 ;  // al_ip/div_signed_gate.v(272)
  wire \u_DIV_SIGNED/al_00000256AA899290 ;  // al_ip/div_signed_gate.v(268)
  wire \u_DIV_SIGNED/al_00000256AA899340 ;  // al_ip/div_signed_gate.v(282)
  wire \u_DIV_SIGNED/al_00000256AA8993F0 ;  // al_ip/div_signed_gate.v(271)
  wire \u_DIV_SIGNED/al_00000256AA8994A0 ;  // al_ip/div_signed_gate.v(275)
  wire \u_DIV_SIGNED/al_00000256AA899550 ;  // al_ip/div_signed_gate.v(286)
  wire \u_DIV_SIGNED/al_00000256AA899600 ;  // al_ip/div_signed_gate.v(289)
  wire \u_DIV_SIGNED/al_00000256AA8996B0 ;  // al_ip/div_signed_gate.v(270)
  wire \u_DIV_SIGNED/al_00000256AA899760 ;  // al_ip/div_signed_gate.v(277)
  wire \u_DIV_SIGNED/al_00000256AA899810 ;  // al_ip/div_signed_gate.v(290)
  wire \u_DIV_SIGNED/al_00000256AA8998C0 ;  // al_ip/div_signed_gate.v(291)
  wire \u_DIV_SIGNED/al_00000256AA899970 ;  // al_ip/div_signed_gate.v(269)
  wire \u_DIV_SIGNED/al_00000256AA899EF0 ;  // al_ip/div_signed_gate.v(267)
  wire \u_DIV_SIGNED/al_00000256AA89A260 ;  // al_ip/div_signed_gate.v(279)
  wire \u_DIV_SIGNED/al_00000256AA89A470 ;  // al_ip/div_signed_gate.v(292)
  wire \u_DIV_SIGNED/al_00000256AA89A520 ;  // al_ip/div_signed_gate.v(273)
  wire \u_DIV_SIGNED/al_00000256AA89A5D0 ;  // al_ip/div_signed_gate.v(266)
  wire \u_DIV_SIGNED/al_00000256AA89A680 ;  // al_ip/div_signed_gate.v(293)
  wire \u_DIV_SIGNED/al_00000256AA89A730 ;  // al_ip/div_signed_gate.v(295)
  wire \u_DIV_SIGNED/al_00000256AA89AC00 ;  // al_ip/div_signed_gate.v(278)
  wire \u_DIV_SIGNED/al_00000256AA89ACB0 ;  // al_ip/div_signed_gate.v(280)
  wire \u_DIV_SIGNED/al_00000256AA89AEC0 ;  // al_ip/div_signed_gate.v(294)
  wire \u_DIV_UNSIGNED/al_00000286E447F1F0 ;  // al_ip/div_unsigned_gate.v(125)
  wire \u_DIV_UNSIGNED/al_00000286E447F350 ;  // al_ip/div_unsigned_gate.v(126)
  wire \u_DIV_UNSIGNED/al_00000286E447F6C0 ;  // al_ip/div_unsigned_gate.v(131)
  wire \u_DIV_UNSIGNED/al_00000286E447FC40 ;  // al_ip/div_unsigned_gate.v(133)
  wire \u_DIV_UNSIGNED/al_00000286E447FCF0 ;  // al_ip/div_unsigned_gate.v(135)
  wire \u_DIV_UNSIGNED/al_00000286E447FDA0 ;  // al_ip/div_unsigned_gate.v(137)
  wire \u_DIV_UNSIGNED/al_00000286E447FE50 ;  // al_ip/div_unsigned_gate.v(139)
  wire \u_DIV_UNSIGNED/al_00000286E447FF00 ;  // al_ip/div_unsigned_gate.v(143)
  wire \u_DIV_UNSIGNED/al_00000286E4480110 ;  // al_ip/div_unsigned_gate.v(144)
  wire \u_DIV_UNSIGNED/al_00000286E4480270 ;  // al_ip/div_unsigned_gate.v(146)
  wire \u_DIV_UNSIGNED/al_00000286E44803D0 ;  // al_ip/div_unsigned_gate.v(138)
  wire \u_DIV_UNSIGNED/al_00000286E4480480 ;  // al_ip/div_unsigned_gate.v(136)
  wire \u_DIV_UNSIGNED/al_00000286E4480530 ;  // al_ip/div_unsigned_gate.v(145)
  wire \u_DIV_UNSIGNED/al_00000286E44805E0 ;  // al_ip/div_unsigned_gate.v(148)
  wire \u_DIV_UNSIGNED/al_00000286E44808A0 ;  // al_ip/div_unsigned_gate.v(132)
  wire \u_DIV_UNSIGNED/al_00000286E4480A00 ;  // al_ip/div_unsigned_gate.v(142)
  wire \u_DIV_UNSIGNED/al_00000286E4480AB0 ;  // al_ip/div_unsigned_gate.v(149)
  wire \u_DIV_UNSIGNED/al_00000286E4480B60 ;  // al_ip/div_unsigned_gate.v(150)
  wire \u_DIV_UNSIGNED/al_00000286E4480CC0 ;  // al_ip/div_unsigned_gate.v(141)
  wire \u_DIV_UNSIGNED/al_00000286E4481030 ;  // al_ip/div_unsigned_gate.v(129)
  wire \u_DIV_UNSIGNED/al_00000286E44810E0 ;  // al_ip/div_unsigned_gate.v(130)
  wire \u_DIV_UNSIGNED/al_00000286E44812F0 ;  // al_ip/div_unsigned_gate.v(147)
  wire \u_DIV_UNSIGNED/al_00000286E4481500 ;  // al_ip/div_unsigned_gate.v(151)
  wire \u_DIV_UNSIGNED/al_00000286E44815B0 ;  // al_ip/div_unsigned_gate.v(152)
  wire \u_DIV_UNSIGNED/al_00000286E4481660 ;  // al_ip/div_unsigned_gate.v(153)
  wire \u_DIV_UNSIGNED/al_00000286E4481710 ;  // al_ip/div_unsigned_gate.v(154)
  wire \u_DIV_UNSIGNED/al_00000286E44817C0 ;  // al_ip/div_unsigned_gate.v(155)
  wire \u_DIV_UNSIGNED/al_00000286E4481920 ;  // al_ip/div_unsigned_gate.v(140)
  wire \u_DIV_UNSIGNED/al_00000286E44819D0 ;  // al_ip/div_unsigned_gate.v(134)
  wire \u_DIV_UNSIGNED/al_00000286E4481B30 ;  // al_ip/div_unsigned_gate.v(128)
  wire \u_DIV_UNSIGNED/al_00000286E4481BE0 ;  // al_ip/div_unsigned_gate.v(127)
  wire \u_DIV_UNSIGNED/al_00000286E44833F0 ;  // al_ip/div_unsigned_gate.v(156)
  wire \u_DIV_UNSIGNED/al_00000286E4688A90 ;  // al_ip/div_unsigned_gate.v(51)
  wire \u_DIV_UNSIGNED/al_00000286E468A980 ;  // al_ip/div_unsigned_gate.v(52)
  wire \u_DIV_UNSIGNED/al_00000286E4A23D20 ;  // al_ip/div_unsigned_gate.v(83)
  wire \u_DIV_UNSIGNED/al_00000286E4A23DD0 ;  // al_ip/div_unsigned_gate.v(60)
  wire \u_DIV_UNSIGNED/al_00000286E4A23E80 ;  // al_ip/div_unsigned_gate.v(66)
  wire \u_DIV_UNSIGNED/al_00000286E4A23F30 ;  // al_ip/div_unsigned_gate.v(65)
  wire \u_DIV_UNSIGNED/al_00000286E4A23FE0 ;  // al_ip/div_unsigned_gate.v(67)
  wire \u_DIV_UNSIGNED/al_00000286E4A24090 ;  // al_ip/div_unsigned_gate.v(68)
  wire \u_DIV_UNSIGNED/al_00000286E4A24560 ;  // al_ip/div_unsigned_gate.v(54)
  wire \u_DIV_UNSIGNED/al_00000286E4A24610 ;  // al_ip/div_unsigned_gate.v(62)
  wire \u_DIV_UNSIGNED/al_00000286E4A24770 ;  // al_ip/div_unsigned_gate.v(116)
  wire \u_DIV_UNSIGNED/al_00000286E4A24820 ;  // al_ip/div_unsigned_gate.v(123)
  wire \u_DIV_UNSIGNED/al_00000286E4A248D0 ;  // al_ip/div_unsigned_gate.v(64)
  wire \u_DIV_UNSIGNED/al_00000286E4A24A30 ;  // al_ip/div_unsigned_gate.v(58)
  wire \u_DIV_UNSIGNED/al_00000286E4A24AE0 ;  // al_ip/div_unsigned_gate.v(72)
  wire \u_DIV_UNSIGNED/al_00000286E4A24DA0 ;  // al_ip/div_unsigned_gate.v(55)
  wire \u_DIV_UNSIGNED/al_00000286E4A24E50 ;  // al_ip/div_unsigned_gate.v(56)
  wire \u_DIV_UNSIGNED/al_00000286E4A24FB0 ;  // al_ip/div_unsigned_gate.v(121)
  wire \u_DIV_UNSIGNED/al_00000286E4A25060 ;  // al_ip/div_unsigned_gate.v(69)
  wire \u_DIV_UNSIGNED/al_00000286E4A25110 ;  // al_ip/div_unsigned_gate.v(73)
  wire \u_DIV_UNSIGNED/al_00000286E4A251C0 ;  // al_ip/div_unsigned_gate.v(75)
  wire \u_DIV_UNSIGNED/al_00000286E4A25270 ;  // al_ip/div_unsigned_gate.v(77)
  wire \u_DIV_UNSIGNED/al_00000286E4A253D0 ;  // al_ip/div_unsigned_gate.v(53)
  wire \u_DIV_UNSIGNED/al_00000286E4A25530 ;  // al_ip/div_unsigned_gate.v(61)
  wire \u_DIV_UNSIGNED/al_00000286E4A25690 ;  // al_ip/div_unsigned_gate.v(105)
  wire \u_DIV_UNSIGNED/al_00000286E4A25740 ;  // al_ip/div_unsigned_gate.v(63)
  wire \u_DIV_UNSIGNED/al_00000286E4A257F0 ;  // al_ip/div_unsigned_gate.v(57)
  wire \u_DIV_UNSIGNED/al_00000286E4A258A0 ;  // al_ip/div_unsigned_gate.v(71)
  wire \u_DIV_UNSIGNED/al_00000286E4A25950 ;  // al_ip/div_unsigned_gate.v(74)
  wire \u_DIV_UNSIGNED/al_00000286E4A25A00 ;  // al_ip/div_unsigned_gate.v(78)
  wire \u_DIV_UNSIGNED/al_00000286E4A25B60 ;  // al_ip/div_unsigned_gate.v(79)
  wire \u_DIV_UNSIGNED/al_00000286E4A25C10 ;  // al_ip/div_unsigned_gate.v(80)
  wire \u_DIV_UNSIGNED/al_00000286E4A25CC0 ;  // al_ip/div_unsigned_gate.v(81)
  wire \u_DIV_UNSIGNED/al_00000286E4A25D70 ;  // al_ip/div_unsigned_gate.v(94)
  wire \u_DIV_UNSIGNED/al_00000286E4A25ED0 ;  // al_ip/div_unsigned_gate.v(76)
  wire \u_DIV_UNSIGNED/al_00000286E4A25F80 ;  // al_ip/div_unsigned_gate.v(82)
  wire \u_DIV_UNSIGNED/al_00000286E4A26030 ;  // al_ip/div_unsigned_gate.v(84)
  wire \u_DIV_UNSIGNED/al_00000286E4A260E0 ;  // al_ip/div_unsigned_gate.v(85)
  wire \u_DIV_UNSIGNED/al_00000286E4A262F0 ;  // al_ip/div_unsigned_gate.v(122)
  wire \u_DIV_UNSIGNED/al_00000286E4A263A0 ;  // al_ip/div_unsigned_gate.v(70)
  wire \u_DIV_UNSIGNED/al_00000286E4A26870 ;  // al_ip/div_unsigned_gate.v(86)
  wire \u_DIV_UNSIGNED/al_00000286E4A26920 ;  // al_ip/div_unsigned_gate.v(88)
  wire \u_DIV_UNSIGNED/al_00000286E4A269D0 ;  // al_ip/div_unsigned_gate.v(90)
  wire \u_DIV_UNSIGNED/al_00000286E4A26A80 ;  // al_ip/div_unsigned_gate.v(91)
  wire \u_DIV_UNSIGNED/al_00000286E4A26B30 ;  // al_ip/div_unsigned_gate.v(108)
  wire \u_DIV_UNSIGNED/al_00000286E4A26BE0 ;  // al_ip/div_unsigned_gate.v(109)
  wire \u_DIV_UNSIGNED/al_00000286E4A26C90 ;  // al_ip/div_unsigned_gate.v(112)
  wire \u_DIV_UNSIGNED/al_00000286E4A26D40 ;  // al_ip/div_unsigned_gate.v(120)
  wire \u_DIV_UNSIGNED/al_00000286E4A26F50 ;  // al_ip/div_unsigned_gate.v(93)
  wire \u_DIV_UNSIGNED/al_00000286E4A270B0 ;  // al_ip/div_unsigned_gate.v(98)
  wire \u_DIV_UNSIGNED/al_00000286E4A27160 ;  // al_ip/div_unsigned_gate.v(118)
  wire \u_DIV_UNSIGNED/al_00000286E4A27210 ;  // al_ip/div_unsigned_gate.v(104)
  wire \u_DIV_UNSIGNED/al_00000286E4A272C0 ;  // al_ip/div_unsigned_gate.v(113)
  wire \u_DIV_UNSIGNED/al_00000286E4A27370 ;  // al_ip/div_unsigned_gate.v(102)
  wire \u_DIV_UNSIGNED/al_00000286E4A27420 ;  // al_ip/div_unsigned_gate.v(92)
  wire \u_DIV_UNSIGNED/al_00000286E4A276E0 ;  // al_ip/div_unsigned_gate.v(96)
  wire \u_DIV_UNSIGNED/al_00000286E4A27790 ;  // al_ip/div_unsigned_gate.v(101)
  wire \u_DIV_UNSIGNED/al_00000286E4A27B00 ;  // al_ip/div_unsigned_gate.v(111)
  wire \u_DIV_UNSIGNED/al_00000286E4A27BB0 ;  // al_ip/div_unsigned_gate.v(87)
  wire \u_DIV_UNSIGNED/al_00000286E4A27C60 ;  // al_ip/div_unsigned_gate.v(100)
  wire \u_DIV_UNSIGNED/al_00000286E4A27FD0 ;  // al_ip/div_unsigned_gate.v(117)
  wire \u_DIV_UNSIGNED/al_00000286E4A28080 ;  // al_ip/div_unsigned_gate.v(114)
  wire \u_DIV_UNSIGNED/al_00000286E4A28290 ;  // al_ip/div_unsigned_gate.v(119)
  wire \u_DIV_UNSIGNED/al_00000286E4A283F0 ;  // al_ip/div_unsigned_gate.v(97)
  wire \u_DIV_UNSIGNED/al_00000286E4A284A0 ;  // al_ip/div_unsigned_gate.v(106)
  wire \u_DIV_UNSIGNED/al_00000286E4A28810 ;  // al_ip/div_unsigned_gate.v(89)
  wire \u_DIV_UNSIGNED/al_00000286E4A28AD0 ;  // al_ip/div_unsigned_gate.v(95)
  wire \u_DIV_UNSIGNED/al_00000286E4A28B80 ;  // al_ip/div_unsigned_gate.v(107)
  wire \u_DIV_UNSIGNED/al_00000286E4A28C30 ;  // al_ip/div_unsigned_gate.v(99)
  wire \u_DIV_UNSIGNED/al_00000286E4A28CE0 ;  // al_ip/div_unsigned_gate.v(103)
  wire \u_DIV_UNSIGNED/al_00000286E4A28D90 ;  // al_ip/div_unsigned_gate.v(110)
  wire \u_DIV_UNSIGNED/al_00000286E4A28E40 ;  // al_ip/div_unsigned_gate.v(115)
  wire \u_DIV_UNSIGNED/al_00000286E5A5D8C0 ;  // al_ip/div_unsigned_gate.v(59)
  wire \u_DIV_UNSIGNED/al_00000286E5A5E1B0 ;  // al_ip/div_unsigned_gate.v(124)
  wire working;  // ../RTL/core/exu_mdu.v(46)

  assign o_mdu_rdidx[4] = o_will_rdidx[4];
  assign o_mdu_rdidx[3] = o_will_rdidx[3];
  assign o_mdu_rdidx[0] = o_will_rdidx[0];
  assign o_will_rdidx[2] = o_mdu_rdidx[2];
  assign o_will_rdidx[1] = o_mdu_rdidx[1];
  add_pu8_pu8_o8 add0 (
    .i0(cnt),
    .i1(8'b00000001),
    .o(n19));  // ../RTL/core/exu_mdu.v(115)
  eq_w8 eq0 (
    .i0(cnt),
    .i1(8'b00000001),
    .o(n18));  // ../RTL/core/exu_mdu.v(109)
  not i_flush_inv (i_flush_neg, i_flush);
  not mdu_finish_inv (mdu_finish_neg, mdu_finish);
  AL_DFF_X mul_finish_reg (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n30),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mul_finish));  // ../RTL/core/exu_mdu.v(96)
  not mul_start_inv (mul_start_neg, mul_start);
  AL_DFF_X mul_vld_reg (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n26),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(mul_vld));  // ../RTL/core/exu_mdu.v(96)
  mult_s32_s32_o64 mult0 (
    .i0(op1),
    .i1(op2),
    .o(mul_ss));  // ../RTL/core/exu_mdu.v(90)
  mult_u32_u32_o64 mult1 (
    .i0(op1),
    .i1(op2),
    .o({mul_uu[63:32],open_n0,open_n1,open_n2,open_n3,open_n4,open_n5,open_n6,open_n7,open_n8,open_n9,open_n10,open_n11,open_n12,open_n13,open_n14,open_n15,open_n16,open_n17,open_n18,open_n19,open_n20,open_n21,open_n22,open_n23,open_n24,open_n25,open_n26,open_n27,open_n28,open_n29,open_n30,open_n31}));  // ../RTL/core/exu_mdu.v(91)
  mult_s32_s33_o64 mult2 (
    .i0(op1),
    .i1({1'b0,op2}),
    .o({mul_su[63:32],open_n32,open_n33,open_n34,open_n35,open_n36,open_n37,open_n38,open_n39,open_n40,open_n41,open_n42,open_n43,open_n44,open_n45,open_n46,open_n47,open_n48,open_n49,open_n50,open_n51,open_n52,open_n53,open_n54,open_n55,open_n56,open_n57,open_n58,open_n59,open_n60,open_n61,open_n62,open_n63}));  // ../RTL/core/exu_mdu.v(92)
  and mux10_b0_sel_is_2 (mux10_b0_sel_is_2_o, i_rstn, mul_start);
  binary_mux_s1_w1 mux11_b0 (
    .i0(1'b0),
    .i1(i_mdu_op2[0]),
    .sel(mdu_vld),
    .o(n34[0]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b1 (
    .i0(1'b0),
    .i1(i_mdu_op2[1]),
    .sel(mdu_vld),
    .o(n34[1]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b10 (
    .i0(1'b0),
    .i1(i_mdu_op2[10]),
    .sel(mdu_vld),
    .o(n34[10]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b11 (
    .i0(1'b0),
    .i1(i_mdu_op2[11]),
    .sel(mdu_vld),
    .o(n34[11]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b12 (
    .i0(1'b0),
    .i1(i_mdu_op2[12]),
    .sel(mdu_vld),
    .o(n34[12]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b13 (
    .i0(1'b0),
    .i1(i_mdu_op2[13]),
    .sel(mdu_vld),
    .o(n34[13]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b14 (
    .i0(1'b0),
    .i1(i_mdu_op2[14]),
    .sel(mdu_vld),
    .o(n34[14]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b15 (
    .i0(1'b0),
    .i1(i_mdu_op2[15]),
    .sel(mdu_vld),
    .o(n34[15]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b16 (
    .i0(1'b0),
    .i1(i_mdu_op2[16]),
    .sel(mdu_vld),
    .o(n34[16]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b17 (
    .i0(1'b0),
    .i1(i_mdu_op2[17]),
    .sel(mdu_vld),
    .o(n34[17]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b18 (
    .i0(1'b0),
    .i1(i_mdu_op2[18]),
    .sel(mdu_vld),
    .o(n34[18]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b19 (
    .i0(1'b0),
    .i1(i_mdu_op2[19]),
    .sel(mdu_vld),
    .o(n34[19]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b2 (
    .i0(1'b0),
    .i1(i_mdu_op2[2]),
    .sel(mdu_vld),
    .o(n34[2]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b20 (
    .i0(1'b0),
    .i1(i_mdu_op2[20]),
    .sel(mdu_vld),
    .o(n34[20]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b21 (
    .i0(1'b0),
    .i1(i_mdu_op2[21]),
    .sel(mdu_vld),
    .o(n34[21]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b22 (
    .i0(1'b0),
    .i1(i_mdu_op2[22]),
    .sel(mdu_vld),
    .o(n34[22]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b23 (
    .i0(1'b0),
    .i1(i_mdu_op2[23]),
    .sel(mdu_vld),
    .o(n34[23]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b24 (
    .i0(1'b0),
    .i1(i_mdu_op2[24]),
    .sel(mdu_vld),
    .o(n34[24]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b25 (
    .i0(1'b0),
    .i1(i_mdu_op2[25]),
    .sel(mdu_vld),
    .o(n34[25]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b26 (
    .i0(1'b0),
    .i1(i_mdu_op2[26]),
    .sel(mdu_vld),
    .o(n34[26]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b27 (
    .i0(1'b0),
    .i1(i_mdu_op2[27]),
    .sel(mdu_vld),
    .o(n34[27]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b28 (
    .i0(1'b0),
    .i1(i_mdu_op2[28]),
    .sel(mdu_vld),
    .o(n34[28]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b29 (
    .i0(1'b0),
    .i1(i_mdu_op2[29]),
    .sel(mdu_vld),
    .o(n34[29]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b3 (
    .i0(1'b0),
    .i1(i_mdu_op2[3]),
    .sel(mdu_vld),
    .o(n34[3]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b30 (
    .i0(1'b0),
    .i1(i_mdu_op2[30]),
    .sel(mdu_vld),
    .o(n34[30]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b31 (
    .i0(1'b0),
    .i1(i_mdu_op2[31]),
    .sel(mdu_vld),
    .o(n34[31]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b4 (
    .i0(1'b0),
    .i1(i_mdu_op2[4]),
    .sel(mdu_vld),
    .o(n34[4]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b5 (
    .i0(1'b0),
    .i1(i_mdu_op2[5]),
    .sel(mdu_vld),
    .o(n34[5]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b6 (
    .i0(1'b0),
    .i1(i_mdu_op2[6]),
    .sel(mdu_vld),
    .o(n34[6]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b7 (
    .i0(1'b0),
    .i1(i_mdu_op2[7]),
    .sel(mdu_vld),
    .o(n34[7]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b8 (
    .i0(1'b0),
    .i1(i_mdu_op2[8]),
    .sel(mdu_vld),
    .o(n34[8]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux11_b9 (
    .i0(1'b0),
    .i1(i_mdu_op2[9]),
    .sel(mdu_vld),
    .o(n34[9]));  // ../RTL/core/exu_mdu.v(130)
  binary_mux_s1_w1 mux12_b0 (
    .i0(1'b0),
    .i1(i_mdu_op1[0]),
    .sel(mdu_vld),
    .o(n35[0]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b1 (
    .i0(1'b0),
    .i1(i_mdu_op1[1]),
    .sel(mdu_vld),
    .o(n35[1]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b10 (
    .i0(1'b0),
    .i1(i_mdu_op1[10]),
    .sel(mdu_vld),
    .o(n35[10]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b11 (
    .i0(1'b0),
    .i1(i_mdu_op1[11]),
    .sel(mdu_vld),
    .o(n35[11]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b12 (
    .i0(1'b0),
    .i1(i_mdu_op1[12]),
    .sel(mdu_vld),
    .o(n35[12]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b13 (
    .i0(1'b0),
    .i1(i_mdu_op1[13]),
    .sel(mdu_vld),
    .o(n35[13]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b14 (
    .i0(1'b0),
    .i1(i_mdu_op1[14]),
    .sel(mdu_vld),
    .o(n35[14]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b15 (
    .i0(1'b0),
    .i1(i_mdu_op1[15]),
    .sel(mdu_vld),
    .o(n35[15]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b16 (
    .i0(1'b0),
    .i1(i_mdu_op1[16]),
    .sel(mdu_vld),
    .o(n35[16]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b17 (
    .i0(1'b0),
    .i1(i_mdu_op1[17]),
    .sel(mdu_vld),
    .o(n35[17]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b18 (
    .i0(1'b0),
    .i1(i_mdu_op1[18]),
    .sel(mdu_vld),
    .o(n35[18]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b19 (
    .i0(1'b0),
    .i1(i_mdu_op1[19]),
    .sel(mdu_vld),
    .o(n35[19]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b2 (
    .i0(1'b0),
    .i1(i_mdu_op1[2]),
    .sel(mdu_vld),
    .o(n35[2]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b20 (
    .i0(1'b0),
    .i1(i_mdu_op1[20]),
    .sel(mdu_vld),
    .o(n35[20]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b21 (
    .i0(1'b0),
    .i1(i_mdu_op1[21]),
    .sel(mdu_vld),
    .o(n35[21]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b22 (
    .i0(1'b0),
    .i1(i_mdu_op1[22]),
    .sel(mdu_vld),
    .o(n35[22]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b23 (
    .i0(1'b0),
    .i1(i_mdu_op1[23]),
    .sel(mdu_vld),
    .o(n35[23]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b24 (
    .i0(1'b0),
    .i1(i_mdu_op1[24]),
    .sel(mdu_vld),
    .o(n35[24]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b25 (
    .i0(1'b0),
    .i1(i_mdu_op1[25]),
    .sel(mdu_vld),
    .o(n35[25]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b26 (
    .i0(1'b0),
    .i1(i_mdu_op1[26]),
    .sel(mdu_vld),
    .o(n35[26]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b27 (
    .i0(1'b0),
    .i1(i_mdu_op1[27]),
    .sel(mdu_vld),
    .o(n35[27]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b28 (
    .i0(1'b0),
    .i1(i_mdu_op1[28]),
    .sel(mdu_vld),
    .o(n35[28]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b29 (
    .i0(1'b0),
    .i1(i_mdu_op1[29]),
    .sel(mdu_vld),
    .o(n35[29]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b3 (
    .i0(1'b0),
    .i1(i_mdu_op1[3]),
    .sel(mdu_vld),
    .o(n35[3]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b30 (
    .i0(1'b0),
    .i1(i_mdu_op1[30]),
    .sel(mdu_vld),
    .o(n35[30]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b31 (
    .i0(1'b0),
    .i1(i_mdu_op1[31]),
    .sel(mdu_vld),
    .o(n35[31]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b4 (
    .i0(1'b0),
    .i1(i_mdu_op1[4]),
    .sel(mdu_vld),
    .o(n35[4]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b5 (
    .i0(1'b0),
    .i1(i_mdu_op1[5]),
    .sel(mdu_vld),
    .o(n35[5]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b6 (
    .i0(1'b0),
    .i1(i_mdu_op1[6]),
    .sel(mdu_vld),
    .o(n35[6]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b7 (
    .i0(1'b0),
    .i1(i_mdu_op1[7]),
    .sel(mdu_vld),
    .o(n35[7]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b8 (
    .i0(1'b0),
    .i1(i_mdu_op1[8]),
    .sel(mdu_vld),
    .o(n35[8]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux12_b9 (
    .i0(1'b0),
    .i1(i_mdu_op1[9]),
    .sel(mdu_vld),
    .o(n35[9]));  // ../RTL/core/exu_mdu.v(131)
  binary_mux_s1_w1 mux13_b0 (
    .i0(div_signed_rem[0]),
    .i1(n37[0]),
    .sel(rem_op1_sym),
    .o(n38[0]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b1 (
    .i0(div_signed_rem[1]),
    .i1(n37[1]),
    .sel(rem_op1_sym),
    .o(n38[1]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b10 (
    .i0(div_signed_rem[10]),
    .i1(n37[10]),
    .sel(rem_op1_sym),
    .o(n38[10]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b11 (
    .i0(div_signed_rem[11]),
    .i1(n37[11]),
    .sel(rem_op1_sym),
    .o(n38[11]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b12 (
    .i0(div_signed_rem[12]),
    .i1(n37[12]),
    .sel(rem_op1_sym),
    .o(n38[12]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b13 (
    .i0(div_signed_rem[13]),
    .i1(n37[13]),
    .sel(rem_op1_sym),
    .o(n38[13]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b14 (
    .i0(div_signed_rem[14]),
    .i1(n37[14]),
    .sel(rem_op1_sym),
    .o(n38[14]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b15 (
    .i0(div_signed_rem[15]),
    .i1(n37[15]),
    .sel(rem_op1_sym),
    .o(n38[15]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b16 (
    .i0(div_signed_rem[16]),
    .i1(n37[16]),
    .sel(rem_op1_sym),
    .o(n38[16]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b17 (
    .i0(div_signed_rem[17]),
    .i1(n37[17]),
    .sel(rem_op1_sym),
    .o(n38[17]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b18 (
    .i0(div_signed_rem[18]),
    .i1(n37[18]),
    .sel(rem_op1_sym),
    .o(n38[18]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b19 (
    .i0(div_signed_rem[19]),
    .i1(n37[19]),
    .sel(rem_op1_sym),
    .o(n38[19]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b2 (
    .i0(div_signed_rem[2]),
    .i1(n37[2]),
    .sel(rem_op1_sym),
    .o(n38[2]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b20 (
    .i0(div_signed_rem[20]),
    .i1(n37[20]),
    .sel(rem_op1_sym),
    .o(n38[20]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b21 (
    .i0(div_signed_rem[21]),
    .i1(n37[21]),
    .sel(rem_op1_sym),
    .o(n38[21]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b22 (
    .i0(div_signed_rem[22]),
    .i1(n37[22]),
    .sel(rem_op1_sym),
    .o(n38[22]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b23 (
    .i0(div_signed_rem[23]),
    .i1(n37[23]),
    .sel(rem_op1_sym),
    .o(n38[23]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b24 (
    .i0(div_signed_rem[24]),
    .i1(n37[24]),
    .sel(rem_op1_sym),
    .o(n38[24]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b25 (
    .i0(div_signed_rem[25]),
    .i1(n37[25]),
    .sel(rem_op1_sym),
    .o(n38[25]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b26 (
    .i0(div_signed_rem[26]),
    .i1(n37[26]),
    .sel(rem_op1_sym),
    .o(n38[26]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b27 (
    .i0(div_signed_rem[27]),
    .i1(n37[27]),
    .sel(rem_op1_sym),
    .o(n38[27]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b28 (
    .i0(div_signed_rem[28]),
    .i1(n37[28]),
    .sel(rem_op1_sym),
    .o(n38[28]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b29 (
    .i0(div_signed_rem[29]),
    .i1(n37[29]),
    .sel(rem_op1_sym),
    .o(n38[29]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b3 (
    .i0(div_signed_rem[3]),
    .i1(n37[3]),
    .sel(rem_op1_sym),
    .o(n38[3]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b30 (
    .i0(div_signed_rem[30]),
    .i1(n37[30]),
    .sel(rem_op1_sym),
    .o(n38[30]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b31 (
    .i0(div_signed_rem[31]),
    .i1(n37[31]),
    .sel(rem_op1_sym),
    .o(n38[31]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b4 (
    .i0(div_signed_rem[4]),
    .i1(n37[4]),
    .sel(rem_op1_sym),
    .o(n38[4]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b5 (
    .i0(div_signed_rem[5]),
    .i1(n37[5]),
    .sel(rem_op1_sym),
    .o(n38[5]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b6 (
    .i0(div_signed_rem[6]),
    .i1(n37[6]),
    .sel(rem_op1_sym),
    .o(n38[6]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b7 (
    .i0(div_signed_rem[7]),
    .i1(n37[7]),
    .sel(rem_op1_sym),
    .o(n38[7]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b8 (
    .i0(div_signed_rem[8]),
    .i1(n37[8]),
    .sel(rem_op1_sym),
    .o(n38[8]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux13_b9 (
    .i0(div_signed_rem[9]),
    .i1(n37[9]),
    .sel(rem_op1_sym),
    .o(n38[9]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux14_b0 (
    .i0(1'b0),
    .i1(div_unsigned_rem[0]),
    .sel(mduinfo[8]),
    .o(n39[0]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b1 (
    .i0(1'b0),
    .i1(div_unsigned_rem[1]),
    .sel(mduinfo[8]),
    .o(n39[1]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b10 (
    .i0(1'b0),
    .i1(div_unsigned_rem[10]),
    .sel(mduinfo[8]),
    .o(n39[10]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b11 (
    .i0(1'b0),
    .i1(div_unsigned_rem[11]),
    .sel(mduinfo[8]),
    .o(n39[11]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b12 (
    .i0(1'b0),
    .i1(div_unsigned_rem[12]),
    .sel(mduinfo[8]),
    .o(n39[12]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b13 (
    .i0(1'b0),
    .i1(div_unsigned_rem[13]),
    .sel(mduinfo[8]),
    .o(n39[13]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b14 (
    .i0(1'b0),
    .i1(div_unsigned_rem[14]),
    .sel(mduinfo[8]),
    .o(n39[14]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b15 (
    .i0(1'b0),
    .i1(div_unsigned_rem[15]),
    .sel(mduinfo[8]),
    .o(n39[15]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b16 (
    .i0(1'b0),
    .i1(div_unsigned_rem[16]),
    .sel(mduinfo[8]),
    .o(n39[16]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b17 (
    .i0(1'b0),
    .i1(div_unsigned_rem[17]),
    .sel(mduinfo[8]),
    .o(n39[17]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b18 (
    .i0(1'b0),
    .i1(div_unsigned_rem[18]),
    .sel(mduinfo[8]),
    .o(n39[18]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b19 (
    .i0(1'b0),
    .i1(div_unsigned_rem[19]),
    .sel(mduinfo[8]),
    .o(n39[19]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b2 (
    .i0(1'b0),
    .i1(div_unsigned_rem[2]),
    .sel(mduinfo[8]),
    .o(n39[2]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b20 (
    .i0(1'b0),
    .i1(div_unsigned_rem[20]),
    .sel(mduinfo[8]),
    .o(n39[20]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b21 (
    .i0(1'b0),
    .i1(div_unsigned_rem[21]),
    .sel(mduinfo[8]),
    .o(n39[21]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b22 (
    .i0(1'b0),
    .i1(div_unsigned_rem[22]),
    .sel(mduinfo[8]),
    .o(n39[22]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b23 (
    .i0(1'b0),
    .i1(div_unsigned_rem[23]),
    .sel(mduinfo[8]),
    .o(n39[23]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b24 (
    .i0(1'b0),
    .i1(div_unsigned_rem[24]),
    .sel(mduinfo[8]),
    .o(n39[24]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b25 (
    .i0(1'b0),
    .i1(div_unsigned_rem[25]),
    .sel(mduinfo[8]),
    .o(n39[25]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b26 (
    .i0(1'b0),
    .i1(div_unsigned_rem[26]),
    .sel(mduinfo[8]),
    .o(n39[26]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b27 (
    .i0(1'b0),
    .i1(div_unsigned_rem[27]),
    .sel(mduinfo[8]),
    .o(n39[27]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b28 (
    .i0(1'b0),
    .i1(div_unsigned_rem[28]),
    .sel(mduinfo[8]),
    .o(n39[28]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b29 (
    .i0(1'b0),
    .i1(div_unsigned_rem[29]),
    .sel(mduinfo[8]),
    .o(n39[29]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b3 (
    .i0(1'b0),
    .i1(div_unsigned_rem[3]),
    .sel(mduinfo[8]),
    .o(n39[3]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b30 (
    .i0(1'b0),
    .i1(div_unsigned_rem[30]),
    .sel(mduinfo[8]),
    .o(n39[30]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b31 (
    .i0(1'b0),
    .i1(div_unsigned_rem[31]),
    .sel(mduinfo[8]),
    .o(n39[31]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b4 (
    .i0(1'b0),
    .i1(div_unsigned_rem[4]),
    .sel(mduinfo[8]),
    .o(n39[4]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b5 (
    .i0(1'b0),
    .i1(div_unsigned_rem[5]),
    .sel(mduinfo[8]),
    .o(n39[5]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b6 (
    .i0(1'b0),
    .i1(div_unsigned_rem[6]),
    .sel(mduinfo[8]),
    .o(n39[6]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b7 (
    .i0(1'b0),
    .i1(div_unsigned_rem[7]),
    .sel(mduinfo[8]),
    .o(n39[7]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b8 (
    .i0(1'b0),
    .i1(div_unsigned_rem[8]),
    .sel(mduinfo[8]),
    .o(n39[8]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux14_b9 (
    .i0(1'b0),
    .i1(div_unsigned_rem[9]),
    .sel(mduinfo[8]),
    .o(n39[9]));  // ../RTL/core/exu_mdu.v(166)
  binary_mux_s1_w1 mux15_b0 (
    .i0(n39[0]),
    .i1(n38[0]),
    .sel(mduinfo[7]),
    .o(n40[0]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b1 (
    .i0(n39[1]),
    .i1(n38[1]),
    .sel(mduinfo[7]),
    .o(n40[1]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b10 (
    .i0(n39[10]),
    .i1(n38[10]),
    .sel(mduinfo[7]),
    .o(n40[10]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b11 (
    .i0(n39[11]),
    .i1(n38[11]),
    .sel(mduinfo[7]),
    .o(n40[11]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b12 (
    .i0(n39[12]),
    .i1(n38[12]),
    .sel(mduinfo[7]),
    .o(n40[12]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b13 (
    .i0(n39[13]),
    .i1(n38[13]),
    .sel(mduinfo[7]),
    .o(n40[13]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b14 (
    .i0(n39[14]),
    .i1(n38[14]),
    .sel(mduinfo[7]),
    .o(n40[14]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b15 (
    .i0(n39[15]),
    .i1(n38[15]),
    .sel(mduinfo[7]),
    .o(n40[15]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b16 (
    .i0(n39[16]),
    .i1(n38[16]),
    .sel(mduinfo[7]),
    .o(n40[16]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b17 (
    .i0(n39[17]),
    .i1(n38[17]),
    .sel(mduinfo[7]),
    .o(n40[17]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b18 (
    .i0(n39[18]),
    .i1(n38[18]),
    .sel(mduinfo[7]),
    .o(n40[18]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b19 (
    .i0(n39[19]),
    .i1(n38[19]),
    .sel(mduinfo[7]),
    .o(n40[19]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b2 (
    .i0(n39[2]),
    .i1(n38[2]),
    .sel(mduinfo[7]),
    .o(n40[2]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b20 (
    .i0(n39[20]),
    .i1(n38[20]),
    .sel(mduinfo[7]),
    .o(n40[20]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b21 (
    .i0(n39[21]),
    .i1(n38[21]),
    .sel(mduinfo[7]),
    .o(n40[21]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b22 (
    .i0(n39[22]),
    .i1(n38[22]),
    .sel(mduinfo[7]),
    .o(n40[22]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b23 (
    .i0(n39[23]),
    .i1(n38[23]),
    .sel(mduinfo[7]),
    .o(n40[23]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b24 (
    .i0(n39[24]),
    .i1(n38[24]),
    .sel(mduinfo[7]),
    .o(n40[24]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b25 (
    .i0(n39[25]),
    .i1(n38[25]),
    .sel(mduinfo[7]),
    .o(n40[25]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b26 (
    .i0(n39[26]),
    .i1(n38[26]),
    .sel(mduinfo[7]),
    .o(n40[26]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b27 (
    .i0(n39[27]),
    .i1(n38[27]),
    .sel(mduinfo[7]),
    .o(n40[27]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b28 (
    .i0(n39[28]),
    .i1(n38[28]),
    .sel(mduinfo[7]),
    .o(n40[28]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b29 (
    .i0(n39[29]),
    .i1(n38[29]),
    .sel(mduinfo[7]),
    .o(n40[29]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b3 (
    .i0(n39[3]),
    .i1(n38[3]),
    .sel(mduinfo[7]),
    .o(n40[3]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b30 (
    .i0(n39[30]),
    .i1(n38[30]),
    .sel(mduinfo[7]),
    .o(n40[30]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b31 (
    .i0(n39[31]),
    .i1(n38[31]),
    .sel(mduinfo[7]),
    .o(n40[31]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b4 (
    .i0(n39[4]),
    .i1(n38[4]),
    .sel(mduinfo[7]),
    .o(n40[4]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b5 (
    .i0(n39[5]),
    .i1(n38[5]),
    .sel(mduinfo[7]),
    .o(n40[5]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b6 (
    .i0(n39[6]),
    .i1(n38[6]),
    .sel(mduinfo[7]),
    .o(n40[6]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b7 (
    .i0(n39[7]),
    .i1(n38[7]),
    .sel(mduinfo[7]),
    .o(n40[7]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b8 (
    .i0(n39[8]),
    .i1(n38[8]),
    .sel(mduinfo[7]),
    .o(n40[8]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux15_b9 (
    .i0(n39[9]),
    .i1(n38[9]),
    .sel(mduinfo[7]),
    .o(n40[9]));  // ../RTL/core/exu_mdu.v(165)
  binary_mux_s1_w1 mux16_b0 (
    .i0(n40[0]),
    .i1(div_unsigned_quo[0]),
    .sel(mduinfo[6]),
    .o(n41[0]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b1 (
    .i0(n40[1]),
    .i1(div_unsigned_quo[1]),
    .sel(mduinfo[6]),
    .o(n41[1]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b10 (
    .i0(n40[10]),
    .i1(div_unsigned_quo[10]),
    .sel(mduinfo[6]),
    .o(n41[10]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b11 (
    .i0(n40[11]),
    .i1(div_unsigned_quo[11]),
    .sel(mduinfo[6]),
    .o(n41[11]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b12 (
    .i0(n40[12]),
    .i1(div_unsigned_quo[12]),
    .sel(mduinfo[6]),
    .o(n41[12]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b13 (
    .i0(n40[13]),
    .i1(div_unsigned_quo[13]),
    .sel(mduinfo[6]),
    .o(n41[13]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b14 (
    .i0(n40[14]),
    .i1(div_unsigned_quo[14]),
    .sel(mduinfo[6]),
    .o(n41[14]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b15 (
    .i0(n40[15]),
    .i1(div_unsigned_quo[15]),
    .sel(mduinfo[6]),
    .o(n41[15]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b16 (
    .i0(n40[16]),
    .i1(div_unsigned_quo[16]),
    .sel(mduinfo[6]),
    .o(n41[16]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b17 (
    .i0(n40[17]),
    .i1(div_unsigned_quo[17]),
    .sel(mduinfo[6]),
    .o(n41[17]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b18 (
    .i0(n40[18]),
    .i1(div_unsigned_quo[18]),
    .sel(mduinfo[6]),
    .o(n41[18]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b19 (
    .i0(n40[19]),
    .i1(div_unsigned_quo[19]),
    .sel(mduinfo[6]),
    .o(n41[19]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b2 (
    .i0(n40[2]),
    .i1(div_unsigned_quo[2]),
    .sel(mduinfo[6]),
    .o(n41[2]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b20 (
    .i0(n40[20]),
    .i1(div_unsigned_quo[20]),
    .sel(mduinfo[6]),
    .o(n41[20]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b21 (
    .i0(n40[21]),
    .i1(div_unsigned_quo[21]),
    .sel(mduinfo[6]),
    .o(n41[21]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b22 (
    .i0(n40[22]),
    .i1(div_unsigned_quo[22]),
    .sel(mduinfo[6]),
    .o(n41[22]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b23 (
    .i0(n40[23]),
    .i1(div_unsigned_quo[23]),
    .sel(mduinfo[6]),
    .o(n41[23]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b24 (
    .i0(n40[24]),
    .i1(div_unsigned_quo[24]),
    .sel(mduinfo[6]),
    .o(n41[24]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b25 (
    .i0(n40[25]),
    .i1(div_unsigned_quo[25]),
    .sel(mduinfo[6]),
    .o(n41[25]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b26 (
    .i0(n40[26]),
    .i1(div_unsigned_quo[26]),
    .sel(mduinfo[6]),
    .o(n41[26]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b27 (
    .i0(n40[27]),
    .i1(div_unsigned_quo[27]),
    .sel(mduinfo[6]),
    .o(n41[27]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b28 (
    .i0(n40[28]),
    .i1(div_unsigned_quo[28]),
    .sel(mduinfo[6]),
    .o(n41[28]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b29 (
    .i0(n40[29]),
    .i1(div_unsigned_quo[29]),
    .sel(mduinfo[6]),
    .o(n41[29]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b3 (
    .i0(n40[3]),
    .i1(div_unsigned_quo[3]),
    .sel(mduinfo[6]),
    .o(n41[3]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b30 (
    .i0(n40[30]),
    .i1(div_unsigned_quo[30]),
    .sel(mduinfo[6]),
    .o(n41[30]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b31 (
    .i0(n40[31]),
    .i1(div_unsigned_quo[31]),
    .sel(mduinfo[6]),
    .o(n41[31]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b4 (
    .i0(n40[4]),
    .i1(div_unsigned_quo[4]),
    .sel(mduinfo[6]),
    .o(n41[4]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b5 (
    .i0(n40[5]),
    .i1(div_unsigned_quo[5]),
    .sel(mduinfo[6]),
    .o(n41[5]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b6 (
    .i0(n40[6]),
    .i1(div_unsigned_quo[6]),
    .sel(mduinfo[6]),
    .o(n41[6]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b7 (
    .i0(n40[7]),
    .i1(div_unsigned_quo[7]),
    .sel(mduinfo[6]),
    .o(n41[7]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b8 (
    .i0(n40[8]),
    .i1(div_unsigned_quo[8]),
    .sel(mduinfo[6]),
    .o(n41[8]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux16_b9 (
    .i0(n40[9]),
    .i1(div_unsigned_quo[9]),
    .sel(mduinfo[6]),
    .o(n41[9]));  // ../RTL/core/exu_mdu.v(164)
  binary_mux_s1_w1 mux17_b0 (
    .i0(n41[0]),
    .i1(div_signed_quo[0]),
    .sel(mduinfo[5]),
    .o(n42[0]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b1 (
    .i0(n41[1]),
    .i1(div_signed_quo[1]),
    .sel(mduinfo[5]),
    .o(n42[1]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b10 (
    .i0(n41[10]),
    .i1(div_signed_quo[10]),
    .sel(mduinfo[5]),
    .o(n42[10]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b11 (
    .i0(n41[11]),
    .i1(div_signed_quo[11]),
    .sel(mduinfo[5]),
    .o(n42[11]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b12 (
    .i0(n41[12]),
    .i1(div_signed_quo[12]),
    .sel(mduinfo[5]),
    .o(n42[12]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b13 (
    .i0(n41[13]),
    .i1(div_signed_quo[13]),
    .sel(mduinfo[5]),
    .o(n42[13]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b14 (
    .i0(n41[14]),
    .i1(div_signed_quo[14]),
    .sel(mduinfo[5]),
    .o(n42[14]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b15 (
    .i0(n41[15]),
    .i1(div_signed_quo[15]),
    .sel(mduinfo[5]),
    .o(n42[15]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b16 (
    .i0(n41[16]),
    .i1(div_signed_quo[16]),
    .sel(mduinfo[5]),
    .o(n42[16]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b17 (
    .i0(n41[17]),
    .i1(div_signed_quo[17]),
    .sel(mduinfo[5]),
    .o(n42[17]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b18 (
    .i0(n41[18]),
    .i1(div_signed_quo[18]),
    .sel(mduinfo[5]),
    .o(n42[18]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b19 (
    .i0(n41[19]),
    .i1(div_signed_quo[19]),
    .sel(mduinfo[5]),
    .o(n42[19]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b2 (
    .i0(n41[2]),
    .i1(div_signed_quo[2]),
    .sel(mduinfo[5]),
    .o(n42[2]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b20 (
    .i0(n41[20]),
    .i1(div_signed_quo[20]),
    .sel(mduinfo[5]),
    .o(n42[20]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b21 (
    .i0(n41[21]),
    .i1(div_signed_quo[21]),
    .sel(mduinfo[5]),
    .o(n42[21]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b22 (
    .i0(n41[22]),
    .i1(div_signed_quo[22]),
    .sel(mduinfo[5]),
    .o(n42[22]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b23 (
    .i0(n41[23]),
    .i1(div_signed_quo[23]),
    .sel(mduinfo[5]),
    .o(n42[23]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b24 (
    .i0(n41[24]),
    .i1(div_signed_quo[24]),
    .sel(mduinfo[5]),
    .o(n42[24]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b25 (
    .i0(n41[25]),
    .i1(div_signed_quo[25]),
    .sel(mduinfo[5]),
    .o(n42[25]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b26 (
    .i0(n41[26]),
    .i1(div_signed_quo[26]),
    .sel(mduinfo[5]),
    .o(n42[26]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b27 (
    .i0(n41[27]),
    .i1(div_signed_quo[27]),
    .sel(mduinfo[5]),
    .o(n42[27]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b28 (
    .i0(n41[28]),
    .i1(div_signed_quo[28]),
    .sel(mduinfo[5]),
    .o(n42[28]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b29 (
    .i0(n41[29]),
    .i1(div_signed_quo[29]),
    .sel(mduinfo[5]),
    .o(n42[29]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b3 (
    .i0(n41[3]),
    .i1(div_signed_quo[3]),
    .sel(mduinfo[5]),
    .o(n42[3]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b30 (
    .i0(n41[30]),
    .i1(div_signed_quo[30]),
    .sel(mduinfo[5]),
    .o(n42[30]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b31 (
    .i0(n41[31]),
    .i1(div_signed_quo[31]),
    .sel(mduinfo[5]),
    .o(n42[31]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b4 (
    .i0(n41[4]),
    .i1(div_signed_quo[4]),
    .sel(mduinfo[5]),
    .o(n42[4]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b5 (
    .i0(n41[5]),
    .i1(div_signed_quo[5]),
    .sel(mduinfo[5]),
    .o(n42[5]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b6 (
    .i0(n41[6]),
    .i1(div_signed_quo[6]),
    .sel(mduinfo[5]),
    .o(n42[6]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b7 (
    .i0(n41[7]),
    .i1(div_signed_quo[7]),
    .sel(mduinfo[5]),
    .o(n42[7]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b8 (
    .i0(n41[8]),
    .i1(div_signed_quo[8]),
    .sel(mduinfo[5]),
    .o(n42[8]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux17_b9 (
    .i0(n41[9]),
    .i1(div_signed_quo[9]),
    .sel(mduinfo[5]),
    .o(n42[9]));  // ../RTL/core/exu_mdu.v(163)
  binary_mux_s1_w1 mux18_b0 (
    .i0(n42[0]),
    .i1(mul_su[32]),
    .sel(mduinfo[3]),
    .o(n43[0]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b1 (
    .i0(n42[1]),
    .i1(mul_su[33]),
    .sel(mduinfo[3]),
    .o(n43[1]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b10 (
    .i0(n42[10]),
    .i1(mul_su[42]),
    .sel(mduinfo[3]),
    .o(n43[10]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b11 (
    .i0(n42[11]),
    .i1(mul_su[43]),
    .sel(mduinfo[3]),
    .o(n43[11]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b12 (
    .i0(n42[12]),
    .i1(mul_su[44]),
    .sel(mduinfo[3]),
    .o(n43[12]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b13 (
    .i0(n42[13]),
    .i1(mul_su[45]),
    .sel(mduinfo[3]),
    .o(n43[13]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b14 (
    .i0(n42[14]),
    .i1(mul_su[46]),
    .sel(mduinfo[3]),
    .o(n43[14]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b15 (
    .i0(n42[15]),
    .i1(mul_su[47]),
    .sel(mduinfo[3]),
    .o(n43[15]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b16 (
    .i0(n42[16]),
    .i1(mul_su[48]),
    .sel(mduinfo[3]),
    .o(n43[16]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b17 (
    .i0(n42[17]),
    .i1(mul_su[49]),
    .sel(mduinfo[3]),
    .o(n43[17]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b18 (
    .i0(n42[18]),
    .i1(mul_su[50]),
    .sel(mduinfo[3]),
    .o(n43[18]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b19 (
    .i0(n42[19]),
    .i1(mul_su[51]),
    .sel(mduinfo[3]),
    .o(n43[19]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b2 (
    .i0(n42[2]),
    .i1(mul_su[34]),
    .sel(mduinfo[3]),
    .o(n43[2]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b20 (
    .i0(n42[20]),
    .i1(mul_su[52]),
    .sel(mduinfo[3]),
    .o(n43[20]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b21 (
    .i0(n42[21]),
    .i1(mul_su[53]),
    .sel(mduinfo[3]),
    .o(n43[21]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b22 (
    .i0(n42[22]),
    .i1(mul_su[54]),
    .sel(mduinfo[3]),
    .o(n43[22]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b23 (
    .i0(n42[23]),
    .i1(mul_su[55]),
    .sel(mduinfo[3]),
    .o(n43[23]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b24 (
    .i0(n42[24]),
    .i1(mul_su[56]),
    .sel(mduinfo[3]),
    .o(n43[24]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b25 (
    .i0(n42[25]),
    .i1(mul_su[57]),
    .sel(mduinfo[3]),
    .o(n43[25]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b26 (
    .i0(n42[26]),
    .i1(mul_su[58]),
    .sel(mduinfo[3]),
    .o(n43[26]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b27 (
    .i0(n42[27]),
    .i1(mul_su[59]),
    .sel(mduinfo[3]),
    .o(n43[27]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b28 (
    .i0(n42[28]),
    .i1(mul_su[60]),
    .sel(mduinfo[3]),
    .o(n43[28]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b29 (
    .i0(n42[29]),
    .i1(mul_su[61]),
    .sel(mduinfo[3]),
    .o(n43[29]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b3 (
    .i0(n42[3]),
    .i1(mul_su[35]),
    .sel(mduinfo[3]),
    .o(n43[3]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b30 (
    .i0(n42[30]),
    .i1(mul_su[62]),
    .sel(mduinfo[3]),
    .o(n43[30]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b31 (
    .i0(n42[31]),
    .i1(mul_su[63]),
    .sel(mduinfo[3]),
    .o(n43[31]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b4 (
    .i0(n42[4]),
    .i1(mul_su[36]),
    .sel(mduinfo[3]),
    .o(n43[4]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b5 (
    .i0(n42[5]),
    .i1(mul_su[37]),
    .sel(mduinfo[3]),
    .o(n43[5]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b6 (
    .i0(n42[6]),
    .i1(mul_su[38]),
    .sel(mduinfo[3]),
    .o(n43[6]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b7 (
    .i0(n42[7]),
    .i1(mul_su[39]),
    .sel(mduinfo[3]),
    .o(n43[7]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b8 (
    .i0(n42[8]),
    .i1(mul_su[40]),
    .sel(mduinfo[3]),
    .o(n43[8]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux18_b9 (
    .i0(n42[9]),
    .i1(mul_su[41]),
    .sel(mduinfo[3]),
    .o(n43[9]));  // ../RTL/core/exu_mdu.v(162)
  binary_mux_s1_w1 mux19_b0 (
    .i0(n43[0]),
    .i1(mul_uu[32]),
    .sel(mduinfo[4]),
    .o(n44[0]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b1 (
    .i0(n43[1]),
    .i1(mul_uu[33]),
    .sel(mduinfo[4]),
    .o(n44[1]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b10 (
    .i0(n43[10]),
    .i1(mul_uu[42]),
    .sel(mduinfo[4]),
    .o(n44[10]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b11 (
    .i0(n43[11]),
    .i1(mul_uu[43]),
    .sel(mduinfo[4]),
    .o(n44[11]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b12 (
    .i0(n43[12]),
    .i1(mul_uu[44]),
    .sel(mduinfo[4]),
    .o(n44[12]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b13 (
    .i0(n43[13]),
    .i1(mul_uu[45]),
    .sel(mduinfo[4]),
    .o(n44[13]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b14 (
    .i0(n43[14]),
    .i1(mul_uu[46]),
    .sel(mduinfo[4]),
    .o(n44[14]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b15 (
    .i0(n43[15]),
    .i1(mul_uu[47]),
    .sel(mduinfo[4]),
    .o(n44[15]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b16 (
    .i0(n43[16]),
    .i1(mul_uu[48]),
    .sel(mduinfo[4]),
    .o(n44[16]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b17 (
    .i0(n43[17]),
    .i1(mul_uu[49]),
    .sel(mduinfo[4]),
    .o(n44[17]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b18 (
    .i0(n43[18]),
    .i1(mul_uu[50]),
    .sel(mduinfo[4]),
    .o(n44[18]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b19 (
    .i0(n43[19]),
    .i1(mul_uu[51]),
    .sel(mduinfo[4]),
    .o(n44[19]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b2 (
    .i0(n43[2]),
    .i1(mul_uu[34]),
    .sel(mduinfo[4]),
    .o(n44[2]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b20 (
    .i0(n43[20]),
    .i1(mul_uu[52]),
    .sel(mduinfo[4]),
    .o(n44[20]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b21 (
    .i0(n43[21]),
    .i1(mul_uu[53]),
    .sel(mduinfo[4]),
    .o(n44[21]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b22 (
    .i0(n43[22]),
    .i1(mul_uu[54]),
    .sel(mduinfo[4]),
    .o(n44[22]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b23 (
    .i0(n43[23]),
    .i1(mul_uu[55]),
    .sel(mduinfo[4]),
    .o(n44[23]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b24 (
    .i0(n43[24]),
    .i1(mul_uu[56]),
    .sel(mduinfo[4]),
    .o(n44[24]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b25 (
    .i0(n43[25]),
    .i1(mul_uu[57]),
    .sel(mduinfo[4]),
    .o(n44[25]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b26 (
    .i0(n43[26]),
    .i1(mul_uu[58]),
    .sel(mduinfo[4]),
    .o(n44[26]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b27 (
    .i0(n43[27]),
    .i1(mul_uu[59]),
    .sel(mduinfo[4]),
    .o(n44[27]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b28 (
    .i0(n43[28]),
    .i1(mul_uu[60]),
    .sel(mduinfo[4]),
    .o(n44[28]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b29 (
    .i0(n43[29]),
    .i1(mul_uu[61]),
    .sel(mduinfo[4]),
    .o(n44[29]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b3 (
    .i0(n43[3]),
    .i1(mul_uu[35]),
    .sel(mduinfo[4]),
    .o(n44[3]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b30 (
    .i0(n43[30]),
    .i1(mul_uu[62]),
    .sel(mduinfo[4]),
    .o(n44[30]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b31 (
    .i0(n43[31]),
    .i1(mul_uu[63]),
    .sel(mduinfo[4]),
    .o(n44[31]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b4 (
    .i0(n43[4]),
    .i1(mul_uu[36]),
    .sel(mduinfo[4]),
    .o(n44[4]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b5 (
    .i0(n43[5]),
    .i1(mul_uu[37]),
    .sel(mduinfo[4]),
    .o(n44[5]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b6 (
    .i0(n43[6]),
    .i1(mul_uu[38]),
    .sel(mduinfo[4]),
    .o(n44[6]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b7 (
    .i0(n43[7]),
    .i1(mul_uu[39]),
    .sel(mduinfo[4]),
    .o(n44[7]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b8 (
    .i0(n43[8]),
    .i1(mul_uu[40]),
    .sel(mduinfo[4]),
    .o(n44[8]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux19_b9 (
    .i0(n43[9]),
    .i1(mul_uu[41]),
    .sel(mduinfo[4]),
    .o(n44[9]));  // ../RTL/core/exu_mdu.v(161)
  binary_mux_s1_w1 mux20_b0 (
    .i0(n44[0]),
    .i1(mul_ss[32]),
    .sel(mduinfo[2]),
    .o(n45[0]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b1 (
    .i0(n44[1]),
    .i1(mul_ss[33]),
    .sel(mduinfo[2]),
    .o(n45[1]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b10 (
    .i0(n44[10]),
    .i1(mul_ss[42]),
    .sel(mduinfo[2]),
    .o(n45[10]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b11 (
    .i0(n44[11]),
    .i1(mul_ss[43]),
    .sel(mduinfo[2]),
    .o(n45[11]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b12 (
    .i0(n44[12]),
    .i1(mul_ss[44]),
    .sel(mduinfo[2]),
    .o(n45[12]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b13 (
    .i0(n44[13]),
    .i1(mul_ss[45]),
    .sel(mduinfo[2]),
    .o(n45[13]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b14 (
    .i0(n44[14]),
    .i1(mul_ss[46]),
    .sel(mduinfo[2]),
    .o(n45[14]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b15 (
    .i0(n44[15]),
    .i1(mul_ss[47]),
    .sel(mduinfo[2]),
    .o(n45[15]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b16 (
    .i0(n44[16]),
    .i1(mul_ss[48]),
    .sel(mduinfo[2]),
    .o(n45[16]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b17 (
    .i0(n44[17]),
    .i1(mul_ss[49]),
    .sel(mduinfo[2]),
    .o(n45[17]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b18 (
    .i0(n44[18]),
    .i1(mul_ss[50]),
    .sel(mduinfo[2]),
    .o(n45[18]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b19 (
    .i0(n44[19]),
    .i1(mul_ss[51]),
    .sel(mduinfo[2]),
    .o(n45[19]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b2 (
    .i0(n44[2]),
    .i1(mul_ss[34]),
    .sel(mduinfo[2]),
    .o(n45[2]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b20 (
    .i0(n44[20]),
    .i1(mul_ss[52]),
    .sel(mduinfo[2]),
    .o(n45[20]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b21 (
    .i0(n44[21]),
    .i1(mul_ss[53]),
    .sel(mduinfo[2]),
    .o(n45[21]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b22 (
    .i0(n44[22]),
    .i1(mul_ss[54]),
    .sel(mduinfo[2]),
    .o(n45[22]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b23 (
    .i0(n44[23]),
    .i1(mul_ss[55]),
    .sel(mduinfo[2]),
    .o(n45[23]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b24 (
    .i0(n44[24]),
    .i1(mul_ss[56]),
    .sel(mduinfo[2]),
    .o(n45[24]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b25 (
    .i0(n44[25]),
    .i1(mul_ss[57]),
    .sel(mduinfo[2]),
    .o(n45[25]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b26 (
    .i0(n44[26]),
    .i1(mul_ss[58]),
    .sel(mduinfo[2]),
    .o(n45[26]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b27 (
    .i0(n44[27]),
    .i1(mul_ss[59]),
    .sel(mduinfo[2]),
    .o(n45[27]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b28 (
    .i0(n44[28]),
    .i1(mul_ss[60]),
    .sel(mduinfo[2]),
    .o(n45[28]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b29 (
    .i0(n44[29]),
    .i1(mul_ss[61]),
    .sel(mduinfo[2]),
    .o(n45[29]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b3 (
    .i0(n44[3]),
    .i1(mul_ss[35]),
    .sel(mduinfo[2]),
    .o(n45[3]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b30 (
    .i0(n44[30]),
    .i1(mul_ss[62]),
    .sel(mduinfo[2]),
    .o(n45[30]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b31 (
    .i0(n44[31]),
    .i1(mul_ss[63]),
    .sel(mduinfo[2]),
    .o(n45[31]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b4 (
    .i0(n44[4]),
    .i1(mul_ss[36]),
    .sel(mduinfo[2]),
    .o(n45[4]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b5 (
    .i0(n44[5]),
    .i1(mul_ss[37]),
    .sel(mduinfo[2]),
    .o(n45[5]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b6 (
    .i0(n44[6]),
    .i1(mul_ss[38]),
    .sel(mduinfo[2]),
    .o(n45[6]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b7 (
    .i0(n44[7]),
    .i1(mul_ss[39]),
    .sel(mduinfo[2]),
    .o(n45[7]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b8 (
    .i0(n44[8]),
    .i1(mul_ss[40]),
    .sel(mduinfo[2]),
    .o(n45[8]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux20_b9 (
    .i0(n44[9]),
    .i1(mul_ss[41]),
    .sel(mduinfo[2]),
    .o(n45[9]));  // ../RTL/core/exu_mdu.v(160)
  binary_mux_s1_w1 mux21_b0 (
    .i0(n45[0]),
    .i1(mul_ss[0]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[0]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b1 (
    .i0(n45[1]),
    .i1(mul_ss[1]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[1]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b10 (
    .i0(n45[10]),
    .i1(mul_ss[10]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[10]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b11 (
    .i0(n45[11]),
    .i1(mul_ss[11]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[11]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b12 (
    .i0(n45[12]),
    .i1(mul_ss[12]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[12]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b13 (
    .i0(n45[13]),
    .i1(mul_ss[13]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[13]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b14 (
    .i0(n45[14]),
    .i1(mul_ss[14]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[14]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b15 (
    .i0(n45[15]),
    .i1(mul_ss[15]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[15]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b16 (
    .i0(n45[16]),
    .i1(mul_ss[16]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[16]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b17 (
    .i0(n45[17]),
    .i1(mul_ss[17]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[17]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b18 (
    .i0(n45[18]),
    .i1(mul_ss[18]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[18]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b19 (
    .i0(n45[19]),
    .i1(mul_ss[19]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[19]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b2 (
    .i0(n45[2]),
    .i1(mul_ss[2]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[2]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b20 (
    .i0(n45[20]),
    .i1(mul_ss[20]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[20]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b21 (
    .i0(n45[21]),
    .i1(mul_ss[21]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[21]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b22 (
    .i0(n45[22]),
    .i1(mul_ss[22]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[22]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b23 (
    .i0(n45[23]),
    .i1(mul_ss[23]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[23]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b24 (
    .i0(n45[24]),
    .i1(mul_ss[24]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[24]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b25 (
    .i0(n45[25]),
    .i1(mul_ss[25]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[25]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b26 (
    .i0(n45[26]),
    .i1(mul_ss[26]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[26]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b27 (
    .i0(n45[27]),
    .i1(mul_ss[27]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[27]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b28 (
    .i0(n45[28]),
    .i1(mul_ss[28]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[28]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b29 (
    .i0(n45[29]),
    .i1(mul_ss[29]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[29]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b3 (
    .i0(n45[3]),
    .i1(mul_ss[3]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[3]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b30 (
    .i0(n45[30]),
    .i1(mul_ss[30]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[30]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b31 (
    .i0(n45[31]),
    .i1(mul_ss[31]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[31]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b4 (
    .i0(n45[4]),
    .i1(mul_ss[4]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[4]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b5 (
    .i0(n45[5]),
    .i1(mul_ss[5]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[5]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b6 (
    .i0(n45[6]),
    .i1(mul_ss[6]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[6]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b7 (
    .i0(n45[7]),
    .i1(mul_ss[7]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[7]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b8 (
    .i0(n45[8]),
    .i1(mul_ss[8]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[8]));  // ../RTL/core/exu_mdu.v(159)
  binary_mux_s1_w1 mux21_b9 (
    .i0(n45[9]),
    .i1(mul_ss[9]),
    .sel(mduinfo[1]),
    .o(o_mdu_rdwdata[9]));  // ../RTL/core/exu_mdu.v(159)
  and mux2_b0_sel_is_2 (mux2_b0_sel_is_2_o, i_rstn, mdu_vld);
  binary_mux_s1_w1 mux4_b0 (
    .i0(n19[0]),
    .i1(1'b0),
    .sel(n18),
    .o(n22[0]));  // ../RTL/core/exu_mdu.v(109)
  binary_mux_s1_w1 mux4_b1 (
    .i0(n19[1]),
    .i1(1'b0),
    .sel(n18),
    .o(n22[1]));  // ../RTL/core/exu_mdu.v(109)
  binary_mux_s1_w1 mux4_b2 (
    .i0(n19[2]),
    .i1(1'b0),
    .sel(n18),
    .o(n22[2]));  // ../RTL/core/exu_mdu.v(109)
  binary_mux_s1_w1 mux4_b3 (
    .i0(n19[3]),
    .i1(1'b0),
    .sel(n18),
    .o(n22[3]));  // ../RTL/core/exu_mdu.v(109)
  binary_mux_s1_w1 mux4_b4 (
    .i0(n19[4]),
    .i1(1'b0),
    .sel(n18),
    .o(n22[4]));  // ../RTL/core/exu_mdu.v(109)
  binary_mux_s1_w1 mux4_b5 (
    .i0(n19[5]),
    .i1(1'b0),
    .sel(n18),
    .o(n22[5]));  // ../RTL/core/exu_mdu.v(109)
  binary_mux_s1_w1 mux4_b6 (
    .i0(n19[6]),
    .i1(1'b0),
    .sel(n18),
    .o(n22[6]));  // ../RTL/core/exu_mdu.v(109)
  binary_mux_s1_w1 mux4_b7 (
    .i0(n19[7]),
    .i1(1'b0),
    .sel(n18),
    .o(n22[7]));  // ../RTL/core/exu_mdu.v(109)
  binary_mux_s1_w1 mux5_b0 (
    .i0(cnt[0]),
    .i1(n22[0]),
    .sel(mul_vld),
    .o(n25[0]));  // ../RTL/core/exu_mdu.v(108)
  binary_mux_s1_w1 mux5_b1 (
    .i0(cnt[1]),
    .i1(n22[1]),
    .sel(mul_vld),
    .o(n25[1]));  // ../RTL/core/exu_mdu.v(108)
  binary_mux_s1_w1 mux5_b2 (
    .i0(cnt[2]),
    .i1(n22[2]),
    .sel(mul_vld),
    .o(n25[2]));  // ../RTL/core/exu_mdu.v(108)
  binary_mux_s1_w1 mux5_b3 (
    .i0(cnt[3]),
    .i1(n22[3]),
    .sel(mul_vld),
    .o(n25[3]));  // ../RTL/core/exu_mdu.v(108)
  binary_mux_s1_w1 mux5_b4 (
    .i0(cnt[4]),
    .i1(n22[4]),
    .sel(mul_vld),
    .o(n25[4]));  // ../RTL/core/exu_mdu.v(108)
  binary_mux_s1_w1 mux5_b5 (
    .i0(cnt[5]),
    .i1(n22[5]),
    .sel(mul_vld),
    .o(n25[5]));  // ../RTL/core/exu_mdu.v(108)
  binary_mux_s1_w1 mux5_b6 (
    .i0(cnt[6]),
    .i1(n22[6]),
    .sel(mul_vld),
    .o(n25[6]));  // ../RTL/core/exu_mdu.v(108)
  binary_mux_s1_w1 mux5_b7 (
    .i0(cnt[7]),
    .i1(n22[7]),
    .sel(mul_vld),
    .o(n25[7]));  // ../RTL/core/exu_mdu.v(108)
  binary_mux_s1_w1 mux8_b0 (
    .i0(n25[0]),
    .i1(1'b0),
    .sel(mul_start),
    .o(n29[0]));  // ../RTL/core/exu_mdu.v(101)
  binary_mux_s1_w1 mux8_b1 (
    .i0(n25[1]),
    .i1(1'b0),
    .sel(mul_start),
    .o(n29[1]));  // ../RTL/core/exu_mdu.v(101)
  binary_mux_s1_w1 mux8_b2 (
    .i0(n25[2]),
    .i1(1'b0),
    .sel(mul_start),
    .o(n29[2]));  // ../RTL/core/exu_mdu.v(101)
  binary_mux_s1_w1 mux8_b3 (
    .i0(n25[3]),
    .i1(1'b0),
    .sel(mul_start),
    .o(n29[3]));  // ../RTL/core/exu_mdu.v(101)
  binary_mux_s1_w1 mux8_b4 (
    .i0(n25[4]),
    .i1(1'b0),
    .sel(mul_start),
    .o(n29[4]));  // ../RTL/core/exu_mdu.v(101)
  binary_mux_s1_w1 mux8_b5 (
    .i0(n25[5]),
    .i1(1'b0),
    .sel(mul_start),
    .o(n29[5]));  // ../RTL/core/exu_mdu.v(101)
  binary_mux_s1_w1 mux8_b6 (
    .i0(n25[6]),
    .i1(1'b0),
    .sel(mul_start),
    .o(n29[6]));  // ../RTL/core/exu_mdu.v(101)
  binary_mux_s1_w1 mux8_b7 (
    .i0(n25[7]),
    .i1(1'b0),
    .sel(mul_start),
    .o(n29[7]));  // ../RTL/core/exu_mdu.v(101)
  add_mu32_o32 neg0 (
    .i0(div_signed_rem),
    .o(n37));  // ../RTL/core/exu_mdu.v(165)
  AL_DFF_X rdwen_reg (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n6),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_will_rdwen));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg0_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_rdidx[0]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_will_rdidx[0]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg0_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_rdidx[1]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_mdu_rdidx[1]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg0_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_rdidx[2]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_mdu_rdidx[2]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg0_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_rdidx[3]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_will_rdidx[3]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg0_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_rdidx[4]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(o_will_rdidx[4]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg1_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mduinfo[1]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(mduinfo[1]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg1_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mduinfo[2]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(mduinfo[2]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg1_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mduinfo[3]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(mduinfo[3]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg1_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mduinfo[4]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(mduinfo[4]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg1_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mduinfo[5]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(mduinfo[5]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg1_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mduinfo[6]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(mduinfo[6]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg1_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mduinfo[7]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(mduinfo[7]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg1_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mduinfo[8]),
    .en(mux2_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(mduinfo[8]));  // ../RTL/core/exu_mdu.v(52)
  AL_DFF_X reg2_b0 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n29[0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(cnt[0]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg2_b1 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n29[1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(cnt[1]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg2_b2 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n29[2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(cnt[2]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg2_b3 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n29[3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(cnt[3]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg2_b4 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n29[4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(cnt[4]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg2_b5 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n29[5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(cnt[5]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg2_b6 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n29[6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(cnt[6]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg2_b7 (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n29[7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(cnt[7]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[0]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[0]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[1]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[1]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[10]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[10]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[11]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[11]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[12]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[12]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[13]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[13]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[14]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[14]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[15]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[15]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[16]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[16]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[17]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[17]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[18]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[18]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[19]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[19]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[2]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[2]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[20]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[20]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[21]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[21]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[22]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[22]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[23]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[23]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[24]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[24]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[25]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[25]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[26]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[26]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[27]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[27]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[28]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[28]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[29]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[29]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[3]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[3]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[30]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[30]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[31]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[31]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[4]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[4]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[5]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[5]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[6]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[6]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[7]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[7]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[8]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[8]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg3_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[9]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op1[9]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[0]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[0]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[1]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[1]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b10 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[10]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[10]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b11 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[11]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[11]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b12 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[12]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[12]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b13 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[13]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[13]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b14 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[14]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[14]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b15 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[15]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[15]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b16 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[16]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[16]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b17 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[17]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[17]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b18 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[18]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[18]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b19 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[19]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[19]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[2]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[2]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b20 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[20]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[20]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b21 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[21]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[21]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b22 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[22]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[22]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b23 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[23]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[23]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b24 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[24]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[24]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b25 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[25]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[25]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b26 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[26]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[26]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b27 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[27]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[27]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b28 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[28]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[28]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b29 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[29]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[29]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[3]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[3]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b30 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[30]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[30]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b31 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[31]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[31]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[4]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[4]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[5]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[5]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[6]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[6]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b7 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[7]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[7]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b8 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[8]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[8]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X reg4_b9 (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op2[9]),
    .en(mux10_b0_sel_is_2_o),
    .sr(1'b0),
    .ss(1'b0),
    .q(op2[9]));  // ../RTL/core/exu_mdu.v(96)
  AL_DFF_X rem_op1_sym_reg (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n10),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(rem_op1_sym));  // ../RTL/core/exu_mdu.v(52)
  AL_MUX u10 (
    .i0(working),
    .i1(1'b0),
    .sel(mdu_finish),
    .o(n4));  // ../RTL/core/exu_mdu.v(66)
  AL_MUX u11 (
    .i0(rem_op1_sym),
    .i1(1'b0),
    .sel(mdu_finish),
    .o(n5));  // ../RTL/core/exu_mdu.v(66)
  AL_MUX u12 (
    .i0(n3),
    .i1(i_mdu_rdwen),
    .sel(mdu_vld),
    .o(n6));  // ../RTL/core/exu_mdu.v(57)
  AL_MUX u13 (
    .i0(n4),
    .i1(1'b1),
    .sel(mdu_vld),
    .o(n8));  // ../RTL/core/exu_mdu.v(57)
  AL_MUX u14 (
    .i0(n5),
    .i1(i_mdu_op1[31]),
    .sel(mdu_vld),
    .o(n10));  // ../RTL/core/exu_mdu.v(57)
  and u16 (o_working, working, mdu_finish_neg);  // ../RTL/core/exu_mdu.v(76)
  or u18 (n14, i_mduinfo[1], i_mduinfo[2]);  // ../RTL/core/exu_mdu.v(94)
  or u19 (n15, n14, i_mduinfo[4]);  // ../RTL/core/exu_mdu.v(94)
  not u2 (n0, o_working);  // ../RTL/core/exu_mdu.v(47)
  or u20 (n16, n15, i_mduinfo[3]);  // ../RTL/core/exu_mdu.v(94)
  and u21 (mul_start, mdu_vld, n16);  // ../RTL/core/exu_mdu.v(93)
  AL_MUX u25 (
    .i0(mul_finish),
    .i1(1'b1),
    .sel(n18),
    .o(n20));  // ../RTL/core/exu_mdu.v(109)
  AL_MUX u28 (
    .i0(mul_vld),
    .i1(1'b0),
    .sel(u28_sel_is_3_o),
    .o(n24));
  and u28_sel_is_3 (u28_sel_is_3_o, mul_vld, n18);
  AL_MUX u29 (
    .i0(n24),
    .i1(1'b1),
    .sel(mul_start),
    .o(n26));  // ../RTL/core/exu_mdu.v(101)
  and u3 (n1, i_decinfo_grp[3], n0);  // ../RTL/core/exu_mdu.v(47)
  AL_MUX u30 (
    .i0(1'b0),
    .i1(n20),
    .sel(u30_sel_is_2_o),
    .o(n30));
  and u30_sel_is_2 (u30_sel_is_2_o, mul_start_neg, mul_vld);
  or u31 (n33, i_mduinfo[5], i_mduinfo[7]);  // ../RTL/core/exu_mdu.v(127)
  and u32 (div_signed_start, mdu_vld, n33);  // ../RTL/core/exu_mdu.v(127)
  or u34 (n36, i_mduinfo[6], i_mduinfo[8]);  // ../RTL/core/exu_mdu.v(142)
  and u35 (div_unsigned_start, mdu_vld, n36);  // ../RTL/core/exu_mdu.v(142)
  or u39 (div_finish, div_unsigned_finish, div_signed_finish);  // ../RTL/core/exu_mdu.v(153)
  and u4 (mdu_vld, n1, i_vld);  // ../RTL/core/exu_mdu.v(47)
  or u40 (mdu_finish, mul_finish, div_finish);  // ../RTL/core/exu_mdu.v(154)
  and u41 (o_mdu_rdwen, mdu_finish, o_will_rdwen);  // ../RTL/core/exu_mdu.v(156)
  AL_MUX u9 (
    .i0(1'b0),
    .i1(o_will_rdwen),
    .sel(u9_sel_is_0_o),
    .o(n3));
  and u9_sel_is_0 (u9_sel_is_0_o, mdu_finish_neg, i_flush_neg);
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F8880  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [8]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [9]));  // al_ip/div_signed_gate.v(4358)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F8990  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [14]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [15]));  // al_ip/div_signed_gate.v(4142)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F8AA0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [19]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [20]));  // al_ip/div_signed_gate.v(4196)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F8CC0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [20]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [21]));  // al_ip/div_signed_gate.v(4205)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F8DD0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [22]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [23]));  // al_ip/div_signed_gate.v(4223)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F8FF0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [18]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [19]));  // al_ip/div_signed_gate.v(4178)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F9210  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [0]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[0]));  // al_ip/div_signed_gate.v(4367)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F9430  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [11]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [12]));  // al_ip/div_signed_gate.v(4115)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F9540  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [23]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [24]));  // al_ip/div_signed_gate.v(4232)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F9650  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [15]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [16]));  // al_ip/div_signed_gate.v(4151)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F9760  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [24]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [25]));  // al_ip/div_signed_gate.v(4241)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F9BA0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [26]));  // al_ip/div_signed_gate.v(3962)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F9CB0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [1]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[1]));  // al_ip/div_signed_gate.v(4376)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F9DC0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [0]));  // al_ip/div_signed_gate.v(4079)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F9ED0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [0]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [1]));  // al_ip/div_signed_gate.v(4088)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66F9FE0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [3]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [4]));  // al_ip/div_signed_gate.v(4313)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FA0F0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [4]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [5]));  // al_ip/div_signed_gate.v(4322)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FA200  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [6]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [7]));  // al_ip/div_signed_gate.v(4340)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FA310  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [2]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[2]));  // al_ip/div_signed_gate.v(4475)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FA420  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [25]));  // al_ip/div_signed_gate.v(3953)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FA530  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [10]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [11]));  // al_ip/div_signed_gate.v(4106)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FA640  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [12]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [13]));  // al_ip/div_signed_gate.v(4124)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FA860  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [2]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [3]));  // al_ip/div_signed_gate.v(4286)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FAB90  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [27]));  // al_ip/div_signed_gate.v(3971)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FACA0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [5]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [6]));  // al_ip/div_signed_gate.v(4331)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FAFD0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [28]));  // al_ip/div_signed_gate.v(3980)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FB1F0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [9]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [10]));  // al_ip/div_signed_gate.v(4097)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FB300  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [13]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [14]));  // al_ip/div_signed_gate.v(4133)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FB410  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [16]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [17]));  // al_ip/div_signed_gate.v(4160)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FB630  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [17]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [18]));  // al_ip/div_signed_gate.v(4169)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FB740  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [21]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [22]));  // al_ip/div_signed_gate.v(4214)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u_DIV_SIGNED/al_00000256A66FB850  (
    .a(1'b0),
    .b(1'b0),
    .c(1'b0),
    .o({\u_DIV_SIGNED/al_00000256AA898580 ,open_n64}));  // al_ip/div_signed_gate.v(5232)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FBA70  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [31]));  // al_ip/div_signed_gate.v(4016)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FC2F0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [23]));  // al_ip/div_signed_gate.v(3935)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FC400  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [30]));  // al_ip/div_signed_gate.v(4007)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FC620  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [29]));  // al_ip/div_signed_gate.v(3989)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FC840  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [24]));  // al_ip/div_signed_gate.v(3944)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FCA60  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [1]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [2]));  // al_ip/div_signed_gate.v(4187)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FCB70  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [7]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [8]));  // al_ip/div_signed_gate.v(4349)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FE0B0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [15]));  // al_ip/div_signed_gate.v(3854)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FE3E0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [16]));  // al_ip/div_signed_gate.v(3863)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FE820  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [17]));  // al_ip/div_signed_gate.v(3872)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FEE80  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [18]));  // al_ip/div_signed_gate.v(3881)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FEF90  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [19]));  // al_ip/div_signed_gate.v(3890)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FF1B0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [20]));  // al_ip/div_signed_gate.v(3908)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FF700  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [21]));  // al_ip/div_signed_gate.v(3917)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FF810  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [22]));  // al_ip/div_signed_gate.v(3926)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FFB40  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [13]));  // al_ip/div_signed_gate.v(3836)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256A66FFD60  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [14]));  // al_ip/div_signed_gate.v(3845)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA39D160  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [25]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [26]));  // al_ip/div_signed_gate.v(4250)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A1780  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [26]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [27]));  // al_ip/div_signed_gate.v(4259)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A1AB0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [11]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [10]));  // al_ip/div_signed_gate.v(3242)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A1CD0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [12]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [11]));  // al_ip/div_signed_gate.v(3251)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A2110  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [17]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [16]));  // al_ip/div_signed_gate.v(3296)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A2550  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [1]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [0]));  // al_ip/div_signed_gate.v(3224)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A2990  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [14]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [13]));  // al_ip/div_signed_gate.v(3269)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A2AA0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [13]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [12]));  // al_ip/div_signed_gate.v(3260)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A2BB0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [18]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [17]));  // al_ip/div_signed_gate.v(3305)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A2CC0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [20]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [19]));  // al_ip/div_signed_gate.v(3323)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A2EE0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [3]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [2]));  // al_ip/div_signed_gate.v(3332)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A3100  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [21]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [20]));  // al_ip/div_signed_gate.v(3341)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A3210  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [4]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [3]));  // al_ip/div_signed_gate.v(3431)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A3320  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [8]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [7]));  // al_ip/div_signed_gate.v(3764)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A3540  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [15]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [14]));  // al_ip/div_signed_gate.v(3278)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A3650  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [22]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [21]));  // al_ip/div_signed_gate.v(3350)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A3760  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [23]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [22]));  // al_ip/div_signed_gate.v(3359)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A3870  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [25]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [24]));  // al_ip/div_signed_gate.v(3377)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A3980  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [9]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [8]));  // al_ip/div_signed_gate.v(3773)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A3ED0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [19]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [18]));  // al_ip/div_signed_gate.v(3314)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A3FE0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [26]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [25]));  // al_ip/div_signed_gate.v(3386)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A40F0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [27]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [26]));  // al_ip/div_signed_gate.v(3395)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A4200  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [28]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [27]));  // al_ip/div_signed_gate.v(3404)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A4310  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [29]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [28]));  // al_ip/div_signed_gate.v(3413)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A4420  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [6]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [5]));  // al_ip/div_signed_gate.v(3629)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A4530  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [30]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [29]));  // al_ip/div_signed_gate.v(3422)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A4640  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [31]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [30]));  // al_ip/div_signed_gate.v(3440)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A4750  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [31]));  // al_ip/div_signed_gate.v(3449)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A4860  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [7]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [6]));  // al_ip/div_signed_gate.v(3728)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A4970  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [16]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [15]));  // al_ip/div_signed_gate.v(3287)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A4A80  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [24]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [23]));  // al_ip/div_signed_gate.v(3368)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A4CA0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [32]));  // al_ip/div_signed_gate.v(3458)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A4DB0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [33]));  // al_ip/div_signed_gate.v(3467)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A50E0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [2]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [1]));  // al_ip/div_signed_gate.v(3233)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A5520  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [10]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [9]));  // al_ip/div_signed_gate.v(3782)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A5850  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [5]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [4]));  // al_ip/div_signed_gate.v(3530)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A5C90  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [29]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [30]));  // al_ip/div_signed_gate.v(4295)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A5DA0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [30]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [31]));  // al_ip/div_signed_gate.v(4304)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A5FC0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [3]));  // al_ip/div_signed_gate.v(3998)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A60D0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [7]));  // al_ip/div_signed_gate.v(4052)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A61E0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [39]));  // al_ip/div_signed_gate.v(3521)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A62F0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [61]));  // al_ip/div_signed_gate.v(3746)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A6510  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [10]));  // al_ip/div_signed_gate.v(3809)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A6620  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [11]));  // al_ip/div_signed_gate.v(3818)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A6730  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [55]));  // al_ip/div_signed_gate.v(3683)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A6840  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [56]));  // al_ip/div_signed_gate.v(3692)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A6950  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [43]));  // al_ip/div_signed_gate.v(3566)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A6A60  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [5]));  // al_ip/div_signed_gate.v(4034)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A6B70  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [8]));  // al_ip/div_signed_gate.v(4061)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A6C80  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [46]));  // al_ip/div_signed_gate.v(3593)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A6D90  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [12]));  // al_ip/div_signed_gate.v(3827)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A6EA0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [42]));  // al_ip/div_signed_gate.v(3557)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A6FB0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [41]));  // al_ip/div_signed_gate.v(3548)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A70C0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [60]));  // al_ip/div_signed_gate.v(3737)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A71D0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [48]));  // al_ip/div_signed_gate.v(3611)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A72E0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [36]));  // al_ip/div_signed_gate.v(3494)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A73F0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [47]));  // al_ip/div_signed_gate.v(3602)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A7500  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [54]));  // al_ip/div_signed_gate.v(3674)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A7610  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D7970 [62]),
    .en(1'b1),
    .sr(~div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [62]));  // al_ip/div_signed_gate.v(3755)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A7720  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [27]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [28]));  // al_ip/div_signed_gate.v(4268)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A7830  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [0]));  // al_ip/div_signed_gate.v(3791)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A7940  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [38]));  // al_ip/div_signed_gate.v(3512)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A7A50  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [57]));  // al_ip/div_signed_gate.v(3701)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A7B60  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [1]));  // al_ip/div_signed_gate.v(3800)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A7C70  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [45]));  // al_ip/div_signed_gate.v(3584)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A7D80  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [40]));  // al_ip/div_signed_gate.v(3539)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A7E90  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [50]));  // al_ip/div_signed_gate.v(3638)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A7FA0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [59]));  // al_ip/div_signed_gate.v(3719)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A80B0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [4]));  // al_ip/div_signed_gate.v(4025)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A81C0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [34]));  // al_ip/div_signed_gate.v(3476)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A82D0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [2]));  // al_ip/div_signed_gate.v(3899)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A83E0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [6]));  // al_ip/div_signed_gate.v(4043)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A84F0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [9]));  // al_ip/div_signed_gate.v(4070)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A8600  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [49]));  // al_ip/div_signed_gate.v(3620)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A8710  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [58]));  // al_ip/div_signed_gate.v(3710)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A8820  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [51]));  // al_ip/div_signed_gate.v(3647)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A8930  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [37]));  // al_ip/div_signed_gate.v(3503)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A8A40  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [52]));  // al_ip/div_signed_gate.v(3656)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A8B50  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [28]),
    .en(1'b1),
    .sr(div_signed_start),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [29]));  // al_ip/div_signed_gate.v(4277)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A8C60  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [44]));  // al_ip/div_signed_gate.v(3575)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A8D70  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [35]));  // al_ip/div_signed_gate.v(3485)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA3A8E80  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [53]));  // al_ip/div_signed_gate.v(3665)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47F090  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [0]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[0]));  // al_ip/div_signed_gate.v(4655)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47F1A0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [3]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[3]));  // al_ip/div_signed_gate.v(4862)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47F2B0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [9]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[9]));  // al_ip/div_signed_gate.v(4646)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47F3C0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [17]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[17]));  // al_ip/div_signed_gate.v(4736)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47F4D0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [19]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[19]));  // al_ip/div_signed_gate.v(4754)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47F5E0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [6]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[6]));  // al_ip/div_signed_gate.v(4619)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47F6F0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D38B0 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CE7C0 [1]));  // al_ip/div_signed_gate.v(4952)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47F800  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [13]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[13]));  // al_ip/div_signed_gate.v(4412)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47F910  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [6]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[6]));  // al_ip/div_signed_gate.v(4907)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47FA20  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [26]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[26]));  // al_ip/div_signed_gate.v(4826)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47FB30  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [27]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[27]));  // al_ip/div_signed_gate.v(4547)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47FC40  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [30]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[30]));  // al_ip/div_signed_gate.v(4583)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47FD50  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [11]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[11]));  // al_ip/div_signed_gate.v(4682)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47FE60  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [12]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[12]));  // al_ip/div_signed_gate.v(4691)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA47FF70  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [20]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[20]));  // al_ip/div_signed_gate.v(4772)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA480080  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [5]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[5]));  // al_ip/div_signed_gate.v(4610)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA480190  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [14]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[14]));  // al_ip/div_signed_gate.v(4421)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4802A0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [7]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[7]));  // al_ip/div_signed_gate.v(4916)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4803B0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [10]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[10]));  // al_ip/div_signed_gate.v(4673)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4804C0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [23]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[23]));  // al_ip/div_signed_gate.v(4799)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4805D0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [26]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[26]));  // al_ip/div_signed_gate.v(4538)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4806E0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [3]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[3]));  // al_ip/div_signed_gate.v(4574)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4807F0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [29]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[29]));  // al_ip/div_signed_gate.v(4565)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA480900  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [28]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[28]));  // al_ip/div_signed_gate.v(4556)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA480A10  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D38B0 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CE7C0 [2]));  // al_ip/div_signed_gate.v(4961)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA480B20  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [14]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[14]));  // al_ip/div_signed_gate.v(4709)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA480C30  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [13]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[13]));  // al_ip/div_signed_gate.v(4700)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA480D40  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [16]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[16]));  // al_ip/div_signed_gate.v(4727)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA480E50  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [8]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[8]));  // al_ip/div_signed_gate.v(4925)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA480F60  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [21]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[21]));  // al_ip/div_signed_gate.v(4781)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA481070  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [24]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[24]));  // al_ip/div_signed_gate.v(4520)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA481180  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [11]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[11]));  // al_ip/div_signed_gate.v(4394)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA481290  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D38B0 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CE7C0 [3]));  // al_ip/div_signed_gate.v(4970)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4813A0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [5]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[5]));  // al_ip/div_signed_gate.v(4898)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4814B0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [9]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[9]));  // al_ip/div_signed_gate.v(4934)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4815C0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [18]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[18]));  // al_ip/div_signed_gate.v(4745)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4816D0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [7]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[7]));  // al_ip/div_signed_gate.v(4628)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4817E0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D38B0 [4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CE7C0 [4]));  // al_ip/div_signed_gate.v(4979)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4818F0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [22]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[22]));  // al_ip/div_signed_gate.v(4790)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA481A00  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D38B0 [5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CE7C0 [5]));  // al_ip/div_signed_gate.v(4988)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA481B10  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [4]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[4]));  // al_ip/div_signed_gate.v(4601)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA481C20  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [15]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[15]));  // al_ip/div_signed_gate.v(4718)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA481D30  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [8]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[8]));  // al_ip/div_signed_gate.v(4637)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA481E40  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [17]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[17]));  // al_ip/div_signed_gate.v(4448)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA481F50  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [20]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[20]));  // al_ip/div_signed_gate.v(4484)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA482060  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [16]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[16]));  // al_ip/div_signed_gate.v(4439)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA482170  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [23]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[23]));  // al_ip/div_signed_gate.v(4511)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA482390  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [12]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[12]));  // al_ip/div_signed_gate.v(4403)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4824A0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [15]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[15]));  // al_ip/div_signed_gate.v(4430)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4825B0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [4]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[4]));  // al_ip/div_signed_gate.v(4889)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4826C0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [24]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[24]));  // al_ip/div_signed_gate.v(4808)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4827D0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [31]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[31]));  // al_ip/div_signed_gate.v(4592)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4828E0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [25]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[25]));  // al_ip/div_signed_gate.v(4817)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA4829F0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [27]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[27]));  // al_ip/div_signed_gate.v(4835)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA482B00  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [18]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[18]));  // al_ip/div_signed_gate.v(4457)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA482C10  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [21]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[21]));  // al_ip/div_signed_gate.v(4493)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA482D20  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [22]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[22]));  // al_ip/div_signed_gate.v(4502)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA482E30  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [25]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[25]));  // al_ip/div_signed_gate.v(4529)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA482F40  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D38B0 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA0CE7C0 [0]));  // al_ip/div_signed_gate.v(4943)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA483050  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [19]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[19]));  // al_ip/div_signed_gate.v(4466)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA483160  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [1]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[1]));  // al_ip/div_signed_gate.v(4664)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA483270  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [2]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[2]));  // al_ip/div_signed_gate.v(4763)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA483380  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [10]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_quo[10]));  // al_ip/div_signed_gate.v(4385)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA483AF0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [30]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[30]));  // al_ip/div_signed_gate.v(4871)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA484150  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [28]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[28]));  // al_ip/div_signed_gate.v(4844)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA485BE0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [29]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[29]));  // al_ip/div_signed_gate.v(4853)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA486570  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [31]),
    .en(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_rem[31]));  // al_ip/div_signed_gate.v(4880)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_SIGNED/al_00000256AA4D31A0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .b(\u_DIV_SIGNED/al_00000256AA8940C0 ),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D29D0 [2]),
    .o(\u_DIV_SIGNED/al_00000256AA0D38B0 [2]));  // al_ip/div_signed_gate.v(975)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_SIGNED/al_00000256AA4D4A10  (
    .a(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .b(\u_DIV_SIGNED/al_00000256AA8940C0 ),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D29D0 [5]),
    .o(\u_DIV_SIGNED/al_00000256AA0D38B0 [5]));  // al_ip/div_signed_gate.v(948)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_SIGNED/al_00000256AA4D4B20  (
    .a(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .b(\u_DIV_SIGNED/al_00000256AA8940C0 ),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D29D0 [1]),
    .o(\u_DIV_SIGNED/al_00000256AA0D38B0 [1]));  // al_ip/div_signed_gate.v(984)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_SIGNED/al_00000256AA4D4E50  (
    .a(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .b(\u_DIV_SIGNED/al_00000256AA8940C0 ),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D29D0 [3]),
    .o(\u_DIV_SIGNED/al_00000256AA0D38B0 [3]));  // al_ip/div_signed_gate.v(966)
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'b0001))
    \u_DIV_SIGNED/al_00000256AA4D58F0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CE7C0 [1]),
    .b(\u_DIV_SIGNED/al_00000256AA0CE7C0 [2]),
    .o(\u_DIV_SIGNED/al_00000256AA895350 ));  // al_ip/div_signed_gate.v(921)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_SIGNED/al_00000256AA4D5E40  (
    .a(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .b(\u_DIV_SIGNED/al_00000256AA8940C0 ),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D29D0 [4]),
    .o(\u_DIV_SIGNED/al_00000256AA0D38B0 [4]));  // al_ip/div_signed_gate.v(957)
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~B*~A))"),
    .INIT(16'b1111000111110000))
    \u_DIV_SIGNED/al_00000256AA4D5F50  (
    .a(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .b(\u_DIV_SIGNED/al_00000256AA8940C0 ),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D29D0 [0]),
    .o(\u_DIV_SIGNED/al_00000256AA0D38B0 [0]));  // al_ip/div_signed_gate.v(1001)
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'b00000000000000000000000000000010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4D6280  (
    .a(\u_DIV_SIGNED/al_00000256AA895350 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CE7C0 [0]),
    .c(\u_DIV_SIGNED/al_00000256AA0CE7C0 [3]),
    .d(\u_DIV_SIGNED/al_00000256AA0CE7C0 [4]),
    .e(\u_DIV_SIGNED/al_00000256AA0CE7C0 [5]),
    .o(\u_DIV_SIGNED/al_00000256AA8940C0 ));  // al_ip/div_signed_gate.v(938)
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'b00000000000010000000000000000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4D6390  (
    .a(\u_DIV_SIGNED/al_00000256AA895350 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CE7C0 [0]),
    .c(\u_DIV_SIGNED/al_00000256AA0CE7C0 [3]),
    .d(\u_DIV_SIGNED/al_00000256AA0CE7C0 [4]),
    .e(\u_DIV_SIGNED/al_00000256AA0CE7C0 [5]),
    .o(\u_DIV_SIGNED/al_00000256AA3DD9A0 ));  // al_ip/div_signed_gate.v(928)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4D6D20  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [9]),
    .b(n35[31]),
    .c(n35[9]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [9]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [9]));  // al_ip/div_signed_gate.v(911)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D7490  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [17]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [17]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [17]));  // al_ip/div_signed_gate.v(1353)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D75A0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [28]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [28]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [28]));  // al_ip/div_signed_gate.v(1065)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D76B0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [5]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [5]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [5]));  // al_ip/div_signed_gate.v(1121)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D77C0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [14]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [14]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [14]));  // al_ip/div_signed_gate.v(1385)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D78D0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [7]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [7]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [7]));  // al_ip/div_signed_gate.v(1177)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D79E0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [10]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [10]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [10]));  // al_ip/div_signed_gate.v(1417)
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'b0110))
    \u_DIV_SIGNED/al_00000256AA4D7AF0  (
    .a(n34[31]),
    .b(n35[31]),
    .o(\u_DIV_SIGNED/al_00000256AA422680 ));  // al_ip/div_signed_gate.v(301)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D7C00  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [31]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [31]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [31]));  // al_ip/div_signed_gate.v(1097)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D7D10  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [0]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [0]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [0]));  // al_ip/div_signed_gate.v(1113)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D7E20  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [9]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [9]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [9]));  // al_ip/div_signed_gate.v(1153)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D7F30  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [21]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [21]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [21]));  // al_ip/div_signed_gate.v(1313)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D8040  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [20]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [20]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [20]));  // al_ip/div_signed_gate.v(1321)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D8150  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [13]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [13]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [13]));  // al_ip/div_signed_gate.v(1393)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D8260  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [13]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [13]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [13]));  // al_ip/div_signed_gate.v(1579)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D8370  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [30]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [30]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [30]));  // al_ip/div_signed_gate.v(1225)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D8480  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [25]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [25]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [25]));  // al_ip/div_signed_gate.v(1273)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D8590  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [26]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [26]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [26]));  // al_ip/div_signed_gate.v(1049)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D86A0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [24]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [24]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [24]));  // al_ip/div_signed_gate.v(1281)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D87B0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [2]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [2]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [2]));  // al_ip/div_signed_gate.v(1329)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D88C0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [12]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [12]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [12]));  // al_ip/div_signed_gate.v(1401)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D89D0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [23]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [23]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [23]));  // al_ip/div_signed_gate.v(1018)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D8AE0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [4]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [4]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [4]));  // al_ip/div_signed_gate.v(1105)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D8BF0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [8]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [8]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [8]));  // al_ip/div_signed_gate.v(1169)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D8D00  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [9]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [9]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [9]));  // al_ip/div_signed_gate.v(1161)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'b1000))
    \u_DIV_SIGNED/al_00000256AA4D8E10  (
    .a(n34[31]),
    .b(\u_DIV_SIGNED/al_00000256AA0D5590 [31]),
    .o(\u_DIV_SIGNED/al_00000256AA0D7970 [62]));  // al_ip/div_signed_gate.v(1026)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D8F20  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [16]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [16]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [16]));  // al_ip/div_signed_gate.v(406)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9030  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [18]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [18]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [18]));  // al_ip/div_signed_gate.v(602)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9140  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [19]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [19]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [19]));  // al_ip/div_signed_gate.v(700)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9250  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [25]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [25]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [25]));  // al_ip/div_signed_gate.v(1041)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9360  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [27]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [27]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [27]));  // al_ip/div_signed_gate.v(1057)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9470  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [1]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [1]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [1]));  // al_ip/div_signed_gate.v(1201)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9580  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [17]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [17]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [17]));  // al_ip/div_signed_gate.v(504)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9690  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [2]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [2]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [2]));  // al_ip/div_signed_gate.v(797)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D97A0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [24]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [24]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [24]));  // al_ip/div_signed_gate.v(1033)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D98B0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [6]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [6]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [6]));  // al_ip/div_signed_gate.v(1185)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D99C0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [31]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [31]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [31]));  // al_ip/div_signed_gate.v(1217)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9AD0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [14]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [14]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [14]));  // al_ip/div_signed_gate.v(1687)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D9BE0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [3]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [3]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [3]));  // al_ip/div_signed_gate.v(1233)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D9CF0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [28]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [28]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [28]));  // al_ip/div_signed_gate.v(1249)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D9E00  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [27]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [27]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [27]));  // al_ip/div_signed_gate.v(1257)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D9F10  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [23]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [23]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [23]));  // al_ip/div_signed_gate.v(1297)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DA020  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [26]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [26]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [26]));  // al_ip/div_signed_gate.v(1265)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DA130  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [22]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [22]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [22]));  // al_ip/div_signed_gate.v(1305)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DA240  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [7]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [7]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [7]));  // al_ip/div_signed_gate.v(1137)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DA350  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [19]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [19]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [19]));  // al_ip/div_signed_gate.v(1337)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DA460  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [3]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [3]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [3]));  // al_ip/div_signed_gate.v(1081)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DA570  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [30]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [30]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [30]));  // al_ip/div_signed_gate.v(1089)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DA680  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [5]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [5]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [5]));  // al_ip/div_signed_gate.v(1193)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DA790  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [22]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [22]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [22]));  // al_ip/div_signed_gate.v(1010)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DA8A0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [18]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [18]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [18]));  // al_ip/div_signed_gate.v(1345)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DA9B0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [15]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [15]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [15]));  // al_ip/div_signed_gate.v(308)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DAAC0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [16]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [16]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [16]));  // al_ip/div_signed_gate.v(1361)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DABD0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [29]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [29]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [29]));  // al_ip/div_signed_gate.v(1073)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DACE0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [12]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [12]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [12]));  // al_ip/div_signed_gate.v(1471)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DADF0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [11]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [11]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [11]));  // al_ip/div_signed_gate.v(1377)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DAF00  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [8]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [8]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [8]));  // al_ip/div_signed_gate.v(1145)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DB010  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [20]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [20]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [20]));  // al_ip/div_signed_gate.v(895)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DB120  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [4]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [4]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [4]));  // al_ip/div_signed_gate.v(1209)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DB230  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [21]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [21]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [21]));  // al_ip/div_signed_gate.v(993)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DB340  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [29]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [29]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [29]));  // al_ip/div_signed_gate.v(1241)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DB450  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [15]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [15]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [15]));  // al_ip/div_signed_gate.v(1369)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DB560  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [11]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [11]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [11]));  // al_ip/div_signed_gate.v(1409)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DB670  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [10]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [10]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [10]));  // al_ip/div_signed_gate.v(1289)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DB780  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [6]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [6]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [6]));  // al_ip/div_signed_gate.v(1129)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DB890  (
    .a(n34[31]),
    .b(n34[5]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [5]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [37]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [36]));  // al_ip/div_signed_gate.v(1725)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DB9A0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [10]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [10]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [10]));  // al_ip/div_signed_gate.v(334)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DBAB0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [14]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [14]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [14]));  // al_ip/div_signed_gate.v(414)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DBBC0  (
    .a(n34[31]),
    .b(n34[15]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [15]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [47]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [46]));  // al_ip/div_signed_gate.v(1519)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DBCD0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [20]),
    .b(n35[31]),
    .c(n35[20]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [20]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [20]));  // al_ip/div_signed_gate.v(556)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DBDE0  (
    .a(n34[31]),
    .b(n34[29]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [29]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [61]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [60]));  // al_ip/div_signed_gate.v(1677)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DBEF0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [16]),
    .b(n35[31]),
    .c(n35[16]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [16]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [16]));  // al_ip/div_signed_gate.v(458)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DC000  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [17]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [17]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [17]));  // al_ip/div_signed_gate.v(468)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DC110  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [19]),
    .b(n35[31]),
    .c(n35[19]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [19]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [19]));  // al_ip/div_signed_gate.v(520)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DC220  (
    .a(n34[31]),
    .b(n34[30]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [30]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [62]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [61]));  // al_ip/div_signed_gate.v(1705)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DC330  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [2]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [2]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [2]));  // al_ip/div_signed_gate.v(530)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DC440  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [20]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [20]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [20]));  // al_ip/div_signed_gate.v(548)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DC550  (
    .a(n34[31]),
    .b(n34[11]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [11]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [43]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [42]));  // al_ip/div_signed_gate.v(1479)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DC660  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [0]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [0]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [0]));  // al_ip/div_signed_gate.v(1775)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DC770  (
    .a(n34[31]),
    .b(n34[1]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [1]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [33]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [32]));  // al_ip/div_signed_gate.v(1451)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DC880  (
    .a(n34[31]),
    .b(n34[8]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [8]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [40]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [39]));  // al_ip/div_signed_gate.v(1755)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DC990  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [15]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [15]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [15]));  // al_ip/div_signed_gate.v(432)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DCAA0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [21]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [21]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [21]));  // al_ip/div_signed_gate.v(566)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DCBB0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [21]),
    .b(n35[31]),
    .c(n35[21]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [21]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [21]));  // al_ip/div_signed_gate.v(574)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DCCC0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [22]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [22]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [22]));  // al_ip/div_signed_gate.v(584)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DCDD0  (
    .a(n34[31]),
    .b(n34[12]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [12]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [44]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [43]));  // al_ip/div_signed_gate.v(1489)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DCEE0  (
    .a(n34[31]),
    .b(n34[10]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [10]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [42]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [41]));  // al_ip/div_signed_gate.v(1461)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DCFF0  (
    .a(n34[31]),
    .b(n34[16]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [16]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [48]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [47]));  // al_ip/div_signed_gate.v(1529)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DD100  (
    .a(n34[31]),
    .b(n34[18]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [18]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [50]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [49]));  // al_ip/div_signed_gate.v(1549)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DD210  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [12]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [12]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [12]));  // al_ip/div_signed_gate.v(370)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DD320  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [1]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [1]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [1]));  // al_ip/div_signed_gate.v(1425)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DD430  (
    .a(n34[31]),
    .b(n34[27]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [27]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [59]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [58]));  // al_ip/div_signed_gate.v(1657)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DD540  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [0]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [0]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [0]));  // al_ip/div_signed_gate.v(1433)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DD650  (
    .a(n34[31]),
    .b(n34[3]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [3]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [35]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [34]));  // al_ip/div_signed_gate.v(1695)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DD760  (
    .a(n34[31]),
    .b(n34[7]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [7]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [39]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [38]));  // al_ip/div_signed_gate.v(1745)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DD870  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [0]),
    .b(n35[31]),
    .c(n35[0]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [0]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [0]));  // al_ip/div_signed_gate.v(1783)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DD980  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [10]),
    .b(n35[31]),
    .c(n35[10]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [10]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [10]));  // al_ip/div_signed_gate.v(342)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DDA90  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [1]),
    .b(n35[31]),
    .c(n35[1]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [1]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [1]));  // al_ip/div_signed_gate.v(324)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DDBA0  (
    .a(n34[31]),
    .b(n34[13]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [13]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [45]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [44]));  // al_ip/div_signed_gate.v(1499)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DDCB0  (
    .a(n34[31]),
    .b(n34[6]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [6]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [38]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [37]));  // al_ip/div_signed_gate.v(1735)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DDDC0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [11]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [11]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [11]));  // al_ip/div_signed_gate.v(352)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DDED0  (
    .a(n34[31]),
    .b(n34[14]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [14]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [46]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [45]));  // al_ip/div_signed_gate.v(1509)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DDFE0  (
    .a(n34[31]),
    .b(n34[17]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [17]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [49]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [48]));  // al_ip/div_signed_gate.v(1539)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE0F0  (
    .a(n34[31]),
    .b(n34[25]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [25]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [57]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [56]));  // al_ip/div_signed_gate.v(1637)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE200  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [12]),
    .b(n35[31]),
    .c(n35[12]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [12]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [12]));  // al_ip/div_signed_gate.v(378)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DE310  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [13]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [13]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [13]));  // al_ip/div_signed_gate.v(388)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE420  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [14]),
    .b(n35[31]),
    .c(n35[14]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [14]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [14]));  // al_ip/div_signed_gate.v(422)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DE530  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [18]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [18]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [18]));  // al_ip/div_signed_gate.v(486)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE640  (
    .a(n34[31]),
    .b(n34[0]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [0]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [32]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [31]));  // al_ip/div_signed_gate.v(1441)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE750  (
    .a(n34[31]),
    .b(n34[19]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [19]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [51]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [50]));  // al_ip/div_signed_gate.v(1559)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE860  (
    .a(n34[31]),
    .b(n34[2]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [2]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [34]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [33]));  // al_ip/div_signed_gate.v(1569)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE970  (
    .a(n34[31]),
    .b(n34[21]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [21]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [53]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [52]));  // al_ip/div_signed_gate.v(1597)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DEA80  (
    .a(n34[31]),
    .b(n34[23]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [23]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [55]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [54]));  // al_ip/div_signed_gate.v(1617)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DEB90  (
    .a(n34[31]),
    .b(n34[22]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [22]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [54]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [53]));  // al_ip/div_signed_gate.v(1607)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DECA0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [1]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [1]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [1]));  // al_ip/div_signed_gate.v(316)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DEDB0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [11]),
    .b(n35[31]),
    .c(n35[11]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [11]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [11]));  // al_ip/div_signed_gate.v(360)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DEEC0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [15]),
    .b(n35[31]),
    .c(n35[15]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [15]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [15]));  // al_ip/div_signed_gate.v(440)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DEFD0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [16]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [16]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [16]));  // al_ip/div_signed_gate.v(450)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF0E0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [17]),
    .b(n35[31]),
    .c(n35[17]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [17]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [17]));  // al_ip/div_signed_gate.v(476)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF1F0  (
    .a(n34[31]),
    .b(n34[24]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [24]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [56]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [55]));  // al_ip/div_signed_gate.v(1627)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF300  (
    .a(n34[31]),
    .b(n34[4]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [4]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [36]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [35]));  // al_ip/div_signed_gate.v(1715)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF410  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [18]),
    .b(n35[31]),
    .c(n35[18]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [18]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [18]));  // al_ip/div_signed_gate.v(494)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF520  (
    .a(n34[31]),
    .b(n34[28]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [28]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [60]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [59]));  // al_ip/div_signed_gate.v(1667)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF630  (
    .a(n34[31]),
    .b(n34[9]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [9]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [41]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [40]));  // al_ip/div_signed_gate.v(1765)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF740  (
    .a(n34[31]),
    .b(n34[20]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [20]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [52]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [51]));  // al_ip/div_signed_gate.v(1587)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF850  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [13]),
    .b(n35[31]),
    .c(n35[13]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [13]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [13]));  // al_ip/div_signed_gate.v(396)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DF960  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [19]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [19]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [19]));  // al_ip/div_signed_gate.v(512)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DFA70  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [2]),
    .b(n35[31]),
    .c(n35[2]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [2]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [2]));  // al_ip/div_signed_gate.v(538)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DFB80  (
    .a(n34[31]),
    .b(n34[26]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [26]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [58]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [57]));  // al_ip/div_signed_gate.v(1647)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DFC90  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [24]),
    .b(n35[31]),
    .c(n35[24]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [24]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [24]));  // al_ip/div_signed_gate.v(636)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DFDA0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [26]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [26]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [26]));  // al_ip/div_signed_gate.v(664)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DFEB0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [27]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [27]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [27]));  // al_ip/div_signed_gate.v(682)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DFFC0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [30]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [30]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [30]));  // al_ip/div_signed_gate.v(762)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E00D0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [29]),
    .b(n35[31]),
    .c(n35[29]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [29]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [29]));  // al_ip/div_signed_gate.v(734)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E02F0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [28]),
    .b(n35[31]),
    .c(n35[28]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [28]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [28]));  // al_ip/div_signed_gate.v(716)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0400  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [25]),
    .b(n35[31]),
    .c(n35[25]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [25]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [25]));  // al_ip/div_signed_gate.v(654)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E0620  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [28]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [28]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [28]));  // al_ip/div_signed_gate.v(708)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E0730  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [3]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [3]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [3]));  // al_ip/div_signed_gate.v(744)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0840  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [30]),
    .b(n35[31]),
    .c(n35[30]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [30]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [30]));  // al_ip/div_signed_gate.v(770)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0950  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [3]),
    .b(n35[31]),
    .c(n35[3]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [3]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [3]));  // al_ip/div_signed_gate.v(752)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E0A60  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [4]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [4]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [4]));  // al_ip/div_signed_gate.v(805)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0B70  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [4]),
    .b(n35[31]),
    .c(n35[4]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [4]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [4]));  // al_ip/div_signed_gate.v(813)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0C80  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [5]),
    .b(n35[31]),
    .c(n35[5]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [5]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [5]));  // al_ip/div_signed_gate.v(831)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0D90  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [6]),
    .b(n35[31]),
    .c(n35[6]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [6]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [6]));  // al_ip/div_signed_gate.v(849)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0EA0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [7]),
    .b(n35[31]),
    .c(n35[7]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [7]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [7]));  // al_ip/div_signed_gate.v(867)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E0FB0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [8]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [8]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [8]));  // al_ip/div_signed_gate.v(877)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E10C0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [9]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [9]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [9]));  // al_ip/div_signed_gate.v(903)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E11D0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [8]),
    .b(n35[31]),
    .c(n35[8]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [8]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [8]));  // al_ip/div_signed_gate.v(885)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E12E0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [29]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [29]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [29]));  // al_ip/div_signed_gate.v(726)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E13F0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [23]),
    .b(n35[31]),
    .c(n35[23]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [23]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [23]));  // al_ip/div_signed_gate.v(618)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E1500  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [26]),
    .b(n35[31]),
    .c(n35[26]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [26]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [26]));  // al_ip/div_signed_gate.v(672)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E1610  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [5]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [5]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [5]));  // al_ip/div_signed_gate.v(823)
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*B))*~(C)+~A*(D*B)*~(C)+~(~A)*(D*B)*C+~A*(D*B)*C)"),
    .INIT(16'b1100010100000101))
    \u_DIV_SIGNED/al_00000256AA4E1720  (
    .a(\u_DIV_SIGNED/al_00000256AA893670 ),
    .b(n35[31]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA3FF0F0 [31]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [31]));  // al_ip/div_signed_gate.v(788)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E1830  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [6]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [6]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [6]));  // al_ip/div_signed_gate.v(841)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E1B60  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [7]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [7]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [7]));  // al_ip/div_signed_gate.v(859)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E1D80  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [23]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [23]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [23]));  // al_ip/div_signed_gate.v(610)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E20B0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [25]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [25]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [25]));  // al_ip/div_signed_gate.v(646)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E21C0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [27]),
    .b(n35[31]),
    .c(n35[27]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [27]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [27]));  // al_ip/div_signed_gate.v(690)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E22D0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [24]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [24]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [24]));  // al_ip/div_signed_gate.v(628)
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b00011011))
    \u_DIV_SIGNED/al_00000256AA4E2710  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [31]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [31]),
    .o(\u_DIV_SIGNED/al_00000256AA893670 ));  // al_ip/div_signed_gate.v(780)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E2B50  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [22]),
    .b(n35[31]),
    .c(n35[22]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [22]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [22]));  // al_ip/div_signed_gate.v(592)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6690A0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [18]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [18]),
    .c(\u_DIV_SIGNED/al_00000256AA8994A0 ),
    .o({\u_DIV_SIGNED/al_00000256AA898DC0 ,\u_DIV_SIGNED/al_00000256AA400D60 [18]}));  // al_ip/div_signed_gate.v(5078)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6691B0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [23]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [23]),
    .c(\u_DIV_SIGNED/al_00000256AA898E70 ),
    .o({\u_DIV_SIGNED/al_00000256AA899340 ,\u_DIV_SIGNED/al_00000256AA400D60 [23]}));  // al_ip/div_signed_gate.v(5120)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6692C0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [25]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [25]),
    .c(\u_DIV_SIGNED/al_00000256AA898D10 ),
    .o({\u_DIV_SIGNED/al_00000256AA898F20 ,\u_DIV_SIGNED/al_00000256AA400D60 [25]}));  // al_ip/div_signed_gate.v(5134)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6693D0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [26]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [26]),
    .c(\u_DIV_SIGNED/al_00000256AA898F20 ),
    .o({\u_DIV_SIGNED/al_00000256AA898630 ,\u_DIV_SIGNED/al_00000256AA400D60 [26]}));  // al_ip/div_signed_gate.v(5141)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6694E0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [22]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [22]),
    .c(\u_DIV_SIGNED/al_00000256AA89ACB0 ),
    .o({\u_DIV_SIGNED/al_00000256AA898E70 ,\u_DIV_SIGNED/al_00000256AA400D60 [22]}));  // al_ip/div_signed_gate.v(5113)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6695F0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [27]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [27]),
    .c(\u_DIV_SIGNED/al_00000256AA898630 ),
    .o({\u_DIV_SIGNED/al_00000256AA899550 ,\u_DIV_SIGNED/al_00000256AA400D60 [27]}));  // al_ip/div_signed_gate.v(5148)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA669700  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [16]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [16]),
    .c(\u_DIV_SIGNED/al_00000256AA89A520 ),
    .o({\u_DIV_SIGNED/al_00000256AA8988F0 ,\u_DIV_SIGNED/al_00000256AA400D60 [16]}));  // al_ip/div_signed_gate.v(5064)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA669810  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [2]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [2]),
    .c(\u_DIV_SIGNED/al_00000256AA899760 ),
    .o({\u_DIV_SIGNED/al_00000256AA898FD0 ,\u_DIV_SIGNED/al_00000256AA400D60 [2]}));  // al_ip/div_signed_gate.v(5092)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA669920  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [14]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [14]),
    .c(\u_DIV_SIGNED/al_00000256AA8993F0 ),
    .o({\u_DIV_SIGNED/al_00000256AA899130 ,\u_DIV_SIGNED/al_00000256AA400D60 [14]}));  // al_ip/div_signed_gate.v(5050)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA669A30  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [28]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [28]),
    .c(\u_DIV_SIGNED/al_00000256AA899550 ),
    .o({\u_DIV_SIGNED/al_00000256AA8986E0 ,\u_DIV_SIGNED/al_00000256AA400D60 [28]}));  // al_ip/div_signed_gate.v(5155)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA669B40  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [29]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [29]),
    .c(\u_DIV_SIGNED/al_00000256AA8986E0 ),
    .o({\u_DIV_SIGNED/al_00000256AA899600 ,\u_DIV_SIGNED/al_00000256AA400D60 [29]}));  // al_ip/div_signed_gate.v(5162)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA669D60  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [12]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [12]),
    .c(\u_DIV_SIGNED/al_00000256AA899970 ),
    .o({\u_DIV_SIGNED/al_00000256AA8996B0 ,\u_DIV_SIGNED/al_00000256AA400D60 [12]}));  // al_ip/div_signed_gate.v(5036)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66A090  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [3]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [3]),
    .c(\u_DIV_SIGNED/al_00000256AA898FD0 ),
    .o({\u_DIV_SIGNED/al_00000256AA8998C0 ,\u_DIV_SIGNED/al_00000256AA400D60 [3]}));  // al_ip/div_signed_gate.v(5169)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA66A1A0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_signed_finish));  // al_ip/div_signed_gate.v(2753)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66A3C0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [30]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [30]),
    .c(\u_DIV_SIGNED/al_00000256AA899600 ),
    .o({\u_DIV_SIGNED/al_00000256AA899810 ,\u_DIV_SIGNED/al_00000256AA400D60 [30]}));  // al_ip/div_signed_gate.v(5176)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66A800  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [15]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [15]),
    .c(\u_DIV_SIGNED/al_00000256AA899130 ),
    .o({\u_DIV_SIGNED/al_00000256AA89A520 ,\u_DIV_SIGNED/al_00000256AA400D60 [15]}));  // al_ip/div_signed_gate.v(5057)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66AD50  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [19]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [19]),
    .c(\u_DIV_SIGNED/al_00000256AA898DC0 ),
    .o({\u_DIV_SIGNED/al_00000256AA89AC00 ,\u_DIV_SIGNED/al_00000256AA400D60 [19]}));  // al_ip/div_signed_gate.v(5085)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66AF70  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [20]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [20]),
    .c(\u_DIV_SIGNED/al_00000256AA89AC00 ),
    .o({\u_DIV_SIGNED/al_00000256AA89A260 ,\u_DIV_SIGNED/al_00000256AA400D60 [20]}));  // al_ip/div_signed_gate.v(5099)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66B080  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [31]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [31]),
    .c(\u_DIV_SIGNED/al_00000256AA899810 ),
    .o({open_n65,\u_DIV_SIGNED/al_00000256AA400D60 [31]}));  // al_ip/div_signed_gate.v(5183)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA66B190  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA422680 ),
    .en(div_signed_start),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA3DC030 ));  // al_ip/div_signed_gate.v(3215)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66B5D0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [21]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [21]),
    .c(\u_DIV_SIGNED/al_00000256AA89A260 ),
    .o({\u_DIV_SIGNED/al_00000256AA89ACB0 ,\u_DIV_SIGNED/al_00000256AA400D60 [21]}));  // al_ip/div_signed_gate.v(5106)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66B6E0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [4]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [4]),
    .c(\u_DIV_SIGNED/al_00000256AA8998C0 ),
    .o({\u_DIV_SIGNED/al_00000256AA89A470 ,\u_DIV_SIGNED/al_00000256AA400D60 [4]}));  // al_ip/div_signed_gate.v(5190)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66B7F0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [0]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [0]),
    .c(\u_DIV_SIGNED/al_00000256AA898580 ),
    .o({\u_DIV_SIGNED/al_00000256AA89A5D0 ,\u_DIV_SIGNED/al_00000256AA400D60 [0]}));  // al_ip/div_signed_gate.v(5008)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66BD40  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [10]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [10]),
    .c(\u_DIV_SIGNED/al_00000256AA899EF0 ),
    .o({\u_DIV_SIGNED/al_00000256AA899290 ,\u_DIV_SIGNED/al_00000256AA400D60 [10]}));  // al_ip/div_signed_gate.v(5022)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66C6D0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [11]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [11]),
    .c(\u_DIV_SIGNED/al_00000256AA899290 ),
    .o({\u_DIV_SIGNED/al_00000256AA899970 ,\u_DIV_SIGNED/al_00000256AA400D60 [11]}));  // al_ip/div_signed_gate.v(5029)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66C7E0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [24]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [24]),
    .c(\u_DIV_SIGNED/al_00000256AA899340 ),
    .o({\u_DIV_SIGNED/al_00000256AA898D10 ,\u_DIV_SIGNED/al_00000256AA400D60 [24]}));  // al_ip/div_signed_gate.v(5127)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66CB10  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [13]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [13]),
    .c(\u_DIV_SIGNED/al_00000256AA8996B0 ),
    .o({\u_DIV_SIGNED/al_00000256AA8993F0 ,\u_DIV_SIGNED/al_00000256AA400D60 [13]}));  // al_ip/div_signed_gate.v(5043)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66D170  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [1]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [1]),
    .c(\u_DIV_SIGNED/al_00000256AA89A5D0 ),
    .o({\u_DIV_SIGNED/al_00000256AA899760 ,\u_DIV_SIGNED/al_00000256AA400D60 [1]}));  // al_ip/div_signed_gate.v(5015)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA66D280  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [17]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [17]),
    .c(\u_DIV_SIGNED/al_00000256AA8988F0 ),
    .o({\u_DIV_SIGNED/al_00000256AA8994A0 ,\u_DIV_SIGNED/al_00000256AA400D60 [17]}));  // al_ip/div_signed_gate.v(5071)
  AL_DFF_0 \u_DIV_SIGNED/al_00000256AA66ED10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(i_mdu_op1[31]),
    .en(1'b1),
    .sr(~mdu_vld),
    .ss(1'b0),
    .q(\u_DIV_SIGNED/al_00000256AA3DC5B0 ));  // al_ip/div_signed_gate.v(4997)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6708B0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [5]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [5]),
    .c(\u_DIV_SIGNED/al_00000256AA89A470 ),
    .o({\u_DIV_SIGNED/al_00000256AA89A680 ,\u_DIV_SIGNED/al_00000256AA400D60 [5]}));  // al_ip/div_signed_gate.v(5197)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_DIV_SIGNED/al_00000256AA672670  (
    .a(1'b0),
    .b(1'b0),
    .c(1'b0),
    .o({\u_DIV_SIGNED/al_00000256AA6537E0 ,open_n66}));  // al_ip/div_signed_gate.v(1834)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_DIV_SIGNED/al_00000256AA672780  (
    .a(\u_DIV_SIGNED/al_00000256AA0CE7C0 [0]),
    .b(1'b1),
    .c(\u_DIV_SIGNED/al_00000256AA6537E0 ),
    .o({\u_DIV_SIGNED/al_00000256AA6547B0 ,\u_DIV_SIGNED/al_00000256AA0D29D0 [0]}));  // al_ip/div_signed_gate.v(1792)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_DIV_SIGNED/al_00000256AA672BC0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CE7C0 [1]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA6547B0 ),
    .o({\u_DIV_SIGNED/al_00000256AA653100 ,\u_DIV_SIGNED/al_00000256AA0D29D0 [1]}));  // al_ip/div_signed_gate.v(1799)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_DIV_SIGNED/al_00000256AA672DE0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CE7C0 [5]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA653E10 ),
    .o({open_n67,\u_DIV_SIGNED/al_00000256AA0D29D0 [5]}));  // al_ip/div_signed_gate.v(1827)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_DIV_SIGNED/al_00000256AA673880  (
    .a(\u_DIV_SIGNED/al_00000256AA0CE7C0 [4]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA6539F0 ),
    .o({\u_DIV_SIGNED/al_00000256AA653E10 ,\u_DIV_SIGNED/al_00000256AA0D29D0 [4]}));  // al_ip/div_signed_gate.v(1820)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_DIV_SIGNED/al_00000256AA675200  (
    .a(\u_DIV_SIGNED/al_00000256AA0CE7C0 [3]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA653890 ),
    .o({\u_DIV_SIGNED/al_00000256AA6539F0 ,\u_DIV_SIGNED/al_00000256AA0D29D0 [3]}));  // al_ip/div_signed_gate.v(1813)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u_DIV_SIGNED/al_00000256AA675530  (
    .a(1'b1),
    .b(1'b0),
    .c(1'b0),
    .o({\u_DIV_SIGNED/al_00000256AA88B690 ,open_n68}));  // al_ip/div_signed_gate.v(3205)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_DIV_SIGNED/al_00000256AA675750  (
    .a(\u_DIV_SIGNED/al_00000256AA0CE7C0 [2]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA653100 ),
    .o({\u_DIV_SIGNED/al_00000256AA653890 ,\u_DIV_SIGNED/al_00000256AA0D29D0 [2]}));  // al_ip/div_signed_gate.v(1806)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA675FD0  (
    .a(1'b0),
    .b(n34[12]),
    .c(\u_DIV_SIGNED/al_00000256AA421760 ),
    .o({\u_DIV_SIGNED/al_00000256AA422E10 ,\u_DIV_SIGNED/al_00000256AA0D5590 [12]}));  // al_ip/div_signed_gate.v(1867)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6760E0  (
    .a(1'b0),
    .b(n34[28]),
    .c(\u_DIV_SIGNED/al_00000256AA421290 ),
    .o({\u_DIV_SIGNED/al_00000256AA4216B0 ,\u_DIV_SIGNED/al_00000256AA0D5590 [28]}));  // al_ip/div_signed_gate.v(1986)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA676520  (
    .a(1'b0),
    .b(n34[7]),
    .c(\u_DIV_SIGNED/al_00000256AA422470 ),
    .o({\u_DIV_SIGNED/al_00000256AA4225D0 ,\u_DIV_SIGNED/al_00000256AA0D5590 [7]}));  // al_ip/div_signed_gate.v(2042)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA676A70  (
    .a(1'b0),
    .b(n34[10]),
    .c(\u_DIV_SIGNED/al_00000256AA423BD0 ),
    .o({\u_DIV_SIGNED/al_00000256AA423390 ,\u_DIV_SIGNED/al_00000256AA0D5590 [10]}));  // al_ip/div_signed_gate.v(1853)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA676B80  (
    .a(1'b0),
    .b(n34[20]),
    .c(\u_DIV_SIGNED/al_00000256AA421810 ),
    .o({\u_DIV_SIGNED/al_00000256AA421550 ,\u_DIV_SIGNED/al_00000256AA0D5590 [20]}));  // al_ip/div_signed_gate.v(1930)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA676C90  (
    .a(1'b0),
    .b(n34[22]),
    .c(\u_DIV_SIGNED/al_00000256AA4221B0 ),
    .o({\u_DIV_SIGNED/al_00000256AA423700 ,\u_DIV_SIGNED/al_00000256AA0D5590 [22]}));  // al_ip/div_signed_gate.v(1944)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA676DA0  (
    .a(1'b0),
    .b(n34[8]),
    .c(\u_DIV_SIGNED/al_00000256AA4225D0 ),
    .o({\u_DIV_SIGNED/al_00000256AA4232E0 ,\u_DIV_SIGNED/al_00000256AA0D5590 [8]}));  // al_ip/div_signed_gate.v(2049)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6771E0  (
    .a(1'b0),
    .b(n34[26]),
    .c(\u_DIV_SIGNED/al_00000256AA423230 ),
    .o({\u_DIV_SIGNED/al_00000256AA421CE0 ,\u_DIV_SIGNED/al_00000256AA0D5590 [26]}));  // al_ip/div_signed_gate.v(1972)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6772F0  (
    .a(1'b0),
    .b(n34[19]),
    .c(\u_DIV_SIGNED/al_00000256AA421130 ),
    .o({\u_DIV_SIGNED/al_00000256AA421810 ,\u_DIV_SIGNED/al_00000256AA0D5590 [19]}));  // al_ip/div_signed_gate.v(1916)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA677400  (
    .a(1'b0),
    .b(n34[16]),
    .c(\u_DIV_SIGNED/al_00000256AA4237B0 ),
    .o({\u_DIV_SIGNED/al_00000256AA421080 ,\u_DIV_SIGNED/al_00000256AA0D5590 [16]}));  // al_ip/div_signed_gate.v(1895)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA677510  (
    .a(1'b0),
    .b(n34[13]),
    .c(\u_DIV_SIGNED/al_00000256AA422E10 ),
    .o({\u_DIV_SIGNED/al_00000256AA423020 ,\u_DIV_SIGNED/al_00000256AA0D5590 [13]}));  // al_ip/div_signed_gate.v(1874)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA677620  (
    .a(1'b0),
    .b(n34[17]),
    .c(\u_DIV_SIGNED/al_00000256AA421080 ),
    .o({\u_DIV_SIGNED/al_00000256AA421EF0 ,\u_DIV_SIGNED/al_00000256AA0D5590 [17]}));  // al_ip/div_signed_gate.v(1902)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u_DIV_SIGNED/al_00000256AA677730  (
    .a(1'b0),
    .b(1'b0),
    .c(1'b0),
    .o({\u_DIV_SIGNED/al_00000256AA423910 ,open_n69}));  // al_ip/div_signed_gate.v(2063)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA677D90  (
    .a(1'b0),
    .b(n34[27]),
    .c(\u_DIV_SIGNED/al_00000256AA421CE0 ),
    .o({\u_DIV_SIGNED/al_00000256AA421290 ,\u_DIV_SIGNED/al_00000256AA0D5590 [27]}));  // al_ip/div_signed_gate.v(1979)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6782E0  (
    .a(1'b0),
    .b(n34[18]),
    .c(\u_DIV_SIGNED/al_00000256AA421EF0 ),
    .o({\u_DIV_SIGNED/al_00000256AA421130 ,\u_DIV_SIGNED/al_00000256AA0D5590 [18]}));  // al_ip/div_signed_gate.v(1909)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6783F0  (
    .a(1'b0),
    .b(n34[5]),
    .c(\u_DIV_SIGNED/al_00000256AA421C30 ),
    .o({\u_DIV_SIGNED/al_00000256AA4223C0 ,\u_DIV_SIGNED/al_00000256AA0D5590 [5]}));  // al_ip/div_signed_gate.v(2028)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA678500  (
    .a(1'b0),
    .b(n34[3]),
    .c(\u_DIV_SIGNED/al_00000256AA4218C0 ),
    .o({\u_DIV_SIGNED/al_00000256AA421B80 ,\u_DIV_SIGNED/al_00000256AA0D5590 [3]}));  // al_ip/div_signed_gate.v(2000)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA678610  (
    .a(1'b0),
    .b(n34[11]),
    .c(\u_DIV_SIGNED/al_00000256AA423390 ),
    .o({\u_DIV_SIGNED/al_00000256AA421760 ,\u_DIV_SIGNED/al_00000256AA0D5590 [11]}));  // al_ip/div_signed_gate.v(1860)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA678720  (
    .a(1'b0),
    .b(n34[21]),
    .c(\u_DIV_SIGNED/al_00000256AA421550 ),
    .o({\u_DIV_SIGNED/al_00000256AA4221B0 ,\u_DIV_SIGNED/al_00000256AA0D5590 [21]}));  // al_ip/div_signed_gate.v(1937)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA678A50  (
    .a(1'b0),
    .b(n34[14]),
    .c(\u_DIV_SIGNED/al_00000256AA423020 ),
    .o({\u_DIV_SIGNED/al_00000256AA422940 ,\u_DIV_SIGNED/al_00000256AA0D5590 [14]}));  // al_ip/div_signed_gate.v(1881)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA678B60  (
    .a(1'b0),
    .b(n34[1]),
    .c(\u_DIV_SIGNED/al_00000256AA423B20 ),
    .o({\u_DIV_SIGNED/al_00000256AA423650 ,\u_DIV_SIGNED/al_00000256AA0D5590 [1]}));  // al_ip/div_signed_gate.v(1846)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA678C70  (
    .a(1'b0),
    .b(n34[2]),
    .c(\u_DIV_SIGNED/al_00000256AA423650 ),
    .o({\u_DIV_SIGNED/al_00000256AA4218C0 ,\u_DIV_SIGNED/al_00000256AA0D5590 [2]}));  // al_ip/div_signed_gate.v(1923)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA678D80  (
    .a(1'b0),
    .b(n34[23]),
    .c(\u_DIV_SIGNED/al_00000256AA423700 ),
    .o({\u_DIV_SIGNED/al_00000256AA422520 ,\u_DIV_SIGNED/al_00000256AA0D5590 [23]}));  // al_ip/div_signed_gate.v(1951)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA678E90  (
    .a(1'b0),
    .b(n34[0]),
    .c(\u_DIV_SIGNED/al_00000256AA423910 ),
    .o({\u_DIV_SIGNED/al_00000256AA423B20 ,\u_DIV_SIGNED/al_00000256AA0D5590 [0]}));  // al_ip/div_signed_gate.v(1839)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA678FA0  (
    .a(1'b0),
    .b(n34[15]),
    .c(\u_DIV_SIGNED/al_00000256AA422940 ),
    .o({\u_DIV_SIGNED/al_00000256AA4237B0 ,\u_DIV_SIGNED/al_00000256AA0D5590 [15]}));  // al_ip/div_signed_gate.v(1888)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6790B0  (
    .a(1'b0),
    .b(n34[25]),
    .c(\u_DIV_SIGNED/al_00000256AA422310 ),
    .o({\u_DIV_SIGNED/al_00000256AA423230 ,\u_DIV_SIGNED/al_00000256AA0D5590 [25]}));  // al_ip/div_signed_gate.v(1965)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6791C0  (
    .a(1'b0),
    .b(n34[30]),
    .c(\u_DIV_SIGNED/al_00000256AA422EC0 ),
    .o({\u_DIV_SIGNED/al_00000256AA421600 ,\u_DIV_SIGNED/al_00000256AA0D5590 [30]}));  // al_ip/div_signed_gate.v(2007)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6792D0  (
    .a(1'b0),
    .b(n34[31]),
    .c(\u_DIV_SIGNED/al_00000256AA421600 ),
    .o({open_n70,\u_DIV_SIGNED/al_00000256AA0D5590 [31]}));  // al_ip/div_signed_gate.v(2014)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6793E0  (
    .a(1'b0),
    .b(n34[24]),
    .c(\u_DIV_SIGNED/al_00000256AA422520 ),
    .o({\u_DIV_SIGNED/al_00000256AA422310 ,\u_DIV_SIGNED/al_00000256AA0D5590 [24]}));  // al_ip/div_signed_gate.v(1958)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6794F0  (
    .a(1'b0),
    .b(n34[4]),
    .c(\u_DIV_SIGNED/al_00000256AA421B80 ),
    .o({\u_DIV_SIGNED/al_00000256AA421C30 ,\u_DIV_SIGNED/al_00000256AA0D5590 [4]}));  // al_ip/div_signed_gate.v(2021)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA679600  (
    .a(1'b0),
    .b(n34[9]),
    .c(\u_DIV_SIGNED/al_00000256AA4232E0 ),
    .o({\u_DIV_SIGNED/al_00000256AA423BD0 ,\u_DIV_SIGNED/al_00000256AA0D5590 [9]}));  // al_ip/div_signed_gate.v(2056)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA679710  (
    .a(1'b0),
    .b(n34[29]),
    .c(\u_DIV_SIGNED/al_00000256AA4216B0 ),
    .o({\u_DIV_SIGNED/al_00000256AA422EC0 ,\u_DIV_SIGNED/al_00000256AA0D5590 [29]}));  // al_ip/div_signed_gate.v(1993)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA679C60  (
    .a(1'b0),
    .b(n34[6]),
    .c(\u_DIV_SIGNED/al_00000256AA4223C0 ),
    .o({\u_DIV_SIGNED/al_00000256AA422470 ,\u_DIV_SIGNED/al_00000256AA0D5590 [6]}));  // al_ip/div_signed_gate.v(2035)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67A1B0  (
    .a(1'b0),
    .b(n35[2]),
    .c(\u_DIV_SIGNED/al_00000256AA3DD4D0 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DD840 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [2]}));  // al_ip/div_signed_gate.v(2152)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67B090  (
    .a(1'b0),
    .b(n35[18]),
    .c(\u_DIV_SIGNED/al_00000256AA3DD370 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DD420 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [18]}));  // al_ip/div_signed_gate.v(2138)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67B5E0  (
    .a(1'b0),
    .b(n35[16]),
    .c(\u_DIV_SIGNED/al_00000256AA3DCB30 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DDA50 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [16]}));  // al_ip/div_signed_gate.v(2124)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67B6F0  (
    .a(1'b0),
    .b(n35[5]),
    .c(\u_DIV_SIGNED/al_00000256AA3DB3D0 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DB060 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [5]}));  // al_ip/div_signed_gate.v(2257)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67B800  (
    .a(1'b0),
    .b(n35[21]),
    .c(\u_DIV_SIGNED/al_00000256AA3DCC90 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DC500 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [21]}));  // al_ip/div_signed_gate.v(2166)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67B910  (
    .a(1'b0),
    .b(n35[17]),
    .c(\u_DIV_SIGNED/al_00000256AA3DDA50 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DD370 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [17]}));  // al_ip/div_signed_gate.v(2131)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67BA20  (
    .a(1'b0),
    .b(n35[6]),
    .c(\u_DIV_SIGNED/al_00000256AA3DB060 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DB480 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [6]}));  // al_ip/div_signed_gate.v(2264)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67BB30  (
    .a(1'b0),
    .b(n35[25]),
    .c(\u_DIV_SIGNED/al_00000256AA3DD580 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DDBB0 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [25]}));  // al_ip/div_signed_gate.v(2194)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67BE60  (
    .a(1'b0),
    .b(n35[19]),
    .c(\u_DIV_SIGNED/al_00000256AA3DD420 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DBF80 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [19]}));  // al_ip/div_signed_gate.v(2145)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67C2A0  (
    .a(1'b0),
    .b(n35[23]),
    .c(\u_DIV_SIGNED/al_00000256AA3DB5E0 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DBCC0 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [23]}));  // al_ip/div_signed_gate.v(2180)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67C6E0  (
    .a(1'b0),
    .b(n35[28]),
    .c(\u_DIV_SIGNED/al_00000256AA3DCD40 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DC9D0 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [28]}));  // al_ip/div_signed_gate.v(2215)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67C7F0  (
    .a(1'b0),
    .b(n35[27]),
    .c(\u_DIV_SIGNED/al_00000256AA3DB320 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DCD40 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [27]}));  // al_ip/div_signed_gate.v(2208)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67C900  (
    .a(1'b0),
    .b(n35[11]),
    .c(\u_DIV_SIGNED/al_00000256AA3DB110 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DC3A0 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [11]}));  // al_ip/div_signed_gate.v(2089)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67CA10  (
    .a(1'b0),
    .b(n35[24]),
    .c(\u_DIV_SIGNED/al_00000256AA3DBCC0 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DD580 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [24]}));  // al_ip/div_signed_gate.v(2187)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67CB20  (
    .a(1'b0),
    .b(n35[7]),
    .c(\u_DIV_SIGNED/al_00000256AA3DB480 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DEB80 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [7]}));  // al_ip/div_signed_gate.v(2271)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67CC30  (
    .a(1'b0),
    .b(n35[22]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC500 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DB5E0 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [22]}));  // al_ip/div_signed_gate.v(2173)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u_DIV_SIGNED/al_00000256AA67CD40  (
    .a(1'b0),
    .b(1'b0),
    .c(1'b0),
    .o({\u_DIV_SIGNED/al_00000256AA3DD210 ,open_n71}));  // al_ip/div_signed_gate.v(2292)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67CE50  (
    .a(1'b0),
    .b(n35[0]),
    .c(\u_DIV_SIGNED/al_00000256AA3DD210 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DD2C0 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [0]}));  // al_ip/div_signed_gate.v(2068)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67D070  (
    .a(1'b0),
    .b(n35[12]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC3A0 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DC870 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [12]}));  // al_ip/div_signed_gate.v(2096)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67D180  (
    .a(1'b0),
    .b(n35[13]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC870 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DBC10 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [13]}));  // al_ip/div_signed_gate.v(2103)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67D290  (
    .a(1'b0),
    .b(n35[20]),
    .c(\u_DIV_SIGNED/al_00000256AA3DBF80 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DCC90 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [20]}));  // al_ip/div_signed_gate.v(2159)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67D4B0  (
    .a(1'b0),
    .b(n35[1]),
    .c(\u_DIV_SIGNED/al_00000256AA3DD2C0 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DD4D0 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [1]}));  // al_ip/div_signed_gate.v(2075)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67D5C0  (
    .a(1'b0),
    .b(n35[15]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC450 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DCB30 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [15]}));  // al_ip/div_signed_gate.v(2117)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67D6D0  (
    .a(1'b0),
    .b(n35[26]),
    .c(\u_DIV_SIGNED/al_00000256AA3DDBB0 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DB320 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [26]}));  // al_ip/div_signed_gate.v(2201)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67D7E0  (
    .a(1'b0),
    .b(n35[14]),
    .c(\u_DIV_SIGNED/al_00000256AA3DBC10 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DC450 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [14]}));  // al_ip/div_signed_gate.v(2110)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67D8F0  (
    .a(1'b0),
    .b(n35[30]),
    .c(\u_DIV_SIGNED/al_00000256AA3DD8F0 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DDB00 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [30]}));  // al_ip/div_signed_gate.v(2236)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67DA00  (
    .a(1'b0),
    .b(n35[31]),
    .c(\u_DIV_SIGNED/al_00000256AA3DDB00 ),
    .o({open_n72,\u_DIV_SIGNED/al_00000256AA3FF0F0 [31]}));  // al_ip/div_signed_gate.v(2243)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67DB10  (
    .a(1'b0),
    .b(n35[10]),
    .c(\u_DIV_SIGNED/al_00000256AA3DBD70 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DB110 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [10]}));  // al_ip/div_signed_gate.v(2082)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67DC20  (
    .a(1'b0),
    .b(n35[4]),
    .c(\u_DIV_SIGNED/al_00000256AA3DCA80 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DB3D0 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [4]}));  // al_ip/div_signed_gate.v(2250)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67DD30  (
    .a(1'b0),
    .b(n35[29]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC9D0 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DD8F0 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [29]}));  // al_ip/div_signed_gate.v(2222)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67DE40  (
    .a(1'b0),
    .b(n35[8]),
    .c(\u_DIV_SIGNED/al_00000256AA3DEB80 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DEA20 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [8]}));  // al_ip/div_signed_gate.v(2278)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67DF50  (
    .a(1'b0),
    .b(n35[9]),
    .c(\u_DIV_SIGNED/al_00000256AA3DEA20 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DBD70 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [9]}));  // al_ip/div_signed_gate.v(2285)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67E170  (
    .a(1'b0),
    .b(n35[3]),
    .c(\u_DIV_SIGNED/al_00000256AA3DD840 ),
    .o({\u_DIV_SIGNED/al_00000256AA3DCA80 ,\u_DIV_SIGNED/al_00000256AA3FF0F0 [3]}));  // al_ip/div_signed_gate.v(2229)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67E5B0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [8]),
    .c(\u_DIV_SIGNED/al_00000256AA444EC0 ),
    .o({\u_DIV_SIGNED/al_00000256AA3E0300 ,\u_DIV_SIGNED/al_00000256AA4072E0 [8]}));  // al_ip/div_signed_gate.v(2507)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67EC10  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [1]),
    .c(\u_DIV_SIGNED/al_00000256AA445230 ),
    .o({\u_DIV_SIGNED/al_00000256AA444050 ,\u_DIV_SIGNED/al_00000256AA4072E0 [1]}));  // al_ip/div_signed_gate.v(2304)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67ED20  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [14]),
    .c(\u_DIV_SIGNED/al_00000256AA445910 ),
    .o({\u_DIV_SIGNED/al_00000256AA443E40 ,\u_DIV_SIGNED/al_00000256AA4072E0 [14]}));  // al_ip/div_signed_gate.v(2339)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67EF40  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [21]),
    .c(\u_DIV_SIGNED/al_00000256AA444680 ),
    .o({\u_DIV_SIGNED/al_00000256AA4452E0 ,\u_DIV_SIGNED/al_00000256AA4072E0 [21]}));  // al_ip/div_signed_gate.v(2395)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67F050  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [19]),
    .c(\u_DIV_SIGNED/al_00000256AA443810 ),
    .o({\u_DIV_SIGNED/al_00000256AA4459C0 ,\u_DIV_SIGNED/al_00000256AA4072E0 [19]}));  // al_ip/div_signed_gate.v(2374)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67F160  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [23]),
    .c(\u_DIV_SIGNED/al_00000256AA444100 ),
    .o({\u_DIV_SIGNED/al_00000256AA445390 ,\u_DIV_SIGNED/al_00000256AA4072E0 [23]}));  // al_ip/div_signed_gate.v(2409)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67F270  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [16]),
    .c(\u_DIV_SIGNED/al_00000256AA443080 ),
    .o({\u_DIV_SIGNED/al_00000256AA443760 ,\u_DIV_SIGNED/al_00000256AA4072E0 [16]}));  // al_ip/div_signed_gate.v(2353)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67F5A0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [2]),
    .c(\u_DIV_SIGNED/al_00000256AA444050 ),
    .o({\u_DIV_SIGNED/al_00000256AA444CB0 ,\u_DIV_SIGNED/al_00000256AA4072E0 [2]}));  // al_ip/div_signed_gate.v(2381)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67F6B0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [20]),
    .c(\u_DIV_SIGNED/al_00000256AA4459C0 ),
    .o({\u_DIV_SIGNED/al_00000256AA444680 ,\u_DIV_SIGNED/al_00000256AA4072E0 [20]}));  // al_ip/div_signed_gate.v(2388)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67F8D0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [24]),
    .c(\u_DIV_SIGNED/al_00000256AA445390 ),
    .o({\u_DIV_SIGNED/al_00000256AA443130 ,\u_DIV_SIGNED/al_00000256AA4072E0 [24]}));  // al_ip/div_signed_gate.v(2416)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67F9E0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [22]),
    .c(\u_DIV_SIGNED/al_00000256AA4452E0 ),
    .o({\u_DIV_SIGNED/al_00000256AA444100 ,\u_DIV_SIGNED/al_00000256AA4072E0 [22]}));  // al_ip/div_signed_gate.v(2402)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67FAF0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [10]),
    .c(\u_DIV_SIGNED/al_00000256AA445860 ),
    .o({\u_DIV_SIGNED/al_00000256AA4436B0 ,\u_DIV_SIGNED/al_00000256AA4072E0 [10]}));  // al_ip/div_signed_gate.v(2311)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67FC00  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [15]),
    .c(\u_DIV_SIGNED/al_00000256AA443E40 ),
    .o({\u_DIV_SIGNED/al_00000256AA443080 ,\u_DIV_SIGNED/al_00000256AA4072E0 [15]}));  // al_ip/div_signed_gate.v(2346)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67FD10  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [13]),
    .c(\u_DIV_SIGNED/al_00000256AA443CE0 ),
    .o({\u_DIV_SIGNED/al_00000256AA445910 ,\u_DIV_SIGNED/al_00000256AA4072E0 [13]}));  // al_ip/div_signed_gate.v(2332)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67FE20  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [11]),
    .c(\u_DIV_SIGNED/al_00000256AA4436B0 ),
    .o({\u_DIV_SIGNED/al_00000256AA444520 ,\u_DIV_SIGNED/al_00000256AA4072E0 [11]}));  // al_ip/div_signed_gate.v(2318)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA67FF30  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [27]),
    .c(\u_DIV_SIGNED/al_00000256AA444B50 ),
    .o({\u_DIV_SIGNED/al_00000256AA445B20 ,\u_DIV_SIGNED/al_00000256AA4072E0 [27]}));  // al_ip/div_signed_gate.v(2437)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA680040  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [29]),
    .c(\u_DIV_SIGNED/al_00000256AA444260 ),
    .o({\u_DIV_SIGNED/al_00000256AA444310 ,\u_DIV_SIGNED/al_00000256AA4072E0 [29]}));  // al_ip/div_signed_gate.v(2451)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA680150  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [30]),
    .c(\u_DIV_SIGNED/al_00000256AA444310 ),
    .o({\u_DIV_SIGNED/al_00000256AA4445D0 ,\u_DIV_SIGNED/al_00000256AA4072E0 [30]}));  // al_ip/div_signed_gate.v(2465)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA680260  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [7]),
    .c(\u_DIV_SIGNED/al_00000256AA444E10 ),
    .o({\u_DIV_SIGNED/al_00000256AA444EC0 ,\u_DIV_SIGNED/al_00000256AA4072E0 [7]}));  // al_ip/div_signed_gate.v(2500)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6807B0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [0]),
    .c(\u_DIV_SIGNED/al_00000256AA443C30 ),
    .o({\u_DIV_SIGNED/al_00000256AA445230 ,\u_DIV_SIGNED/al_00000256AA4072E0 [0]}));  // al_ip/div_signed_gate.v(2297)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA680AE0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [6]),
    .c(\u_DIV_SIGNED/al_00000256AA444D60 ),
    .o({\u_DIV_SIGNED/al_00000256AA444E10 ,\u_DIV_SIGNED/al_00000256AA4072E0 [6]}));  // al_ip/div_signed_gate.v(2493)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA680E10  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [28]),
    .c(\u_DIV_SIGNED/al_00000256AA445B20 ),
    .o({\u_DIV_SIGNED/al_00000256AA444260 ,\u_DIV_SIGNED/al_00000256AA4072E0 [28]}));  // al_ip/div_signed_gate.v(2444)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA680F20  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [12]),
    .c(\u_DIV_SIGNED/al_00000256AA444520 ),
    .o({\u_DIV_SIGNED/al_00000256AA443CE0 ,\u_DIV_SIGNED/al_00000256AA4072E0 [12]}));  // al_ip/div_signed_gate.v(2325)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA681030  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [31]),
    .c(\u_DIV_SIGNED/al_00000256AA4445D0 ),
    .o({open_n73,\u_DIV_SIGNED/al_00000256AA4072E0 [31]}));  // al_ip/div_signed_gate.v(2472)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6817A0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [26]),
    .c(\u_DIV_SIGNED/al_00000256AA445020 ),
    .o({\u_DIV_SIGNED/al_00000256AA444B50 ,\u_DIV_SIGNED/al_00000256AA4072E0 [26]}));  // al_ip/div_signed_gate.v(2430)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6818B0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [17]),
    .c(\u_DIV_SIGNED/al_00000256AA443760 ),
    .o({\u_DIV_SIGNED/al_00000256AA443EF0 ,\u_DIV_SIGNED/al_00000256AA4072E0 [17]}));  // al_ip/div_signed_gate.v(2360)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6819C0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [4]),
    .c(\u_DIV_SIGNED/al_00000256AA444730 ),
    .o({\u_DIV_SIGNED/al_00000256AA444940 ,\u_DIV_SIGNED/al_00000256AA4072E0 [4]}));  // al_ip/div_signed_gate.v(2479)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA681CF0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [9]),
    .c(\u_DIV_SIGNED/al_00000256AA3E0300 ),
    .o({\u_DIV_SIGNED/al_00000256AA445860 ,\u_DIV_SIGNED/al_00000256AA4072E0 [9]}));  // al_ip/div_signed_gate.v(2514)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA682020  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [18]),
    .c(\u_DIV_SIGNED/al_00000256AA443EF0 ),
    .o({\u_DIV_SIGNED/al_00000256AA443810 ,\u_DIV_SIGNED/al_00000256AA4072E0 [18]}));  // al_ip/div_signed_gate.v(2367)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA682130  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [5]),
    .c(\u_DIV_SIGNED/al_00000256AA444940 ),
    .o({\u_DIV_SIGNED/al_00000256AA444D60 ,\u_DIV_SIGNED/al_00000256AA4072E0 [5]}));  // al_ip/div_signed_gate.v(2486)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u_DIV_SIGNED/al_00000256AA682240  (
    .a(1'b0),
    .b(1'b0),
    .c(1'b0),
    .o({\u_DIV_SIGNED/al_00000256AA443C30 ,open_n74}));  // al_ip/div_signed_gate.v(2521)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA682350  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [3]),
    .c(\u_DIV_SIGNED/al_00000256AA444CB0 ),
    .o({\u_DIV_SIGNED/al_00000256AA444730 ,\u_DIV_SIGNED/al_00000256AA4072E0 [3]}));  // al_ip/div_signed_gate.v(2458)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA682460  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [25]),
    .c(\u_DIV_SIGNED/al_00000256AA443130 ),
    .o({\u_DIV_SIGNED/al_00000256AA445020 ,\u_DIV_SIGNED/al_00000256AA4072E0 [25]}));  // al_ip/div_signed_gate.v(2423)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA6828A0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [4]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [4]),
    .c(\u_DIV_SIGNED/al_00000256AA88D000 ),
    .o({\u_DIV_SIGNED/al_00000256AA88ADA0 ,open_n75}));  // al_ip/div_signed_gate.v(3002)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA682AC0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [7]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [7]),
    .c(\u_DIV_SIGNED/al_00000256AA88D0B0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88AAE0 ,open_n76}));  // al_ip/div_signed_gate.v(3184)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA682BD0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [9]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [9]),
    .c(\u_DIV_SIGNED/al_00000256AA88A980 ),
    .o({\u_DIV_SIGNED/al_00000256AA88AA30 ,open_n77}));  // al_ip/div_signed_gate.v(3198)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA682CE0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [12]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [12]),
    .c(\u_DIV_SIGNED/al_00000256AA88D160 ),
    .o({\u_DIV_SIGNED/al_00000256AA88A8D0 ,open_n78}));  // al_ip/div_signed_gate.v(2792)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA682DF0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [13]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [13]),
    .c(\u_DIV_SIGNED/al_00000256AA88A8D0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88AFB0 ,open_n79}));  // al_ip/div_signed_gate.v(2799)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA682F00  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [17]),
    .c(\u_DIV_SIGNED/al_00000256AA88BED0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C2F0 ,\u_DIV_SIGNED/al_00000256AA40B170 [17]}));  // al_ip/div_signed_gate.v(2589)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA683010  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [16]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [16]),
    .c(\u_DIV_SIGNED/al_00000256AA88AB90 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B110 ,open_n80}));  // al_ip/div_signed_gate.v(2820)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA683120  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [17]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [17]),
    .c(\u_DIV_SIGNED/al_00000256AA88B110 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B3D0 ,open_n81}));  // al_ip/div_signed_gate.v(2827)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA683230  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [9]),
    .c(\u_DIV_SIGNED/al_00000256AA88AF00 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C920 ,\u_DIV_SIGNED/al_00000256AA40B170 [9]}));  // al_ip/div_signed_gate.v(2743)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA683340  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [18]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [18]),
    .c(\u_DIV_SIGNED/al_00000256AA88B3D0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B480 ,open_n82}));  // al_ip/div_signed_gate.v(2834)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA683450  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [6]),
    .c(\u_DIV_SIGNED/al_00000256AA88CC90 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B530 ,\u_DIV_SIGNED/al_00000256AA40B170 [6]}));  // al_ip/div_signed_gate.v(2722)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA683560  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [19]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [19]),
    .c(\u_DIV_SIGNED/al_00000256AA88B480 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B740 ,open_n83}));  // al_ip/div_signed_gate.v(2841)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA683670  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [7]),
    .c(\u_DIV_SIGNED/al_00000256AA88B530 ),
    .o({\u_DIV_SIGNED/al_00000256AA88CD40 ,\u_DIV_SIGNED/al_00000256AA40B170 [7]}));  // al_ip/div_signed_gate.v(2729)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA683780  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [13]),
    .c(\u_DIV_SIGNED/al_00000256AA88C240 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C9D0 ,\u_DIV_SIGNED/al_00000256AA40B170 [13]}));  // al_ip/div_signed_gate.v(2561)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA683890  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [2]),
    .c(\u_DIV_SIGNED/al_00000256AA88B1C0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88AC40 ,\u_DIV_SIGNED/al_00000256AA40B170 [2]}));  // al_ip/div_signed_gate.v(2610)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA6839A0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [8]),
    .c(\u_DIV_SIGNED/al_00000256AA88CD40 ),
    .o({\u_DIV_SIGNED/al_00000256AA88AF00 ,\u_DIV_SIGNED/al_00000256AA40B170 [8]}));  // al_ip/div_signed_gate.v(2736)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA683AB0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [18]),
    .c(\u_DIV_SIGNED/al_00000256AA88C2F0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88CEA0 ,\u_DIV_SIGNED/al_00000256AA40B170 [18]}));  // al_ip/div_signed_gate.v(2596)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA683BC0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [6]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [6]),
    .c(\u_DIV_SIGNED/al_00000256AA88AE50 ),
    .o({\u_DIV_SIGNED/al_00000256AA88D0B0 ,open_n84}));  // al_ip/div_signed_gate.v(3156)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA683CD0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [15]),
    .c(\u_DIV_SIGNED/al_00000256AA88C660 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B8A0 ,\u_DIV_SIGNED/al_00000256AA40B170 [15]}));  // al_ip/div_signed_gate.v(2575)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA683EF0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [21]),
    .c(\u_DIV_SIGNED/al_00000256AA88CBE0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B320 ,\u_DIV_SIGNED/al_00000256AA40B170 [21]}));  // al_ip/div_signed_gate.v(2624)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA684000  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [10]),
    .c(\u_DIV_SIGNED/al_00000256AA88C920 ),
    .o({\u_DIV_SIGNED/al_00000256AA88D420 ,\u_DIV_SIGNED/al_00000256AA40B170 [10]}));  // al_ip/div_signed_gate.v(2540)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA684110  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [26]),
    .c(\u_DIV_SIGNED/al_00000256AA88D2C0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B950 ,\u_DIV_SIGNED/al_00000256AA40B170 [26]}));  // al_ip/div_signed_gate.v(2659)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA684440  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [22]),
    .c(\u_DIV_SIGNED/al_00000256AA88B320 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C5B0 ,\u_DIV_SIGNED/al_00000256AA40B170 [22]}));  // al_ip/div_signed_gate.v(2631)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA684550  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [4]),
    .c(\u_DIV_SIGNED/al_00000256AA88ACF0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B270 ,\u_DIV_SIGNED/al_00000256AA40B170 [4]}));  // al_ip/div_signed_gate.v(2708)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u_DIV_SIGNED/al_00000256AA684660  (
    .a(1'b0),
    .b(1'b0),
    .c(1'b0),
    .o({\u_DIV_SIGNED/al_00000256AA88D210 ,open_n85}));  // al_ip/div_signed_gate.v(2750)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA684880  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [11]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [11]),
    .c(\u_DIV_SIGNED/al_00000256AA88BCC0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88D160 ,open_n86}));  // al_ip/div_signed_gate.v(2785)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA684990  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [14]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [14]),
    .c(\u_DIV_SIGNED/al_00000256AA88AFB0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C3A0 ,open_n87}));  // al_ip/div_signed_gate.v(2806)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA684AA0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [14]),
    .c(\u_DIV_SIGNED/al_00000256AA88C9D0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C660 ,\u_DIV_SIGNED/al_00000256AA40B170 [14]}));  // al_ip/div_signed_gate.v(2568)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA684BB0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [5]),
    .c(\u_DIV_SIGNED/al_00000256AA88B270 ),
    .o({\u_DIV_SIGNED/al_00000256AA88CC90 ,\u_DIV_SIGNED/al_00000256AA40B170 [5]}));  // al_ip/div_signed_gate.v(2715)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA684CC0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [15]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [15]),
    .c(\u_DIV_SIGNED/al_00000256AA88C3A0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88AB90 ,open_n88}));  // al_ip/div_signed_gate.v(2813)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA684DD0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [25]),
    .c(\u_DIV_SIGNED/al_00000256AA88CA80 ),
    .o({\u_DIV_SIGNED/al_00000256AA88D2C0 ,\u_DIV_SIGNED/al_00000256AA40B170 [25]}));  // al_ip/div_signed_gate.v(2652)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA684EE0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [19]),
    .c(\u_DIV_SIGNED/al_00000256AA88CEA0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B5E0 ,\u_DIV_SIGNED/al_00000256AA40B170 [19]}));  // al_ip/div_signed_gate.v(2603)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA685100  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [20]),
    .c(\u_DIV_SIGNED/al_00000256AA88B5E0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88CBE0 ,\u_DIV_SIGNED/al_00000256AA40B170 [20]}));  // al_ip/div_signed_gate.v(2617)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA685210  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [29]),
    .c(\u_DIV_SIGNED/al_00000256AA88B060 ),
    .o({\u_DIV_SIGNED/al_00000256AA88CB30 ,\u_DIV_SIGNED/al_00000256AA40B170 [29]}));  // al_ip/div_signed_gate.v(2680)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA685430  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [0]),
    .c(\u_DIV_SIGNED/al_00000256AA88D210 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C190 ,\u_DIV_SIGNED/al_00000256AA40B170 [0]}));  // al_ip/div_signed_gate.v(2526)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA685540  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [23]),
    .c(\u_DIV_SIGNED/al_00000256AA88C5B0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88D370 ,\u_DIV_SIGNED/al_00000256AA40B170 [23]}));  // al_ip/div_signed_gate.v(2638)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA685650  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [27]),
    .c(\u_DIV_SIGNED/al_00000256AA88B950 ),
    .o({\u_DIV_SIGNED/al_00000256AA88CF50 ,\u_DIV_SIGNED/al_00000256AA40B170 [27]}));  // al_ip/div_signed_gate.v(2666)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA685760  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [2]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [2]),
    .c(\u_DIV_SIGNED/al_00000256AA88CDF0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C450 ,open_n89}));  // al_ip/div_signed_gate.v(2848)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA685870  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [5]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [5]),
    .c(\u_DIV_SIGNED/al_00000256AA88ADA0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88AE50 ,open_n90}));  // al_ip/div_signed_gate.v(3079)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA685980  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [10]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [10]),
    .c(\u_DIV_SIGNED/al_00000256AA88AA30 ),
    .o({\u_DIV_SIGNED/al_00000256AA88BCC0 ,open_n91}));  // al_ip/div_signed_gate.v(2778)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA685A90  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [24]),
    .c(\u_DIV_SIGNED/al_00000256AA88D370 ),
    .o({\u_DIV_SIGNED/al_00000256AA88CA80 ,\u_DIV_SIGNED/al_00000256AA40B170 [24]}));  // al_ip/div_signed_gate.v(2645)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA685BA0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [16]),
    .c(\u_DIV_SIGNED/al_00000256AA88B8A0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88BED0 ,\u_DIV_SIGNED/al_00000256AA40B170 [16]}));  // al_ip/div_signed_gate.v(2582)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA685CB0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [3]),
    .c(\u_DIV_SIGNED/al_00000256AA88AC40 ),
    .o({\u_DIV_SIGNED/al_00000256AA88ACF0 ,\u_DIV_SIGNED/al_00000256AA40B170 [3]}));  // al_ip/div_signed_gate.v(2687)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA685ED0  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [30]),
    .c(\u_DIV_SIGNED/al_00000256AA88CB30 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C710 ,\u_DIV_SIGNED/al_00000256AA40B170 [30]}));  // al_ip/div_signed_gate.v(2694)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA686200  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [31]),
    .c(\u_DIV_SIGNED/al_00000256AA88C710 ),
    .o({open_n92,\u_DIV_SIGNED/al_00000256AA40B170 [31]}));  // al_ip/div_signed_gate.v(2701)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA686310  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [1]),
    .c(\u_DIV_SIGNED/al_00000256AA88C190 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B1C0 ,\u_DIV_SIGNED/al_00000256AA40B170 [1]}));  // al_ip/div_signed_gate.v(2533)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA686420  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [1]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [1]),
    .c(\u_DIV_SIGNED/al_00000256AA88C500 ),
    .o({\u_DIV_SIGNED/al_00000256AA88CDF0 ,open_n93}));  // al_ip/div_signed_gate.v(2771)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA686530  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [3]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [3]),
    .c(\u_DIV_SIGNED/al_00000256AA88C450 ),
    .o({\u_DIV_SIGNED/al_00000256AA88D000 ,open_n94}));  // al_ip/div_signed_gate.v(2925)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA686640  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [8]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [8]),
    .c(\u_DIV_SIGNED/al_00000256AA88AAE0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88A980 ,open_n95}));  // al_ip/div_signed_gate.v(3191)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA686860  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [12]),
    .c(\u_DIV_SIGNED/al_00000256AA88C870 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C240 ,\u_DIV_SIGNED/al_00000256AA40B170 [12]}));  // al_ip/div_signed_gate.v(2554)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA686970  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [11]),
    .c(\u_DIV_SIGNED/al_00000256AA88D420 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C870 ,\u_DIV_SIGNED/al_00000256AA40B170 [11]}));  // al_ip/div_signed_gate.v(2547)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA686A80  (
    .a(1'b0),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [28]),
    .c(\u_DIV_SIGNED/al_00000256AA88CF50 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B060 ,\u_DIV_SIGNED/al_00000256AA40B170 [28]}));  // al_ip/div_signed_gate.v(2673)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA686B90  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [0]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [0]),
    .c(\u_DIV_SIGNED/al_00000256AA88B690 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C500 ,open_n96}));  // al_ip/div_signed_gate.v(2764)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA686CA0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [56]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88FCB0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88F680 ,open_n97}));  // al_ip/div_signed_gate.v(3128)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA686DB0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [26]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [26]),
    .c(\u_DIV_SIGNED/al_00000256AA88BD70 ),
    .o({\u_DIV_SIGNED/al_00000256AA88BE20 ,open_n98}));  // al_ip/div_signed_gate.v(2897)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA686EC0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [58]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88E810 ),
    .o({\u_DIV_SIGNED/al_00000256AA88E340 ,open_n99}));  // al_ip/div_signed_gate.v(3142)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA686FD0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [61]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88F730 ),
    .o({\u_DIV_SIGNED/al_00000256AA88EA20 ,open_n100}));  // al_ip/div_signed_gate.v(3170)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA6870E0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [42]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88FAA0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88E130 ,open_n101}));  // al_ip/div_signed_gate.v(3023)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA6871F0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [62]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88EA20 ),
    .o({\u_DIV_SIGNED/al_00000256AA88D630 ,open_n102}));  // al_ip/div_signed_gate.v(3177)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA687300  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [38]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88E970 ),
    .o({\u_DIV_SIGNED/al_00000256AA88F3C0 ,open_n103}));  // al_ip/div_signed_gate.v(2988)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA687410  (
    .a(1'b0),
    .b(1'b1),
    .c(\u_DIV_SIGNED/al_00000256AA88D630 ),
    .o({open_n104,\u_DIV_SIGNED/al_00000256AA3DB7F0 }));  // al_ip/div_signed_gate.v(3210)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA687520  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [33]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88DB00 ),
    .o({\u_DIV_SIGNED/al_00000256AA88EC30 ,open_n105}));  // al_ip/div_signed_gate.v(2953)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA687630  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [6]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [6]),
    .c(\u_DIV_SIGNED/al_00000256AA89A680 ),
    .o({\u_DIV_SIGNED/al_00000256AA89AEC0 ,\u_DIV_SIGNED/al_00000256AA400D60 [6]}));  // al_ip/div_signed_gate.v(5204)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA687740  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [7]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [7]),
    .c(\u_DIV_SIGNED/al_00000256AA89AEC0 ),
    .o({\u_DIV_SIGNED/al_00000256AA89A730 ,\u_DIV_SIGNED/al_00000256AA400D60 [7]}));  // al_ip/div_signed_gate.v(5211)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA687850  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [57]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88F680 ),
    .o({\u_DIV_SIGNED/al_00000256AA88E810 ,open_n106}));  // al_ip/div_signed_gate.v(3135)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA687960  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [8]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [8]),
    .c(\u_DIV_SIGNED/al_00000256AA89A730 ),
    .o({\u_DIV_SIGNED/al_00000256AA899080 ,\u_DIV_SIGNED/al_00000256AA400D60 [8]}));  // al_ip/div_signed_gate.v(5218)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_SIGNED/al_00000256AA687A70  (
    .a(\u_DIV_SIGNED/al_00000256AA0CF470 [9]),
    .b(\u_DIV_SIGNED/al_00000256AA0D0BA0 [9]),
    .c(\u_DIV_SIGNED/al_00000256AA899080 ),
    .o({\u_DIV_SIGNED/al_00000256AA899EF0 ,\u_DIV_SIGNED/al_00000256AA400D60 [9]}));  // al_ip/div_signed_gate.v(5225)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA687B80  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [29]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [29]),
    .c(\u_DIV_SIGNED/al_00000256AA88C030 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C0E0 ,open_n107}));  // al_ip/div_signed_gate.v(2918)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA687C90  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [20]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [20]),
    .c(\u_DIV_SIGNED/al_00000256AA88B740 ),
    .o({\u_DIV_SIGNED/al_00000256AA88BA00 ,open_n108}));  // al_ip/div_signed_gate.v(2855)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA687DA0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [22]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [22]),
    .c(\u_DIV_SIGNED/al_00000256AA88B7F0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88BAB0 ,open_n109}));  // al_ip/div_signed_gate.v(2869)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA687EB0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [23]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [23]),
    .c(\u_DIV_SIGNED/al_00000256AA88BAB0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88BB60 ,open_n110}));  // al_ip/div_signed_gate.v(2876)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA687FC0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [27]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [27]),
    .c(\u_DIV_SIGNED/al_00000256AA88BE20 ),
    .o({\u_DIV_SIGNED/al_00000256AA88BF80 ,open_n111}));  // al_ip/div_signed_gate.v(2904)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA6880D0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [24]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [24]),
    .c(\u_DIV_SIGNED/al_00000256AA88BB60 ),
    .o({\u_DIV_SIGNED/al_00000256AA88BC10 ,open_n112}));  // al_ip/div_signed_gate.v(2883)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA6881E0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [34]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88EC30 ),
    .o({\u_DIV_SIGNED/al_00000256AA88EE40 ,open_n113}));  // al_ip/div_signed_gate.v(2960)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA6882F0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [28]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [28]),
    .c(\u_DIV_SIGNED/al_00000256AA88BF80 ),
    .o({\u_DIV_SIGNED/al_00000256AA88C030 ,open_n114}));  // al_ip/div_signed_gate.v(2911)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA688400  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [40]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88FD60 ),
    .o({\u_DIV_SIGNED/al_00000256AA88F890 ,open_n115}));  // al_ip/div_signed_gate.v(3009)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA688510  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [43]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88E130 ),
    .o({\u_DIV_SIGNED/al_00000256AA88F260 ,open_n116}));  // al_ip/div_signed_gate.v(3030)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA688620  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [31]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [31]),
    .c(\u_DIV_SIGNED/al_00000256AA88FC00 ),
    .o({\u_DIV_SIGNED/al_00000256AA88F5D0 ,open_n117}));  // al_ip/div_signed_gate.v(2939)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA688730  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [41]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88F890 ),
    .o({\u_DIV_SIGNED/al_00000256AA88FAA0 ,open_n118}));  // al_ip/div_signed_gate.v(3016)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA688840  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [46]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88FB50 ),
    .o({\u_DIV_SIGNED/al_00000256AA88E1E0 ,open_n119}));  // al_ip/div_signed_gate.v(3051)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA688950  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [47]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88E1E0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88F310 ,open_n120}));  // al_ip/div_signed_gate.v(3058)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA688A60  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [32]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88F5D0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88DB00 ,open_n121}));  // al_ip/div_signed_gate.v(2946)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA688B70  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [37]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88F470 ),
    .o({\u_DIV_SIGNED/al_00000256AA88E970 ,open_n122}));  // al_ip/div_signed_gate.v(2981)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA688C80  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [45]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88DE70 ),
    .o({\u_DIV_SIGNED/al_00000256AA88FB50 ,open_n123}));  // al_ip/div_signed_gate.v(3044)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA688D90  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [49]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88DF20 ),
    .o({\u_DIV_SIGNED/al_00000256AA88F940 ,open_n124}));  // al_ip/div_signed_gate.v(3072)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA688EA0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [50]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88F940 ),
    .o({\u_DIV_SIGNED/al_00000256AA88F520 ,open_n125}));  // al_ip/div_signed_gate.v(3086)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA688FB0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [44]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88F260 ),
    .o({\u_DIV_SIGNED/al_00000256AA88DE70 ,open_n126}));  // al_ip/div_signed_gate.v(3037)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA6890C0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [25]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [25]),
    .c(\u_DIV_SIGNED/al_00000256AA88BC10 ),
    .o({\u_DIV_SIGNED/al_00000256AA88BD70 ,open_n127}));  // al_ip/div_signed_gate.v(2890)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA6891D0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [48]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88F310 ),
    .o({\u_DIV_SIGNED/al_00000256AA88DF20 ,open_n128}));  // al_ip/div_signed_gate.v(3065)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA6892E0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [21]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [21]),
    .c(\u_DIV_SIGNED/al_00000256AA88BA00 ),
    .o({\u_DIV_SIGNED/al_00000256AA88B7F0 ,open_n129}));  // al_ip/div_signed_gate.v(2862)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA6893F0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [52]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88ECE0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88F9F0 ,open_n130}));  // al_ip/div_signed_gate.v(3100)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA689500  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [53]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88F9F0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88E290 ,open_n131}));  // al_ip/div_signed_gate.v(3107)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA689610  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [54]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88E290 ),
    .o({\u_DIV_SIGNED/al_00000256AA88DFD0 ,open_n132}));  // al_ip/div_signed_gate.v(3114)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA689720  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [36]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88DD10 ),
    .o({\u_DIV_SIGNED/al_00000256AA88F470 ,open_n133}));  // al_ip/div_signed_gate.v(2974)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA689830  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [59]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88E340 ),
    .o({\u_DIV_SIGNED/al_00000256AA88DA50 ,open_n134}));  // al_ip/div_signed_gate.v(3149)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA689940  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [30]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [30]),
    .c(\u_DIV_SIGNED/al_00000256AA88C0E0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88FC00 ,open_n135}));  // al_ip/div_signed_gate.v(2932)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA689A50  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [60]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88DA50 ),
    .o({\u_DIV_SIGNED/al_00000256AA88F730 ,open_n136}));  // al_ip/div_signed_gate.v(3163)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA689B60  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [55]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88DFD0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88FCB0 ,open_n137}));  // al_ip/div_signed_gate.v(3121)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA689C70  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [39]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88F3C0 ),
    .o({\u_DIV_SIGNED/al_00000256AA88FD60 ,open_n138}));  // al_ip/div_signed_gate.v(2995)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA689D80  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [51]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88F520 ),
    .o({\u_DIV_SIGNED/al_00000256AA88ECE0 ,open_n139}));  // al_ip/div_signed_gate.v(3093)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_SIGNED/al_00000256AA689E90  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [35]),
    .b(1'b0),
    .c(\u_DIV_SIGNED/al_00000256AA88EE40 ),
    .o({\u_DIV_SIGNED/al_00000256AA88DD10 ,open_n140}));  // al_ip/div_signed_gate.v(2967)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE91F6C0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [30]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [30]));  // al_ip/div_unsigned_gate.v(2099)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE91F7D0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [6]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [7]));  // al_ip/div_unsigned_gate.v(2432)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE91F8E0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [5]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [6]));  // al_ip/div_unsigned_gate.v(2423)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE91F9F0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [7]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [8]));  // al_ip/div_unsigned_gate.v(2441)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE91FB00  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [8]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [9]));  // al_ip/div_unsigned_gate.v(2450)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE91FC10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [20]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [21]));  // al_ip/div_unsigned_gate.v(2297)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE91FD20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [22]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [23]));  // al_ip/div_unsigned_gate.v(2315)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE91FF40  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [13]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [14]));  // al_ip/div_unsigned_gate.v(2225)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE920050  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [16]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [16]));  // al_ip/div_unsigned_gate.v(1955)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE920160  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [19]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [19]));  // al_ip/div_unsigned_gate.v(1982)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE920270  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [27]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [27]));  // al_ip/div_unsigned_gate.v(2063)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE920490  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [21]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [22]));  // al_ip/div_unsigned_gate.v(2306)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9205A0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [23]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [24]));  // al_ip/div_unsigned_gate.v(2324)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9206B0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [24]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [25]));  // al_ip/div_unsigned_gate.v(2333)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9207C0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [27]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [28]));  // al_ip/div_unsigned_gate.v(2360)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9208D0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [28]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [29]));  // al_ip/div_unsigned_gate.v(2369)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9209E0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [28]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [28]));  // al_ip/div_unsigned_gate.v(2072)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE920D10  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [1]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[1]));  // al_ip/div_unsigned_gate.v(2468)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE920E20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [3]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [4]));  // al_ip/div_unsigned_gate.v(2405)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE920F30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [26]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [26]));  // al_ip/div_unsigned_gate.v(2054)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE921040  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [14]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [15]));  // al_ip/div_unsigned_gate.v(2234)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE921150  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [29]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [30]));  // al_ip/div_unsigned_gate.v(2387)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE921260  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [0]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [1]));  // al_ip/div_unsigned_gate.v(2180)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE921370  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [26]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [27]));  // al_ip/div_unsigned_gate.v(2351)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE921480  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [30]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [31]));  // al_ip/div_unsigned_gate.v(2396)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE921590  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [15]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [15]));  // al_ip/div_unsigned_gate.v(1946)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9216A0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [12]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [13]));  // al_ip/div_unsigned_gate.v(2216)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9217B0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [15]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [16]));  // al_ip/div_unsigned_gate.v(2243)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9218C0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [19]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [20]));  // al_ip/div_unsigned_gate.v(2288)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE921AE0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [4]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[4]));  // al_ip/div_unsigned_gate.v(2693)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE921BF0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [5]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[5]));  // al_ip/div_unsigned_gate.v(2702)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE921D00  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [20]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [20]));  // al_ip/div_unsigned_gate.v(2000)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE921E10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [24]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [24]));  // al_ip/div_unsigned_gate.v(2036)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE921F20  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [10]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [11]));  // al_ip/div_unsigned_gate.v(2198)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE922030  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [17]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [17]));  // al_ip/div_unsigned_gate.v(1964)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE922140  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [2]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [3]));  // al_ip/div_unsigned_gate.v(2378)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE922250  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [4]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [5]));  // al_ip/div_unsigned_gate.v(2414)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE922360  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [1]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [2]));  // al_ip/div_unsigned_gate.v(2279)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE922470  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [11]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [12]));  // al_ip/div_unsigned_gate.v(2207)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9227A0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [0]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[0]));  // al_ip/div_unsigned_gate.v(2459)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9228B0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [25]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [25]));  // al_ip/div_unsigned_gate.v(2045)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9229C0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [6]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[6]));  // al_ip/div_unsigned_gate.v(2711)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE922AD0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [23]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [23]));  // al_ip/div_unsigned_gate.v(2027)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE922BE0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [3]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[3]));  // al_ip/div_unsigned_gate.v(2666)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE922CF0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [7]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[7]));  // al_ip/div_unsigned_gate.v(2720)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE922E00  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [21]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [21]));  // al_ip/div_unsigned_gate.v(2009)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE922F10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [16]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [17]));  // al_ip/div_unsigned_gate.v(2252)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE923020  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [17]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [18]));  // al_ip/div_unsigned_gate.v(2261)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE923130  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [31]));  // al_ip/div_unsigned_gate.v(2108)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE923240  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [0]));  // al_ip/div_unsigned_gate.v(2171)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE923350  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [25]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [26]));  // al_ip/div_unsigned_gate.v(2342)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE923460  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [29]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [29]));  // al_ip/div_unsigned_gate.v(2081)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE923570  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [2]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[2]));  // al_ip/div_unsigned_gate.v(2567)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE923680  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [22]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [22]));  // al_ip/div_unsigned_gate.v(2018)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE923790  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [9]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [10]));  // al_ip/div_unsigned_gate.v(2189)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9238A0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [18]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [19]));  // al_ip/div_unsigned_gate.v(2270)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9239B0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [18]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [18]));  // al_ip/div_unsigned_gate.v(1973)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE923AC0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [2]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[2]));  // al_ip/div_unsigned_gate.v(2855)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE923CE0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [12]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[12]));  // al_ip/div_unsigned_gate.v(2495)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE923DF0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [14]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[14]));  // al_ip/div_unsigned_gate.v(2513)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE923F00  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [16]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[16]));  // al_ip/div_unsigned_gate.v(2531)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE924230  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [28]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[28]));  // al_ip/div_unsigned_gate.v(2648)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE924450  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [0]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[0]));  // al_ip/div_unsigned_gate.v(2747)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE924560  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [7]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[7]));  // al_ip/div_unsigned_gate.v(3008)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE924890  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [13]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[13]));  // al_ip/div_unsigned_gate.v(2504)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE924DE0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [15]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[15]));  // al_ip/div_unsigned_gate.v(2522)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE925000  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [19]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[19]));  // al_ip/div_unsigned_gate.v(2558)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE925110  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [23]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[23]));  // al_ip/div_unsigned_gate.v(2603)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE925220  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [24]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[24]));  // al_ip/div_unsigned_gate.v(2612)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE925330  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [27]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[27]));  // al_ip/div_unsigned_gate.v(2639)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE925550  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [8]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[8]));  // al_ip/div_unsigned_gate.v(2729)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE925660  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [9]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[9]));  // al_ip/div_unsigned_gate.v(2738)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE925770  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [17]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[17]));  // al_ip/div_unsigned_gate.v(2540)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE925880  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [30]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[30]));  // al_ip/div_unsigned_gate.v(2675)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE925AA0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [31]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[31]));  // al_ip/div_unsigned_gate.v(2684)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE925BB0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [25]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[25]));  // al_ip/div_unsigned_gate.v(2621)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE925CC0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [22]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[22]));  // al_ip/div_unsigned_gate.v(2594)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE926430  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [26]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[26]));  // al_ip/div_unsigned_gate.v(2630)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE926540  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [18]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[18]));  // al_ip/div_unsigned_gate.v(2549)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE926650  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [20]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[20]));  // al_ip/div_unsigned_gate.v(2576)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE926870  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [3]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[3]));  // al_ip/div_unsigned_gate.v(2954)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE926980  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [4]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[4]));  // al_ip/div_unsigned_gate.v(2981)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE926A90  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [5]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[5]));  // al_ip/div_unsigned_gate.v(2990)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE926CB0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [6]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[6]));  // al_ip/div_unsigned_gate.v(2999)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE926ED0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [11]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[11]));  // al_ip/div_unsigned_gate.v(2486)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE926FE0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [21]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[21]));  // al_ip/div_unsigned_gate.v(2585)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE9270F0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [29]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[29]));  // al_ip/div_unsigned_gate.v(2657)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE927200  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [10]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_quo[10]));  // al_ip/div_unsigned_gate.v(2477)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DE927420  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [1]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[1]));  // al_ip/div_unsigned_gate.v(2756)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA92230  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [11]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[11]));  // al_ip/div_unsigned_gate.v(2774)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA92340  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [25]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[25]));  // al_ip/div_unsigned_gate.v(2909)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA92450  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E04A0 [4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [4]));  // al_ip/div_unsigned_gate.v(3071)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA92AB0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [9]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[9]));  // al_ip/div_unsigned_gate.v(3026)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA92BC0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [20]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[20]));  // al_ip/div_unsigned_gate.v(2864)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA93220  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [18]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[18]));  // al_ip/div_unsigned_gate.v(2837)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA93330  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [23]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[23]));  // al_ip/div_unsigned_gate.v(2891)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA93550  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [17]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[17]));  // al_ip/div_unsigned_gate.v(2828)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA93660  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [29]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[29]));  // al_ip/div_unsigned_gate.v(2945)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA93880  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [8]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[8]));  // al_ip/div_unsigned_gate.v(3017)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA93AA0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E04A0 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [2]));  // al_ip/div_unsigned_gate.v(3053)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA93DD0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [16]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[16]));  // al_ip/div_unsigned_gate.v(2819)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA94320  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [19]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[19]));  // al_ip/div_unsigned_gate.v(2846)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA94540  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [13]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[13]));  // al_ip/div_unsigned_gate.v(2792)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA94870  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [10]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[10]));  // al_ip/div_unsigned_gate.v(2765)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA94980  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [12]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[12]));  // al_ip/div_unsigned_gate.v(2783)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA94A90  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [15]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[15]));  // al_ip/div_unsigned_gate.v(2810)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA94CB0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [14]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[14]));  // al_ip/div_unsigned_gate.v(2801)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA94DC0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [21]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[21]));  // al_ip/div_unsigned_gate.v(2873)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA94ED0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [22]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[22]));  // al_ip/div_unsigned_gate.v(2882)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA94FE0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [26]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[26]));  // al_ip/div_unsigned_gate.v(2918)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA950F0  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [28]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[28]));  // al_ip/div_unsigned_gate.v(2936)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA95200  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [30]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[30]));  // al_ip/div_unsigned_gate.v(2963)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA95310  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E04A0 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [0]));  // al_ip/div_unsigned_gate.v(3035)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA95420  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E04A0 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [1]));  // al_ip/div_unsigned_gate.v(3044)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA95530  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E04A0 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [3]));  // al_ip/div_unsigned_gate.v(3062)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA95640  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E04A0 [5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [5]));  // al_ip/div_unsigned_gate.v(3080)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA95750  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [24]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[24]));  // al_ip/div_unsigned_gate.v(2900)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA95860  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [31]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[31]));  // al_ip/div_unsigned_gate.v(2972)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286DEA95970  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [27]),
    .en(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_rem[27]));  // al_ip/div_unsigned_gate.v(2927)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443B780  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [10]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [10]),
    .c(\u_DIV_UNSIGNED/al_00000286E4481BE0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4481B30 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [10]}));  // al_ip/div_unsigned_gate.v(3105)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443B9A0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [12]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [12]),
    .c(\u_DIV_UNSIGNED/al_00000286E4481030 ),
    .o({\u_DIV_UNSIGNED/al_00000286E44810E0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [12]}));  // al_ip/div_unsigned_gate.v(3119)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443BAB0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [14]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [14]),
    .c(\u_DIV_UNSIGNED/al_00000286E447F6C0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E44808A0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [14]}));  // al_ip/div_unsigned_gate.v(3133)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443BBC0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [15]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [15]),
    .c(\u_DIV_UNSIGNED/al_00000286E44808A0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E447FC40 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [15]}));  // al_ip/div_unsigned_gate.v(3140)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443BCD0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [18]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [18]),
    .c(\u_DIV_UNSIGNED/al_00000286E447FCF0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4480480 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [18]}));  // al_ip/div_unsigned_gate.v(3161)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443C000  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [1]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [1]),
    .c(\u_DIV_UNSIGNED/al_00000286E447F350 ),
    .o({\u_DIV_UNSIGNED/al_00000286E447FDA0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [1]}));  // al_ip/div_unsigned_gate.v(3098)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443C110  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [2]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [2]),
    .c(\u_DIV_UNSIGNED/al_00000286E447FDA0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E44805E0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [2]}));  // al_ip/div_unsigned_gate.v(3175)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443C220  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [0]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [0]),
    .c(\u_DIV_UNSIGNED/al_00000286E447F1F0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E447F350 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [0]}));  // al_ip/div_unsigned_gate.v(3091)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443C330  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [25]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [25]),
    .c(\u_DIV_UNSIGNED/al_00000286E447FF00 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4480110 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [25]}));  // al_ip/div_unsigned_gate.v(3217)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443C440  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [26]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [26]),
    .c(\u_DIV_UNSIGNED/al_00000286E4480110 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4480530 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [26]}));  // al_ip/div_unsigned_gate.v(3224)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443C550  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [27]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [27]),
    .c(\u_DIV_UNSIGNED/al_00000286E4480530 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4480270 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [27]}));  // al_ip/div_unsigned_gate.v(3231)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443C990  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [11]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [11]),
    .c(\u_DIV_UNSIGNED/al_00000286E4481B30 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4481030 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [11]}));  // al_ip/div_unsigned_gate.v(3112)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443CAA0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [16]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [16]),
    .c(\u_DIV_UNSIGNED/al_00000286E447FC40 ),
    .o({\u_DIV_UNSIGNED/al_00000286E44819D0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [16]}));  // al_ip/div_unsigned_gate.v(3147)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443CFF0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [17]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [17]),
    .c(\u_DIV_UNSIGNED/al_00000286E44819D0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E447FCF0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [17]}));  // al_ip/div_unsigned_gate.v(3154)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443D100  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [23]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [23]),
    .c(\u_DIV_UNSIGNED/al_00000286E4480CC0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4480A00 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [23]}));  // al_ip/div_unsigned_gate.v(3203)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443D210  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [28]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [28]),
    .c(\u_DIV_UNSIGNED/al_00000286E4480270 ),
    .o({\u_DIV_UNSIGNED/al_00000286E44812F0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [28]}));  // al_ip/div_unsigned_gate.v(3238)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443D320  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [19]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [19]),
    .c(\u_DIV_UNSIGNED/al_00000286E4480480 ),
    .o({\u_DIV_UNSIGNED/al_00000286E44803D0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [19]}));  // al_ip/div_unsigned_gate.v(3168)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443D430  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [29]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [29]),
    .c(\u_DIV_UNSIGNED/al_00000286E44812F0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4480AB0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [29]}));  // al_ip/div_unsigned_gate.v(3245)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443D540  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [3]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [3]),
    .c(\u_DIV_UNSIGNED/al_00000286E44805E0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4481500 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [3]}));  // al_ip/div_unsigned_gate.v(3252)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443DCB0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [20]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [20]),
    .c(\u_DIV_UNSIGNED/al_00000286E44803D0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E447FE50 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [20]}));  // al_ip/div_unsigned_gate.v(3182)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443DDC0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [21]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [21]),
    .c(\u_DIV_UNSIGNED/al_00000286E447FE50 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4481920 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [21]}));  // al_ip/div_unsigned_gate.v(3189)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443DED0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [24]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [24]),
    .c(\u_DIV_UNSIGNED/al_00000286E4480A00 ),
    .o({\u_DIV_UNSIGNED/al_00000286E447FF00 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [24]}));  // al_ip/div_unsigned_gate.v(3210)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443DFE0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [30]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [30]),
    .c(\u_DIV_UNSIGNED/al_00000286E4480AB0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4480B60 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [30]}));  // al_ip/div_unsigned_gate.v(3259)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443E0F0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [31]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [31]),
    .c(\u_DIV_UNSIGNED/al_00000286E4480B60 ),
    .o({open_n141,\u_DIV_UNSIGNED/al_00000286E57E1690 [31]}));  // al_ip/div_unsigned_gate.v(3266)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443E200  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [4]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [4]),
    .c(\u_DIV_UNSIGNED/al_00000286E4481500 ),
    .o({\u_DIV_UNSIGNED/al_00000286E44815B0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [4]}));  // al_ip/div_unsigned_gate.v(3273)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443E310  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [5]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [5]),
    .c(\u_DIV_UNSIGNED/al_00000286E44815B0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4481660 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [5]}));  // al_ip/div_unsigned_gate.v(3280)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443E530  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [6]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [6]),
    .c(\u_DIV_UNSIGNED/al_00000286E4481660 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4481710 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [6]}));  // al_ip/div_unsigned_gate.v(3287)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443E970  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [13]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [13]),
    .c(\u_DIV_UNSIGNED/al_00000286E44810E0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E447F6C0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [13]}));  // al_ip/div_unsigned_gate.v(3126)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E443EA80  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [22]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [22]),
    .c(\u_DIV_UNSIGNED/al_00000286E4481920 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4480CC0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [22]}));  // al_ip/div_unsigned_gate.v(3196)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E443ECA0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [8]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [8]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A262F0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A24820 ,open_n142}));  // al_ip/div_unsigned_gate.v(1292)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E443EDB0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [9]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [9]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A24820 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A24610 ,open_n143}));  // al_ip/div_unsigned_gate.v(1299)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E443EEC0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [12]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [12]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A248D0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A23F30 ,open_n144}));  // al_ip/div_unsigned_gate.v(893)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E443EFD0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [13]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [13]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A23F30 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A23E80 ,open_n145}));  // al_ip/div_unsigned_gate.v(900)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_DIV_UNSIGNED/al_00000286E443F300  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [0]),
    .b(1'b1),
    .c(\u_DIV_UNSIGNED/al_00000286E4A253D0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A24560 ,\u_DIV_UNSIGNED/al_00000286E57E03C0 [0]}));  // al_ip/div_unsigned_gate.v(809)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E443F630  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [14]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [14]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A23E80 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A23FE0 ,open_n146}));  // al_ip/div_unsigned_gate.v(907)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E443F850  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [15]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [15]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A23FE0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A24090 ,open_n147}));  // al_ip/div_unsigned_gate.v(914)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E443F960  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [17]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [17]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25060 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A263A0 ,open_n148}));  // al_ip/div_unsigned_gate.v(928)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E443FA70  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [18]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [18]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A263A0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A258A0 ,open_n149}));  // al_ip/div_unsigned_gate.v(935)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E443FB80  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [19]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [19]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A258A0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25110 ,open_n150}));  // al_ip/div_unsigned_gate.v(942)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_DIV_UNSIGNED/al_00000286E443FC90  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [4]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A257F0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A24A30 ,\u_DIV_UNSIGNED/al_00000286E57E03C0 [4]}));  // al_ip/div_unsigned_gate.v(837)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E443FDA0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [1]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [1]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25530 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A24AE0 ,open_n151}));  // al_ip/div_unsigned_gate.v(872)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E443FEB0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [21]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [21]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25950 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A251C0 ,open_n152}));  // al_ip/div_unsigned_gate.v(963)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E443FFC0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [22]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [22]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A251C0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25ED0 ,open_n153}));  // al_ip/div_unsigned_gate.v(970)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44400D0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [23]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [23]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25ED0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25270 ,open_n154}));  // al_ip/div_unsigned_gate.v(977)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44401E0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [24]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [24]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25270 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25A00 ,open_n155}));  // al_ip/div_unsigned_gate.v(984)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44402F0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [26]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [26]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25B60 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25C10 ,open_n156}));  // al_ip/div_unsigned_gate.v(998)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4440400  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [27]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [27]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25C10 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25CC0 ,open_n157}));  // al_ip/div_unsigned_gate.v(1005)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4440510  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [29]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [29]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25F80 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A26030 ,open_n158}));  // al_ip/div_unsigned_gate.v(1019)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4440620  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [30]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [30]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A26030 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A260E0 ,open_n159}));  // al_ip/div_unsigned_gate.v(1033)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4440730  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [31]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [31]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A260E0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A26870 ,open_n160}));  // al_ip/div_unsigned_gate.v(1040)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4440840  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [2]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [2]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A24AE0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A23D20 ,open_n161}));  // al_ip/div_unsigned_gate.v(949)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4440950  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [33]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A27BB0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A26920 ,open_n162}));  // al_ip/div_unsigned_gate.v(1054)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4440A60  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [34]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A26920 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A28810 ,open_n163}));  // al_ip/div_unsigned_gate.v(1061)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4440D90  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [28]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [28]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25CC0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25F80 ,open_n164}));  // al_ip/div_unsigned_gate.v(1012)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4440EA0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [35]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A28810 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A269D0 ,open_n165}));  // al_ip/div_unsigned_gate.v(1068)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4440FB0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [32]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A26870 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A27BB0 ,open_n166}));  // al_ip/div_unsigned_gate.v(1047)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44410C0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [36]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A269D0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A26A80 ,open_n167}));  // al_ip/div_unsigned_gate.v(1075)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD_CARRY"))
    \u_DIV_UNSIGNED/al_00000286E44411D0  (
    .a(1'b0),
    .b(1'b0),
    .c(1'b0),
    .o({\u_DIV_UNSIGNED/al_00000286E4A253D0 ,open_n168}));  // al_ip/div_unsigned_gate.v(851)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44412E0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [11]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [11]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25740 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A248D0 ,open_n169}));  // al_ip/div_unsigned_gate.v(886)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44413F0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [0]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [0]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A23DD0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25530 ,open_n170}));  // al_ip/div_unsigned_gate.v(865)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4441500  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [25]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [25]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25A00 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25B60 ,open_n171}));  // al_ip/div_unsigned_gate.v(991)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4441720  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [37]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A26A80 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A27420 ,open_n172}));  // al_ip/div_unsigned_gate.v(1082)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4441830  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [6]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [6]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A24770 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A24FB0 ,open_n173}));  // al_ip/div_unsigned_gate.v(1257)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4441A50  (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(div_unsigned_finish));  // al_ip/div_unsigned_gate.v(854)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_DIV_UNSIGNED/al_00000286E4441D80  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [1]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A24560 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A24DA0 ,\u_DIV_UNSIGNED/al_00000286E57E03C0 [1]}));  // al_ip/div_unsigned_gate.v(816)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_DIV_UNSIGNED/al_00000286E4441E90  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [2]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A24DA0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A24E50 ,\u_DIV_UNSIGNED/al_00000286E57E03C0 [2]}));  // al_ip/div_unsigned_gate.v(823)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_DIV_UNSIGNED/al_00000286E4441FA0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [5]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A24A30 ),
    .o({open_n174,\u_DIV_UNSIGNED/al_00000286E57E03C0 [5]}));  // al_ip/div_unsigned_gate.v(844)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44420B0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [10]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [10]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A24610 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25740 ,open_n175}));  // al_ip/div_unsigned_gate.v(879)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44422D0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [16]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [16]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A24090 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25060 ,open_n176}));  // al_ip/div_unsigned_gate.v(921)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44423E0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [20]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [20]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25110 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25950 ,open_n177}));  // al_ip/div_unsigned_gate.v(956)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44424F0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [7]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [7]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A24FB0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A262F0 ,open_n178}));  // al_ip/div_unsigned_gate.v(1285)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B_CARRY"))
    \u_DIV_UNSIGNED/al_00000286E4442600  (
    .a(1'b1),
    .b(1'b0),
    .c(1'b0),
    .o({\u_DIV_UNSIGNED/al_00000286E4A23DD0 ,open_n179}));  // al_ip/div_unsigned_gate.v(1306)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4442820  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [3]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [3]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A23D20 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25D70 ,open_n180}));  // al_ip/div_unsigned_gate.v(1026)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4442930  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [5]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [5]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25690 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A24770 ,open_n181}));  // al_ip/div_unsigned_gate.v(1180)
  AL_MAP_ADDER #(
    .ALUTYPE("ADD"))
    \u_DIV_UNSIGNED/al_00000286E4442D70  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [3]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A24E50 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A257F0 ,\u_DIV_UNSIGNED/al_00000286E57E03C0 [3]}));  // al_ip/div_unsigned_gate.v(830)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4442F90  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [4]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [4]),
    .c(\u_DIV_UNSIGNED/al_00000286E4A25D70 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A25690 ,open_n182}));  // al_ip/div_unsigned_gate.v(1103)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44432C0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [58]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A28080 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A28E40 ,open_n183}));  // al_ip/div_unsigned_gate.v(1243)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44433D0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [46]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A27790 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A27370 ,open_n184}));  // al_ip/div_unsigned_gate.v(1152)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44434E0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [49]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A27210 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A284A0 ,open_n185}));  // al_ip/div_unsigned_gate.v(1173)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44435F0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [52]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A26B30 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A26BE0 ,open_n186}));  // al_ip/div_unsigned_gate.v(1201)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4443700  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [45]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A27C60 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A27790 ,open_n187}));  // al_ip/div_unsigned_gate.v(1145)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4443810  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [61]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A27160 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A28290 ,open_n188}));  // al_ip/div_unsigned_gate.v(1271)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4443A30  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [38]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A27420 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A26F50 ,open_n189}));  // al_ip/div_unsigned_gate.v(1089)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4443B40  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [55]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A27B00 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A26C90 ,open_n190}));  // al_ip/div_unsigned_gate.v(1222)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4443C50  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [40]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A28AD0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A276E0 ,open_n191}));  // al_ip/div_unsigned_gate.v(1110)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44443C0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [44]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A28C30 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A27C60 ,open_n192}));  // al_ip/div_unsigned_gate.v(1138)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44444D0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [53]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A26BE0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A28D90 ,open_n193}));  // al_ip/div_unsigned_gate.v(1208)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44445E0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [60]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A27FD0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A27160 ,open_n194}));  // al_ip/div_unsigned_gate.v(1264)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB_CARRY"))
    \u_DIV_UNSIGNED/al_00000286E44446F0  (
    .a(1'b0),
    .b(1'b0),
    .c(1'b0),
    .o({\u_DIV_UNSIGNED/al_00000286E447F1F0 ,open_n195}));  // al_ip/div_unsigned_gate.v(3315)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4444800  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [41]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A276E0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A283F0 ,open_n196}));  // al_ip/div_unsigned_gate.v(1117)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4444910  (
    .a(1'b0),
    .b(1'b1),
    .c(\u_DIV_UNSIGNED/al_00000286E4A26D40 ),
    .o({open_n197,\u_DIV_UNSIGNED/al_00000286E5A5D8C0 }));  // al_ip/div_unsigned_gate.v(1311)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E4444F70  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [9]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [9]),
    .c(\u_DIV_UNSIGNED/al_00000286E44833F0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4481BE0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [9]}));  // al_ip/div_unsigned_gate.v(3308)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44453B0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [47]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A27370 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A28CE0 ,open_n198}));  // al_ip/div_unsigned_gate.v(1159)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44454C0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [42]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A283F0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A270B0 ,open_n199}));  // al_ip/div_unsigned_gate.v(1124)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44455D0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [59]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A28E40 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A27FD0 ,open_n200}));  // al_ip/div_unsigned_gate.v(1250)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44457F0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [39]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A26F50 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A28AD0 ,open_n201}));  // al_ip/div_unsigned_gate.v(1096)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4445F60  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [43]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A270B0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A28C30 ,open_n202}));  // al_ip/div_unsigned_gate.v(1131)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4446070  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [51]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A28B80 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A26B30 ,open_n203}));  // al_ip/div_unsigned_gate.v(1194)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4446180  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [57]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A272C0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A28080 ,open_n204}));  // al_ip/div_unsigned_gate.v(1236)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E44464B0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [48]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A28CE0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A27210 ,open_n205}));  // al_ip/div_unsigned_gate.v(1166)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4446C20  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [50]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A284A0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A28B80 ,open_n206}));  // al_ip/div_unsigned_gate.v(1187)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4446E40  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [62]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A28290 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A26D40 ,open_n207}));  // al_ip/div_unsigned_gate.v(1278)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4447060  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [54]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A28D90 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A27B00 ,open_n208}));  // al_ip/div_unsigned_gate.v(1215)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E4447170  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [7]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [7]),
    .c(\u_DIV_UNSIGNED/al_00000286E4481710 ),
    .o({\u_DIV_UNSIGNED/al_00000286E44817C0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [7]}));  // al_ip/div_unsigned_gate.v(3294)
  AL_MAP_ADDER #(
    .ALUTYPE("SUB"))
    \u_DIV_UNSIGNED/al_00000286E4447280  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [8]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [8]),
    .c(\u_DIV_UNSIGNED/al_00000286E44817C0 ),
    .o({\u_DIV_UNSIGNED/al_00000286E44833F0 ,\u_DIV_UNSIGNED/al_00000286E57E1690 [8]}));  // al_ip/div_unsigned_gate.v(3301)
  AL_MAP_ADDER #(
    .ALUTYPE("A_LE_B"))
    \u_DIV_UNSIGNED/al_00000286E4447390  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [56]),
    .b(1'b0),
    .c(\u_DIV_UNSIGNED/al_00000286E4A26C90 ),
    .o({\u_DIV_UNSIGNED/al_00000286E4A272C0 ,open_n209}));  // al_ip/div_unsigned_gate.v(1229)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC86D0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [55]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [55]));  // al_ip/div_unsigned_gate.v(1775)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC87E0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [5]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [5]));  // al_ip/div_unsigned_gate.v(2126)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC8B10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [57]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [57]));  // al_ip/div_unsigned_gate.v(1793)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC8D30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [3]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [3]));  // al_ip/div_unsigned_gate.v(2090)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC8E40  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [7]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [7]));  // al_ip/div_unsigned_gate.v(2144)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC8F50  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [8]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [8]));  // al_ip/div_unsigned_gate.v(2153)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC94A0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [4]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [4]));  // al_ip/div_unsigned_gate.v(2117)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC95B0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [2]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [2]));  // al_ip/div_unsigned_gate.v(1991)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC96C0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [6]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [6]));  // al_ip/div_unsigned_gate.v(2135)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC97D0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [9]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [9]));  // al_ip/div_unsigned_gate.v(2162)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC99F0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [56]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [56]));  // al_ip/div_unsigned_gate.v(1784)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC9B00  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [10]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [10]));  // al_ip/div_unsigned_gate.v(1901)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC9E30  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [11]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [11]));  // al_ip/div_unsigned_gate.v(1910)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BC9F40  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [12]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [12]));  // al_ip/div_unsigned_gate.v(1919)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BCA050  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [13]));  // al_ip/div_unsigned_gate.v(1928)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BCA270  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [14]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [14]));  // al_ip/div_unsigned_gate.v(1937)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BCB7B0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [58]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [58]));  // al_ip/div_unsigned_gate.v(1802)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BCB8C0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [59]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [59]));  // al_ip/div_unsigned_gate.v(1811)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BCB9D0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [60]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [60]));  // al_ip/div_unsigned_gate.v(1829)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BCBAE0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [61]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [61]));  // al_ip/div_unsigned_gate.v(1838)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BCBBF0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(n34[31]),
    .en(1'b1),
    .sr(~div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [62]));  // al_ip/div_unsigned_gate.v(1847)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BCBD00  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [0]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [0]));  // al_ip/div_unsigned_gate.v(1883)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BCC580  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [1]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [1]));  // al_ip/div_unsigned_gate.v(1892)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDD8B0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [47]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [47]));  // al_ip/div_unsigned_gate.v(1694)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDD9C0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [20]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [19]));  // al_ip/div_unsigned_gate.v(1415)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDDAD0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [52]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [52]));  // al_ip/div_unsigned_gate.v(1748)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDDBE0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [53]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [53]));  // al_ip/div_unsigned_gate.v(1757)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDDE00  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [54]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [54]));  // al_ip/div_unsigned_gate.v(1766)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDDF10  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [28]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [27]));  // al_ip/div_unsigned_gate.v(1496)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDE020  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [38]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [38]));  // al_ip/div_unsigned_gate.v(1604)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDE130  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [9]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [8]));  // al_ip/div_unsigned_gate.v(1865)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDE460  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [12]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [11]));  // al_ip/div_unsigned_gate.v(1343)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDE570  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [21]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [20]));  // al_ip/div_unsigned_gate.v(1433)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDE790  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [48]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [48]));  // al_ip/div_unsigned_gate.v(1703)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDE8A0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [2]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [1]));  // al_ip/div_unsigned_gate.v(1325)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDE9B0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [4]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [3]));  // al_ip/div_unsigned_gate.v(1523)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDEAC0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [7]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [6]));  // al_ip/div_unsigned_gate.v(1820)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDEBD0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [8]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [7]));  // al_ip/div_unsigned_gate.v(1856)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDECE0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [11]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [10]));  // al_ip/div_unsigned_gate.v(1334)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDEDF0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [35]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [35]));  // al_ip/div_unsigned_gate.v(1577)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDEF00  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [27]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [26]));  // al_ip/div_unsigned_gate.v(1487)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDF010  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [34]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [34]));  // al_ip/div_unsigned_gate.v(1568)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDF120  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [32]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [32]));  // al_ip/div_unsigned_gate.v(1550)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDF230  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [39]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [39]));  // al_ip/div_unsigned_gate.v(1613)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDF340  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [24]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [23]));  // al_ip/div_unsigned_gate.v(1460)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDF450  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [45]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [45]));  // al_ip/div_unsigned_gate.v(1676)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDF560  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [49]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [49]));  // al_ip/div_unsigned_gate.v(1712)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDF670  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [36]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [36]));  // al_ip/div_unsigned_gate.v(1586)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDF780  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [50]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [50]));  // al_ip/div_unsigned_gate.v(1730)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDF890  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [51]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [51]));  // al_ip/div_unsigned_gate.v(1739)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDF9A0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [22]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [21]));  // al_ip/div_unsigned_gate.v(1442)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDFAB0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [17]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [16]));  // al_ip/div_unsigned_gate.v(1388)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDFCD0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [1]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [0]));  // al_ip/div_unsigned_gate.v(1316)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDFDE0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [6]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [5]));  // al_ip/div_unsigned_gate.v(1721)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BDFEF0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [5]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [4]));  // al_ip/div_unsigned_gate.v(1622)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0110  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [30]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [29]));  // al_ip/div_unsigned_gate.v(1514)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0220  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [25]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [24]));  // al_ip/div_unsigned_gate.v(1469)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0330  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [15]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [14]));  // al_ip/div_unsigned_gate.v(1370)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0440  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [26]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [25]));  // al_ip/div_unsigned_gate.v(1478)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0550  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [31]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [30]));  // al_ip/div_unsigned_gate.v(1532)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0660  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [37]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [37]));  // al_ip/div_unsigned_gate.v(1595)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0770  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [3]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [2]));  // al_ip/div_unsigned_gate.v(1424)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0990  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [14]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [13]));  // al_ip/div_unsigned_gate.v(1361)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0AA0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [29]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [28]));  // al_ip/div_unsigned_gate.v(1505)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0BB0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [10]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [9]));  // al_ip/div_unsigned_gate.v(1874)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0CC0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [33]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [33]));  // al_ip/div_unsigned_gate.v(1559)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0DD0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [40]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [40]));  // al_ip/div_unsigned_gate.v(1631)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0EE0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [42]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [42]));  // al_ip/div_unsigned_gate.v(1649)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE0FF0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [19]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [18]));  // al_ip/div_unsigned_gate.v(1406)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE1100  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [43]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [43]));  // al_ip/div_unsigned_gate.v(1658)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE1210  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [23]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [22]));  // al_ip/div_unsigned_gate.v(1451)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE1320  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [44]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [44]));  // al_ip/div_unsigned_gate.v(1667)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE1430  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [46]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [46]));  // al_ip/div_unsigned_gate.v(1685)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE1540  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [16]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [15]));  // al_ip/div_unsigned_gate.v(1379)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE1650  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [41]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [41]));  // al_ip/div_unsigned_gate.v(1640)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE1760  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [13]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [12]));  // al_ip/div_unsigned_gate.v(1352)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE1A90  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [18]),
    .en(1'b1),
    .sr(div_unsigned_start),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [17]));  // al_ip/div_unsigned_gate.v(1397)
  AL_DFF_0 \u_DIV_UNSIGNED/al_00000286E4BE1BA0  (
    .ar(1'b0),
    .as(1'b0),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [31]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [31]));  // al_ip/div_unsigned_gate.v(1541)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E578F490  (
    .a(n35[16]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [16]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [16]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [16]));  // al_ip/div_unsigned_gate.v(441)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E578F5A0  (
    .a(n35[19]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [19]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [19]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [19]));  // al_ip/div_unsigned_gate.v(479)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E578F6B0  (
    .a(n35[2]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [2]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [2]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [2]));  // al_ip/div_unsigned_gate.v(489)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E578F7C0  (
    .a(n34[6]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [38]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [37]));  // al_ip/div_unsigned_gate.v(667)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E578F8D0  (
    .a(n34[18]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [50]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [49]));  // al_ip/div_unsigned_gate.v(241)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E578F9E0  (
    .a(n35[21]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [21]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [21]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [21]));  // al_ip/div_unsigned_gate.v(509)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E578FAF0  (
    .a(n34[9]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [41]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [40]));  // al_ip/div_unsigned_gate.v(802)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E578FC00  (
    .a(n34[10]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [42]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [41]));  // al_ip/div_unsigned_gate.v(177)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E578FD10  (
    .a(n34[22]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [54]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [53]));  // al_ip/div_unsigned_gate.v(281)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E578FE20  (
    .a(n35[3]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [3]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [3]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [3]));  // al_ip/div_unsigned_gate.v(607)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E578FF30  (
    .a(n35[4]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [4]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [4]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [4]));  // al_ip/div_unsigned_gate.v(637)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5790040  (
    .a(n34[14]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [46]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [45]));  // al_ip/div_unsigned_gate.v(209)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5790150  (
    .a(n35[5]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [5]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [5]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [5]));  // al_ip/div_unsigned_gate.v(647)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5790260  (
    .a(n35[20]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [20]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [20]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [20]));  // al_ip/div_unsigned_gate.v(499)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5790370  (
    .a(n34[16]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [48]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [47]));  // al_ip/div_unsigned_gate.v(225)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5790480  (
    .a(n34[20]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [52]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [51]));  // al_ip/div_unsigned_gate.v(265)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5790590  (
    .a(n34[24]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [56]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [55]));  // al_ip/div_unsigned_gate.v(297)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E57906A0  (
    .a(n34[29]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [61]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [60]));  // al_ip/div_unsigned_gate.v(337)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E57907B0  (
    .a(n34[30]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [62]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [61]));  // al_ip/div_unsigned_gate.v(353)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E57908C0  (
    .a(n34[7]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [39]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [38]));  // al_ip/div_unsigned_gate.v(768)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E57909D0  (
    .a(n35[11]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [11]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [11]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [11]));  // al_ip/div_unsigned_gate.v(391)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5790AE0  (
    .a(n34[21]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [53]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [52]));  // al_ip/div_unsigned_gate.v(273)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5790BF0  (
    .a(n35[17]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [17]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [17]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [17]));  // al_ip/div_unsigned_gate.v(459)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5790D00  (
    .a(n35[26]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [26]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [26]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [26]));  // al_ip/div_unsigned_gate.v(567)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5790E10  (
    .a(n34[15]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [47]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [46]));  // al_ip/div_unsigned_gate.v(217)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5790F20  (
    .a(n35[28]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [28]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [28]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [28]));  // al_ip/div_unsigned_gate.v(587)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791030  (
    .a(n35[7]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [7]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [7]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [7]));  // al_ip/div_unsigned_gate.v(675)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5791140  (
    .a(n34[3]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [35]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [34]));  // al_ip/div_unsigned_gate.v(345)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5791250  (
    .a(n34[2]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [34]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [33]));  // al_ip/div_unsigned_gate.v(257)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791360  (
    .a(n35[1]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [1]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [1]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [1]));  // al_ip/div_unsigned_gate.v(371)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5791470  (
    .a(n34[4]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [36]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [35]));  // al_ip/div_unsigned_gate.v(451)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5791580  (
    .a(n34[17]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [49]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [48]));  // al_ip/div_unsigned_gate.v(233)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791690  (
    .a(n35[22]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [22]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [22]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [22]));  // al_ip/div_unsigned_gate.v(519)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E57917A0  (
    .a(n35[23]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [23]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [23]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [23]));  // al_ip/div_unsigned_gate.v(529)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E57918B0  (
    .a(n34[5]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [37]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [36]));  // al_ip/div_unsigned_gate.v(559)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E57919C0  (
    .a(n35[24]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [24]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [24]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [24]));  // al_ip/div_unsigned_gate.v(539)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791AD0  (
    .a(n35[30]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [30]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [30]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [30]));  // al_ip/div_unsigned_gate.v(617)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791BE0  (
    .a(n35[10]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [10]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [10]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [10]));  // al_ip/div_unsigned_gate.v(381)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791CF0  (
    .a(n35[31]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [31]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [31]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [31]));  // al_ip/div_unsigned_gate.v(627)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791E00  (
    .a(n35[8]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [8]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [8]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [8]));  // al_ip/div_unsigned_gate.v(685)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791F10  (
    .a(n35[18]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [18]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [18]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [18]));  // al_ip/div_unsigned_gate.v(469)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792020  (
    .a(n34[26]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [58]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [57]));  // al_ip/div_unsigned_gate.v(313)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792130  (
    .a(n34[27]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [59]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [58]));  // al_ip/div_unsigned_gate.v(321)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792240  (
    .a(n34[12]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [44]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [43]));  // al_ip/div_unsigned_gate.v(193)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792350  (
    .a(n34[25]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [57]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [56]));  // al_ip/div_unsigned_gate.v(305)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5792460  (
    .a(n35[14]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [14]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [14]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [14]));  // al_ip/div_unsigned_gate.v(421)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5792570  (
    .a(n35[25]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [25]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [25]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [25]));  // al_ip/div_unsigned_gate.v(549)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5792680  (
    .a(n35[27]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [27]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [27]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [27]));  // al_ip/div_unsigned_gate.v(577)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5792790  (
    .a(n35[9]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [9]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [9]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [9]));  // al_ip/div_unsigned_gate.v(695)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E57928A0  (
    .a(n35[6]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [6]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [6]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [6]));  // al_ip/div_unsigned_gate.v(657)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E57929B0  (
    .a(n34[0]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [32]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [31]));  // al_ip/div_unsigned_gate.v(161)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5792AC0  (
    .a(n35[0]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [0]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [0]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [0]));  // al_ip/div_unsigned_gate.v(361)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5792BD0  (
    .a(n35[13]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [13]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [13]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [13]));  // al_ip/div_unsigned_gate.v(411)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792CE0  (
    .a(n34[13]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [45]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [44]));  // al_ip/div_unsigned_gate.v(201)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792DF0  (
    .a(n34[28]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [60]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [59]));  // al_ip/div_unsigned_gate.v(329)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792F00  (
    .a(n34[19]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [51]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [50]));  // al_ip/div_unsigned_gate.v(249)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5793010  (
    .a(n34[23]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [55]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [54]));  // al_ip/div_unsigned_gate.v(289)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5793120  (
    .a(n35[15]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [15]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [15]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [15]));  // al_ip/div_unsigned_gate.v(431)
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'b0001))
    \u_DIV_UNSIGNED/al_00000286E5793230  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [1]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [2]),
    .o(\u_DIV_UNSIGNED/al_00000286E4688A90 ));  // al_ip/div_unsigned_gate.v(705)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5793340  (
    .a(n35[29]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [29]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [29]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [29]));  // al_ip/div_unsigned_gate.v(597)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5793450  (
    .a(n34[1]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [33]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [32]));  // al_ip/div_unsigned_gate.v(169)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5793560  (
    .a(n34[11]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [43]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [42]));  // al_ip/div_unsigned_gate.v(185)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5793670  (
    .a(n34[8]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [40]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [39]));  // al_ip/div_unsigned_gate.v(794)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5793780  (
    .a(n35[12]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [12]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [12]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [12]));  // al_ip/div_unsigned_gate.v(401)
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'b00000000000000000000000000000010),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5794000  (
    .a(\u_DIV_UNSIGNED/al_00000286E4688A90 ),
    .b(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [0]),
    .c(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [3]),
    .d(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [4]),
    .e(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [5]),
    .o(\u_DIV_UNSIGNED/al_00000286E468A980 ));  // al_ip/div_unsigned_gate.v(722)
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'b00000000000010000000000000000000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5794220  (
    .a(\u_DIV_UNSIGNED/al_00000286E4688A90 ),
    .b(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [0]),
    .c(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [3]),
    .d(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [4]),
    .e(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [5]),
    .o(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ));  // al_ip/div_unsigned_gate.v(712)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_UNSIGNED/al_00000286E5794770  (
    .a(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .b(\u_DIV_UNSIGNED/al_00000286E468A980 ),
    .c(div_unsigned_start),
    .d(\u_DIV_UNSIGNED/al_00000286E57E03C0 [5]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E04A0 [5]));  // al_ip/div_unsigned_gate.v(732)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_UNSIGNED/al_00000286E5795540  (
    .a(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .b(\u_DIV_UNSIGNED/al_00000286E468A980 ),
    .c(div_unsigned_start),
    .d(\u_DIV_UNSIGNED/al_00000286E57E03C0 [3]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E04A0 [3]));  // al_ip/div_unsigned_gate.v(750)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_UNSIGNED/al_00000286E5796530  (
    .a(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .b(\u_DIV_UNSIGNED/al_00000286E468A980 ),
    .c(div_unsigned_start),
    .d(\u_DIV_UNSIGNED/al_00000286E57E03C0 [1]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E04A0 [1]));  // al_ip/div_unsigned_gate.v(776)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_UNSIGNED/al_00000286E5796A80  (
    .a(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .b(\u_DIV_UNSIGNED/al_00000286E468A980 ),
    .c(div_unsigned_start),
    .d(\u_DIV_UNSIGNED/al_00000286E57E03C0 [4]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E04A0 [4]));  // al_ip/div_unsigned_gate.v(741)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_UNSIGNED/al_00000286E5797740  (
    .a(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .b(\u_DIV_UNSIGNED/al_00000286E468A980 ),
    .c(div_unsigned_start),
    .d(\u_DIV_UNSIGNED/al_00000286E57E03C0 [2]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E04A0 [2]));  // al_ip/div_unsigned_gate.v(759)
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~B*~A))"),
    .INIT(16'b1111000111110000))
    \u_DIV_UNSIGNED/al_00000286E5797B80  (
    .a(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .b(\u_DIV_UNSIGNED/al_00000286E468A980 ),
    .c(div_unsigned_start),
    .d(\u_DIV_UNSIGNED/al_00000286E57E03C0 [0]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E04A0 [0]));  // al_ip/div_unsigned_gate.v(785)
  AL_DFF_X working_reg (
    .ar(~i_rstn),
    .as(1'b0),
    .clk(i_clk),
    .d(n8),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(working));  // ../RTL/core/exu_mdu.v(52)

endmodule 

module binary_mux_s5_w1
  (
  i0,
  i1,
  i10,
  i11,
  i12,
  i13,
  i14,
  i15,
  i16,
  i17,
  i18,
  i19,
  i2,
  i20,
  i21,
  i22,
  i23,
  i24,
  i25,
  i26,
  i27,
  i28,
  i29,
  i3,
  i30,
  i31,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  sel,
  o
  );

  input i0;
  input i1;
  input i10;
  input i11;
  input i12;
  input i13;
  input i14;
  input i15;
  input i16;
  input i17;
  input i18;
  input i19;
  input i2;
  input i20;
  input i21;
  input i22;
  input i23;
  input i24;
  input i25;
  input i26;
  input i27;
  input i28;
  input i29;
  input i3;
  input i30;
  input i31;
  input i4;
  input i5;
  input i6;
  input i7;
  input i8;
  input i9;
  input [4:0] sel;
  output o;

  wire  B0_0;
  wire  B0_1;
  wire  B0_10;
  wire  B0_11;
  wire  B0_12;
  wire  B0_13;
  wire  B0_14;
  wire  B0_15;
  wire  B0_2;
  wire  B0_3;
  wire  B0_4;
  wire  B0_5;
  wire  B0_6;
  wire  B0_7;
  wire  B0_8;
  wire  B0_9;
  wire  B1_0;
  wire  B1_1;
  wire  B1_2;
  wire  B1_3;
  wire  B1_4;
  wire  B1_5;
  wire  B1_6;
  wire  B1_7;
  wire  B2_0;
  wire  B2_1;
  wire  B2_2;
  wire  B2_3;
  wire  B3_0;
  wire  B3_1;

  AL_MUX al_mux_b0_0_0 (
    .i0(i0),
    .i1(i1),
    .sel(sel[0]),
    .o(B0_0));
  AL_MUX al_mux_b0_0_1 (
    .i0(i2),
    .i1(i3),
    .sel(sel[0]),
    .o(B0_1));
  AL_MUX al_mux_b0_0_10 (
    .i0(i20),
    .i1(i21),
    .sel(sel[0]),
    .o(B0_10));
  AL_MUX al_mux_b0_0_11 (
    .i0(i22),
    .i1(i23),
    .sel(sel[0]),
    .o(B0_11));
  AL_MUX al_mux_b0_0_12 (
    .i0(i24),
    .i1(i25),
    .sel(sel[0]),
    .o(B0_12));
  AL_MUX al_mux_b0_0_13 (
    .i0(i26),
    .i1(i27),
    .sel(sel[0]),
    .o(B0_13));
  AL_MUX al_mux_b0_0_14 (
    .i0(i28),
    .i1(i29),
    .sel(sel[0]),
    .o(B0_14));
  AL_MUX al_mux_b0_0_15 (
    .i0(i30),
    .i1(i31),
    .sel(sel[0]),
    .o(B0_15));
  AL_MUX al_mux_b0_0_2 (
    .i0(i4),
    .i1(i5),
    .sel(sel[0]),
    .o(B0_2));
  AL_MUX al_mux_b0_0_3 (
    .i0(i6),
    .i1(i7),
    .sel(sel[0]),
    .o(B0_3));
  AL_MUX al_mux_b0_0_4 (
    .i0(i8),
    .i1(i9),
    .sel(sel[0]),
    .o(B0_4));
  AL_MUX al_mux_b0_0_5 (
    .i0(i10),
    .i1(i11),
    .sel(sel[0]),
    .o(B0_5));
  AL_MUX al_mux_b0_0_6 (
    .i0(i12),
    .i1(i13),
    .sel(sel[0]),
    .o(B0_6));
  AL_MUX al_mux_b0_0_7 (
    .i0(i14),
    .i1(i15),
    .sel(sel[0]),
    .o(B0_7));
  AL_MUX al_mux_b0_0_8 (
    .i0(i16),
    .i1(i17),
    .sel(sel[0]),
    .o(B0_8));
  AL_MUX al_mux_b0_0_9 (
    .i0(i18),
    .i1(i19),
    .sel(sel[0]),
    .o(B0_9));
  AL_MUX al_mux_b0_1_0 (
    .i0(B0_0),
    .i1(B0_1),
    .sel(sel[1]),
    .o(B1_0));
  AL_MUX al_mux_b0_1_1 (
    .i0(B0_2),
    .i1(B0_3),
    .sel(sel[1]),
    .o(B1_1));
  AL_MUX al_mux_b0_1_2 (
    .i0(B0_4),
    .i1(B0_5),
    .sel(sel[1]),
    .o(B1_2));
  AL_MUX al_mux_b0_1_3 (
    .i0(B0_6),
    .i1(B0_7),
    .sel(sel[1]),
    .o(B1_3));
  AL_MUX al_mux_b0_1_4 (
    .i0(B0_8),
    .i1(B0_9),
    .sel(sel[1]),
    .o(B1_4));
  AL_MUX al_mux_b0_1_5 (
    .i0(B0_10),
    .i1(B0_11),
    .sel(sel[1]),
    .o(B1_5));
  AL_MUX al_mux_b0_1_6 (
    .i0(B0_12),
    .i1(B0_13),
    .sel(sel[1]),
    .o(B1_6));
  AL_MUX al_mux_b0_1_7 (
    .i0(B0_14),
    .i1(B0_15),
    .sel(sel[1]),
    .o(B1_7));
  AL_MUX al_mux_b0_2_0 (
    .i0(B1_0),
    .i1(B1_1),
    .sel(sel[2]),
    .o(B2_0));
  AL_MUX al_mux_b0_2_1 (
    .i0(B1_2),
    .i1(B1_3),
    .sel(sel[2]),
    .o(B2_1));
  AL_MUX al_mux_b0_2_2 (
    .i0(B1_4),
    .i1(B1_5),
    .sel(sel[2]),
    .o(B2_2));
  AL_MUX al_mux_b0_2_3 (
    .i0(B1_6),
    .i1(B1_7),
    .sel(sel[2]),
    .o(B2_3));
  AL_MUX al_mux_b0_3_0 (
    .i0(B2_0),
    .i1(B2_1),
    .sel(sel[3]),
    .o(B3_0));
  AL_MUX al_mux_b0_3_1 (
    .i0(B2_2),
    .i1(B2_3),
    .sel(sel[3]),
    .o(B3_1));
  AL_MUX al_mux_b0_4_0 (
    .i0(B3_0),
    .i1(B3_1),
    .sel(sel[4]),
    .o(o));

endmodule 

module add_sub_1  // ../RTL/core/fpu.v(83)
  (
  n1,
  n2,
  sub,
  Exception,
  Overflow,
  Underflow,
  result
  );

  input [31:0] n1;  // ../RTL/core/fpu.v(84)
  input [31:0] n2;  // ../RTL/core/fpu.v(85)
  input sub;  // ../RTL/core/fpu.v(87)
  output Exception;  // ../RTL/core/fpu.v(90)
  output Overflow;  // ../RTL/core/fpu.v(88)
  output Underflow;  // ../RTL/core/fpu.v(89)
  output [31:0] result;  // ../RTL/core/fpu.v(86)

  wire [7:0] \C023/outtemp ;  // ../RTL/core/fpu_utils.v(93)
  wire [23:0] \C03/outtemp ;  // ../RTL/core/fpu_utils.v(99)
  wire [7:0] E;  // ../RTL/core/fpu.v(95)
  wire [23:0] M1;  // ../RTL/core/fpu.v(97)
  wire [23:0] M2;  // ../RTL/core/fpu.v(97)
  wire [23:0] M_result;  // ../RTL/core/fpu.v(97)
  wire [23:0] M_result2;  // ../RTL/core/fpu.v(97)
  wire [22:0] \NM/n122 ;
  wire [22:0] \NM/n4 ;
  wire  \NM/sel0_b1/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b1/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B13_al_b40 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B12_al_b39 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B13_al_b40 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B11_al_b38 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B12_al_b39 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B13_al_b40 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B10_al_b37 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B11_al_b38 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B12_al_b39 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B13_al_b40 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B10_al_b37 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B11_al_b38 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B12_al_b39 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B13_al_b40 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B9_al_b36 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B10_al_b37 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B11_al_b38 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B12_al_b39 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B13_al_b40 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B8_al_b35 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B9_al_b36 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B10_al_b37 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B11_al_b38 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B12_al_b39 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B13_al_b40 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B7_al_b34 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B8_al_b35 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B9_al_b36 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B10_al_b37 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B11_al_b38 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B12_al_b39 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B13_al_b40 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B6_al_b33 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B7_al_b34 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B8_al_b35 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B9_al_b36 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B10_al_b37 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B11_al_b38 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B12_al_b39 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B13_al_b40 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B5_al_b32 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B6_al_b33 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B7_al_b34 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B8_al_b35 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B9_al_b36 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b2/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b2/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b2/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B10_al_b37 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B11_al_b38 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B12_al_b39 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B13_al_b40 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B4_al_b31 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B5_al_b32 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B6_al_b33 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B7_al_b34 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B8_al_b35 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B9_al_b36 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B10_al_b37 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B11_al_b38 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B12_al_b39 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B13_al_b40 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B3_al_b30 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B4_al_b31 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B5_al_b32 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B6_al_b33 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B7_al_b34 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B8_al_b35 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B9_al_b36 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B10_al_b37 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B11_al_b38 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B12_al_b39 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B13_al_b40 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B14_al_b41 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B2_al_b29 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B3_al_b30 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B4_al_b31 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B5_al_b32 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B6_al_b33 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B7_al_b34 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B8_al_b35 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B9_al_b36 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b3/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b3/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b3/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b3/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b4/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b4/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b4/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b4/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b4/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b5/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b5/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b5/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b5/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b5/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b5/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B15_al_b42 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B16_al_b43 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B17_al_b44 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B18_al_b45 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B19_al_b46 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B20_al_b47 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B21_al_b48 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B22_al_b49 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B23_al_b50 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B24_al_b51 ;  // ../RTL/core/fpu_utils.v(163)
  wire [7:0] One_Added_E;  // ../RTL/core/fpu.v(95)
  wire [7:0] complemented_E2;  // ../RTL/core/fpu.v(95)
  wire [23:0] complemented_M_result;  // ../RTL/core/fpu.v(97)
  wire [7:0] complemented_shift_E;  // ../RTL/core/fpu.v(95)
  wire [7:0] complemented_temp_exp_diff;  // ../RTL/core/fpu.v(95)
  wire [7:0] exp_diff;  // ../RTL/core/fpu.v(95)
  wire [23:0] n37;
  wire [23:0] n62;
  wire [7:0] new_E;  // ../RTL/core/fpu.v(95)
  wire [23:0] new_M2;  // ../RTL/core/fpu.v(97)
  wire [4:0] shift_E;  // ../RTL/core/fpu.v(100)
  wire [7:0] temp_exp_diff;  // ../RTL/core/fpu.v(95)
  wire \ADD01/ADD01/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/n1 ;
  wire \ADD01/ADD01/n10 ;
  wire \ADD01/ADD01/n12 ;
  wire \ADD01/ADD01/n13 ;
  wire \ADD01/ADD01/n14 ;
  wire \ADD01/ADD01/n15 ;
  wire \ADD01/ADD01/n16 ;
  wire \ADD01/ADD01/n17 ;
  wire \ADD01/ADD01/n18 ;
  wire \ADD01/ADD01/n19 ;
  wire \ADD01/ADD01/n2 ;
  wire \ADD01/ADD01/n20 ;
  wire \ADD01/ADD01/n3 ;
  wire \ADD01/ADD01/n5 ;
  wire \ADD01/ADD01/n6 ;
  wire \ADD01/ADD01/n7 ;
  wire \ADD01/ADD01/n8 ;
  wire \ADD01/ADD01/n9 ;
  wire \ADD01/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/p0_neg ;
  wire \ADD01/ADD01/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/n0 ;
  wire \ADD01/ADD02/n1 ;
  wire \ADD01/ADD02/n10 ;
  wire \ADD01/ADD02/n11 ;
  wire \ADD01/ADD02/n12 ;
  wire \ADD01/ADD02/n13 ;
  wire \ADD01/ADD02/n14 ;
  wire \ADD01/ADD02/n15 ;
  wire \ADD01/ADD02/n16 ;
  wire \ADD01/ADD02/n17 ;
  wire \ADD01/ADD02/n18 ;
  wire \ADD01/ADD02/n19 ;
  wire \ADD01/ADD02/n2 ;
  wire \ADD01/ADD02/n20 ;
  wire \ADD01/ADD02/n21 ;
  wire \ADD01/ADD02/n3 ;
  wire \ADD01/ADD02/n4 ;
  wire \ADD01/ADD02/n5 ;
  wire \ADD01/ADD02/n6 ;
  wire \ADD01/ADD02/n7 ;
  wire \ADD01/ADD02/n8 ;
  wire \ADD01/ADD02/n9 ;
  wire \ADD01/ADD02/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ctemp ;  // ../RTL/core/fpu_utils.v(76)
  wire \ADD02/ADD01/ADD01/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/n0 ;
  wire \ADD02/ADD01/ADD01/n1 ;
  wire \ADD02/ADD01/ADD01/n10 ;
  wire \ADD02/ADD01/ADD01/n11 ;
  wire \ADD02/ADD01/ADD01/n12 ;
  wire \ADD02/ADD01/ADD01/n13 ;
  wire \ADD02/ADD01/ADD01/n14 ;
  wire \ADD02/ADD01/ADD01/n15 ;
  wire \ADD02/ADD01/ADD01/n16 ;
  wire \ADD02/ADD01/ADD01/n17 ;
  wire \ADD02/ADD01/ADD01/n18 ;
  wire \ADD02/ADD01/ADD01/n19 ;
  wire \ADD02/ADD01/ADD01/n2 ;
  wire \ADD02/ADD01/ADD01/n20 ;
  wire \ADD02/ADD01/ADD01/n21 ;
  wire \ADD02/ADD01/ADD01/n3 ;
  wire \ADD02/ADD01/ADD01/n4 ;
  wire \ADD02/ADD01/ADD01/n5 ;
  wire \ADD02/ADD01/ADD01/n6 ;
  wire \ADD02/ADD01/ADD01/n7 ;
  wire \ADD02/ADD01/ADD01/n8 ;
  wire \ADD02/ADD01/ADD01/n9 ;
  wire \ADD02/ADD01/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/n0 ;
  wire \ADD02/ADD01/ADD02/n1 ;
  wire \ADD02/ADD01/ADD02/n10 ;
  wire \ADD02/ADD01/ADD02/n11 ;
  wire \ADD02/ADD01/ADD02/n12 ;
  wire \ADD02/ADD01/ADD02/n13 ;
  wire \ADD02/ADD01/ADD02/n14 ;
  wire \ADD02/ADD01/ADD02/n15 ;
  wire \ADD02/ADD01/ADD02/n16 ;
  wire \ADD02/ADD01/ADD02/n17 ;
  wire \ADD02/ADD01/ADD02/n18 ;
  wire \ADD02/ADD01/ADD02/n19 ;
  wire \ADD02/ADD01/ADD02/n2 ;
  wire \ADD02/ADD01/ADD02/n20 ;
  wire \ADD02/ADD01/ADD02/n21 ;
  wire \ADD02/ADD01/ADD02/n3 ;
  wire \ADD02/ADD01/ADD02/n4 ;
  wire \ADD02/ADD01/ADD02/n5 ;
  wire \ADD02/ADD01/ADD02/n6 ;
  wire \ADD02/ADD01/ADD02/n7 ;
  wire \ADD02/ADD01/ADD02/n8 ;
  wire \ADD02/ADD01/ADD02/n9 ;
  wire \ADD02/ADD01/ADD02/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ctemp ;  // ../RTL/core/fpu_utils.v(76)
  wire \ADD02/ADD02/ADD01/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/n0 ;
  wire \ADD02/ADD02/ADD01/n1 ;
  wire \ADD02/ADD02/ADD01/n10 ;
  wire \ADD02/ADD02/ADD01/n11 ;
  wire \ADD02/ADD02/ADD01/n12 ;
  wire \ADD02/ADD02/ADD01/n13 ;
  wire \ADD02/ADD02/ADD01/n14 ;
  wire \ADD02/ADD02/ADD01/n15 ;
  wire \ADD02/ADD02/ADD01/n16 ;
  wire \ADD02/ADD02/ADD01/n17 ;
  wire \ADD02/ADD02/ADD01/n18 ;
  wire \ADD02/ADD02/ADD01/n19 ;
  wire \ADD02/ADD02/ADD01/n2 ;
  wire \ADD02/ADD02/ADD01/n20 ;
  wire \ADD02/ADD02/ADD01/n21 ;
  wire \ADD02/ADD02/ADD01/n3 ;
  wire \ADD02/ADD02/ADD01/n4 ;
  wire \ADD02/ADD02/ADD01/n5 ;
  wire \ADD02/ADD02/ADD01/n6 ;
  wire \ADD02/ADD02/ADD01/n7 ;
  wire \ADD02/ADD02/ADD01/n8 ;
  wire \ADD02/ADD02/ADD01/n9 ;
  wire \ADD02/ADD02/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/n0 ;
  wire \ADD02/ADD02/ADD02/n1 ;
  wire \ADD02/ADD02/ADD02/n10 ;
  wire \ADD02/ADD02/ADD02/n11 ;
  wire \ADD02/ADD02/ADD02/n12 ;
  wire \ADD02/ADD02/ADD02/n13 ;
  wire \ADD02/ADD02/ADD02/n14 ;
  wire \ADD02/ADD02/ADD02/n15 ;
  wire \ADD02/ADD02/ADD02/n16 ;
  wire \ADD02/ADD02/ADD02/n17 ;
  wire \ADD02/ADD02/ADD02/n18 ;
  wire \ADD02/ADD02/ADD02/n19 ;
  wire \ADD02/ADD02/ADD02/n2 ;
  wire \ADD02/ADD02/ADD02/n20 ;
  wire \ADD02/ADD02/ADD02/n21 ;
  wire \ADD02/ADD02/ADD02/n3 ;
  wire \ADD02/ADD02/ADD02/n4 ;
  wire \ADD02/ADD02/ADD02/n5 ;
  wire \ADD02/ADD02/ADD02/n6 ;
  wire \ADD02/ADD02/ADD02/n7 ;
  wire \ADD02/ADD02/ADD02/n8 ;
  wire \ADD02/ADD02/ADD02/n9 ;
  wire \ADD02/ADD02/ADD02/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ctemp ;  // ../RTL/core/fpu_utils.v(76)
  wire \ADD02/ADD03/ADD01/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/n0 ;
  wire \ADD02/ADD03/ADD01/n1 ;
  wire \ADD02/ADD03/ADD01/n10 ;
  wire \ADD02/ADD03/ADD01/n11 ;
  wire \ADD02/ADD03/ADD01/n12 ;
  wire \ADD02/ADD03/ADD01/n13 ;
  wire \ADD02/ADD03/ADD01/n14 ;
  wire \ADD02/ADD03/ADD01/n15 ;
  wire \ADD02/ADD03/ADD01/n16 ;
  wire \ADD02/ADD03/ADD01/n17 ;
  wire \ADD02/ADD03/ADD01/n18 ;
  wire \ADD02/ADD03/ADD01/n19 ;
  wire \ADD02/ADD03/ADD01/n2 ;
  wire \ADD02/ADD03/ADD01/n20 ;
  wire \ADD02/ADD03/ADD01/n21 ;
  wire \ADD02/ADD03/ADD01/n3 ;
  wire \ADD02/ADD03/ADD01/n4 ;
  wire \ADD02/ADD03/ADD01/n5 ;
  wire \ADD02/ADD03/ADD01/n6 ;
  wire \ADD02/ADD03/ADD01/n7 ;
  wire \ADD02/ADD03/ADD01/n8 ;
  wire \ADD02/ADD03/ADD01/n9 ;
  wire \ADD02/ADD03/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/n0 ;
  wire \ADD02/ADD03/ADD02/n1 ;
  wire \ADD02/ADD03/ADD02/n10 ;
  wire \ADD02/ADD03/ADD02/n11 ;
  wire \ADD02/ADD03/ADD02/n12 ;
  wire \ADD02/ADD03/ADD02/n13 ;
  wire \ADD02/ADD03/ADD02/n14 ;
  wire \ADD02/ADD03/ADD02/n15 ;
  wire \ADD02/ADD03/ADD02/n16 ;
  wire \ADD02/ADD03/ADD02/n17 ;
  wire \ADD02/ADD03/ADD02/n18 ;
  wire \ADD02/ADD03/ADD02/n19 ;
  wire \ADD02/ADD03/ADD02/n2 ;
  wire \ADD02/ADD03/ADD02/n20 ;
  wire \ADD02/ADD03/ADD02/n21 ;
  wire \ADD02/ADD03/ADD02/n3 ;
  wire \ADD02/ADD03/ADD02/n4 ;
  wire \ADD02/ADD03/ADD02/n5 ;
  wire \ADD02/ADD03/ADD02/n6 ;
  wire \ADD02/ADD03/ADD02/n7 ;
  wire \ADD02/ADD03/ADD02/n8 ;
  wire \ADD02/ADD03/ADD02/n9 ;
  wire \ADD02/ADD03/ADD02/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ctemp ;  // ../RTL/core/fpu_utils.v(76)
  wire \ADD02/ctemp1 ;  // ../RTL/core/fpu_utils.v(87)
  wire \ADD02/ctemp2 ;  // ../RTL/core/fpu_utils.v(88)
  wire \ADD0212/ADD01/n1 ;
  wire \ADD0212/ADD01/n14 ;
  wire \ADD0212/ADD01/n17 ;
  wire \ADD0212/ADD01/n18 ;
  wire \ADD0212/ADD01/n7 ;
  wire \ADD0212/ADD01/n8 ;
  wire \ADD0212/ADD02/n0 ;
  wire \ADD0212/ADD02/n10 ;
  wire \ADD0212/ADD02/n11 ;
  wire \ADD0212/ADD02/n3 ;
  wire \ADD0212/ADD02/n4 ;
  wire \ADD0212/ADD02/n7 ;
  wire \ADD03/ADD01/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/n1 ;
  wire \ADD03/ADD01/n10 ;
  wire \ADD03/ADD01/n12 ;
  wire \ADD03/ADD01/n13 ;
  wire \ADD03/ADD01/n14 ;
  wire \ADD03/ADD01/n15 ;
  wire \ADD03/ADD01/n16 ;
  wire \ADD03/ADD01/n17 ;
  wire \ADD03/ADD01/n18 ;
  wire \ADD03/ADD01/n19 ;
  wire \ADD03/ADD01/n2 ;
  wire \ADD03/ADD01/n20 ;
  wire \ADD03/ADD01/n3 ;
  wire \ADD03/ADD01/n5 ;
  wire \ADD03/ADD01/n6 ;
  wire \ADD03/ADD01/n7 ;
  wire \ADD03/ADD01/n8 ;
  wire \ADD03/ADD01/n9 ;
  wire \ADD03/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/p0_neg ;
  wire \ADD03/ADD01/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD02/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD02/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD02/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD02/n0 ;
  wire \ADD03/ADD02/n1 ;
  wire \ADD03/ADD02/n10 ;
  wire \ADD03/ADD02/n11 ;
  wire \ADD03/ADD02/n2 ;
  wire \ADD03/ADD02/n3 ;
  wire \ADD03/ADD02/n4 ;
  wire \ADD03/ADD02/n5 ;
  wire \ADD03/ADD02/n6 ;
  wire \ADD03/ADD02/n7 ;
  wire \ADD03/ADD02/n8 ;
  wire \ADD03/ADD02/n9 ;
  wire \ADD03/ADD02/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ctemp ;  // ../RTL/core/fpu_utils.v(76)
  wire \C023/ADD01/ADD01/n1 ;
  wire \C023/ADD01/ADD01/n14 ;
  wire \C023/ADD01/ADD01/n17 ;
  wire \C023/ADD01/ADD01/n18 ;
  wire \C023/ADD01/ADD01/n7 ;
  wire \C023/ADD01/ADD01/n8 ;
  wire \C023/ADD01/ADD02/n0 ;
  wire \C023/ADD01/ADD02/n10 ;
  wire \C023/ADD01/ADD02/n11 ;
  wire \C023/ADD01/ADD02/n3 ;
  wire \C023/ADD01/ADD02/n4 ;
  wire \C023/ADD01/ADD02/n7 ;
  wire \C03/ADD01/ADD01/ADD01/n1 ;
  wire \C03/ADD01/ADD01/ADD01/n14 ;
  wire \C03/ADD01/ADD01/ADD01/n17 ;
  wire \C03/ADD01/ADD01/ADD01/n18 ;
  wire \C03/ADD01/ADD01/ADD01/n7 ;
  wire \C03/ADD01/ADD01/ADD01/n8 ;
  wire \C03/ADD01/ADD01/ADD02/n0 ;
  wire \C03/ADD01/ADD01/ADD02/n10 ;
  wire \C03/ADD01/ADD01/ADD02/n11 ;
  wire \C03/ADD01/ADD01/ADD02/n14 ;
  wire \C03/ADD01/ADD01/ADD02/n17 ;
  wire \C03/ADD01/ADD01/ADD02/n20 ;
  wire \C03/ADD01/ADD01/ADD02/n21 ;
  wire \C03/ADD01/ADD01/ADD02/n3 ;
  wire \C03/ADD01/ADD01/ADD02/n4 ;
  wire \C03/ADD01/ADD01/ADD02/n7 ;
  wire \C03/ADD01/ADD02/ADD01/n0 ;
  wire \C03/ADD01/ADD02/ADD01/n10 ;
  wire \C03/ADD01/ADD02/ADD01/n11 ;
  wire \C03/ADD01/ADD02/ADD01/n14 ;
  wire \C03/ADD01/ADD02/ADD01/n17 ;
  wire \C03/ADD01/ADD02/ADD01/n20 ;
  wire \C03/ADD01/ADD02/ADD01/n21 ;
  wire \C03/ADD01/ADD02/ADD01/n3 ;
  wire \C03/ADD01/ADD02/ADD01/n4 ;
  wire \C03/ADD01/ADD02/ADD01/n7 ;
  wire \C03/ADD01/ADD02/ADD02/n0 ;
  wire \C03/ADD01/ADD02/ADD02/n10 ;
  wire \C03/ADD01/ADD02/ADD02/n11 ;
  wire \C03/ADD01/ADD02/ADD02/n14 ;
  wire \C03/ADD01/ADD02/ADD02/n17 ;
  wire \C03/ADD01/ADD02/ADD02/n20 ;
  wire \C03/ADD01/ADD02/ADD02/n21 ;
  wire \C03/ADD01/ADD02/ADD02/n3 ;
  wire \C03/ADD01/ADD02/ADD02/n4 ;
  wire \C03/ADD01/ADD02/ADD02/n7 ;
  wire \C03/ADD01/ADD03/ADD01/n0 ;
  wire \C03/ADD01/ADD03/ADD01/n10 ;
  wire \C03/ADD01/ADD03/ADD01/n11 ;
  wire \C03/ADD01/ADD03/ADD01/n14 ;
  wire \C03/ADD01/ADD03/ADD01/n17 ;
  wire \C03/ADD01/ADD03/ADD01/n20 ;
  wire \C03/ADD01/ADD03/ADD01/n21 ;
  wire \C03/ADD01/ADD03/ADD01/n3 ;
  wire \C03/ADD01/ADD03/ADD01/n4 ;
  wire \C03/ADD01/ADD03/ADD01/n7 ;
  wire \C03/ADD01/ADD03/ADD02/n0 ;
  wire \C03/ADD01/ADD03/ADD02/n10 ;
  wire \C03/ADD01/ADD03/ADD02/n11 ;
  wire \C03/ADD01/ADD03/ADD02/n3 ;
  wire \C03/ADD01/ADD03/ADD02/n4 ;
  wire \C03/ADD01/ADD03/ADD02/n7 ;
  wire \M031/M01/invSL ;  // ../RTL/core/fpu_utils.v(105)
  wire \M04/M01/M01/invSL ;  // ../RTL/core/fpu_utils.v(105)
  wire M_carry;  // ../RTL/core/fpu.v(93)
  wire \NM/mux1_b0_sel_is_2_o ;
  wire \NM/mux1_b1_sel_is_2_o ;
  wire \NM/mux1_b2_sel_is_2_o ;
  wire \NM/mux1_b3_sel_is_2_o ;
  wire \NM/mux1_b4_sel_is_2_o ;
  wire \NM/n10 ;
  wire \NM/n100 ;
  wire \NM/n101 ;
  wire \NM/n102 ;
  wire \NM/n103 ;
  wire \NM/n104 ;
  wire \NM/n105 ;
  wire \NM/n106 ;
  wire \NM/n107 ;
  wire \NM/n108 ;
  wire \NM/n109 ;
  wire \NM/n11 ;
  wire \NM/n110 ;
  wire \NM/n111 ;
  wire \NM/n112 ;
  wire \NM/n113 ;
  wire \NM/n114 ;
  wire \NM/n115 ;
  wire \NM/n116 ;
  wire \NM/n117 ;
  wire \NM/n118 ;
  wire \NM/n119 ;
  wire \NM/n12 ;
  wire \NM/n124 ;
  wire \NM/n125 ;
  wire \NM/n126 ;
  wire \NM/n127 ;
  wire \NM/n128 ;
  wire \NM/n129 ;
  wire \NM/n13 ;
  wire \NM/n130 ;
  wire \NM/n132 ;
  wire \NM/n133 ;
  wire \NM/n134 ;
  wire \NM/n14 ;
  wire \NM/n142 ;
  wire \NM/n143 ;
  wire \NM/n146 ;
  wire \NM/n15 ;
  wire \NM/n153 ;
  wire \NM/n156 ;
  wire \NM/n158 ;
  wire \NM/n16 ;
  wire \NM/n165 ;
  wire \NM/n166 ;
  wire \NM/n168 ;
  wire \NM/n17 ;
  wire \NM/n170 ;
  wire \NM/n171 ;
  wire \NM/n175 ;
  wire \NM/n176 ;
  wire \NM/n177 ;
  wire \NM/n179 ;
  wire \NM/n18 ;
  wire \NM/n180 ;
  wire \NM/n182 ;
  wire \NM/n183 ;
  wire \NM/n184 ;
  wire \NM/n185 ;
  wire \NM/n186 ;
  wire \NM/n187 ;
  wire \NM/n188 ;
  wire \NM/n189 ;
  wire \NM/n19 ;
  wire \NM/n190 ;
  wire \NM/n191 ;
  wire \NM/n193 ;
  wire \NM/n194 ;
  wire \NM/n195 ;
  wire \NM/n2 ;
  wire \NM/n20 ;
  wire \NM/n202 ;
  wire \NM/n207 ;
  wire \NM/n209 ;
  wire \NM/n21 ;
  wire \NM/n210 ;
  wire \NM/n211 ;
  wire \NM/n213 ;
  wire \NM/n214 ;
  wire \NM/n215 ;
  wire \NM/n216 ;
  wire \NM/n22 ;
  wire \NM/n222 ;
  wire \NM/n227 ;
  wire \NM/n23 ;
  wire \NM/n230 ;
  wire \NM/n232 ;
  wire \NM/n234 ;
  wire \NM/n236 ;
  wire \NM/n24 ;
  wire \NM/n240 ;
  wire \NM/n242 ;
  wire \NM/n243 ;
  wire \NM/n244 ;
  wire \NM/n246 ;
  wire \NM/n247 ;
  wire \NM/n248 ;
  wire \NM/n249 ;
  wire \NM/n25 ;
  wire \NM/n251 ;
  wire \NM/n253 ;
  wire \NM/n257 ;
  wire \NM/n258 ;
  wire \NM/n26 ;
  wire \NM/n260 ;
  wire \NM/n261 ;
  wire \NM/n262 ;
  wire \NM/n263 ;
  wire \NM/n265 ;
  wire \NM/n268 ;
  wire \NM/n269 ;
  wire \NM/n27 ;
  wire \NM/n271 ;
  wire \NM/n273 ;
  wire \NM/n274 ;
  wire \NM/n276 ;
  wire \NM/n278 ;
  wire \NM/n279 ;
  wire \NM/n28 ;
  wire \NM/n280 ;
  wire \NM/n281 ;
  wire \NM/n283 ;
  wire \NM/n284 ;
  wire \NM/n286 ;
  wire \NM/n29 ;
  wire \NM/n296 ;
  wire \NM/n30 ;
  wire \NM/n300 ;
  wire \NM/n304 ;
  wire \NM/n306 ;
  wire \NM/n308 ;
  wire \NM/n31 ;
  wire \NM/n310 ;
  wire \NM/n311 ;
  wire \NM/n312 ;
  wire \NM/n313 ;
  wire \NM/n314 ;
  wire \NM/n315 ;
  wire \NM/n316 ;
  wire \NM/n318 ;
  wire \NM/n319 ;
  wire \NM/n32 ;
  wire \NM/n320 ;
  wire \NM/n321 ;
  wire \NM/n322 ;
  wire \NM/n325 ;
  wire \NM/n33 ;
  wire \NM/n331 ;
  wire \NM/n332 ;
  wire \NM/n335 ;
  wire \NM/n34 ;
  wire \NM/n340 ;
  wire \NM/n341 ;
  wire \NM/n343 ;
  wire \NM/n348 ;
  wire \NM/n349 ;
  wire \NM/n35 ;
  wire \NM/n351 ;
  wire \NM/n355 ;
  wire \NM/n357 ;
  wire \NM/n36 ;
  wire \NM/n361 ;
  wire \NM/n363 ;
  wire \NM/n366 ;
  wire \NM/n367 ;
  wire \NM/n37 ;
  wire \NM/n370 ;
  wire \NM/n371 ;
  wire \NM/n373 ;
  wire \NM/n374 ;
  wire \NM/n375 ;
  wire \NM/n376 ;
  wire \NM/n38 ;
  wire \NM/n39 ;
  wire \NM/n40 ;
  wire \NM/n41 ;
  wire \NM/n42 ;
  wire \NM/n44 ;
  wire \NM/n45 ;
  wire \NM/n46 ;
  wire \NM/n47 ;
  wire \NM/n48 ;
  wire \NM/n49 ;
  wire \NM/n50 ;
  wire \NM/n51 ;
  wire \NM/n52 ;
  wire \NM/n53 ;
  wire \NM/n54 ;
  wire \NM/n55 ;
  wire \NM/n56 ;
  wire \NM/n57 ;
  wire \NM/n58 ;
  wire \NM/n59 ;
  wire \NM/n6 ;
  wire \NM/n60 ;
  wire \NM/n61 ;
  wire \NM/n62 ;
  wire \NM/n63 ;
  wire \NM/n64 ;
  wire \NM/n65 ;
  wire \NM/n66 ;
  wire \NM/n67 ;
  wire \NM/n68 ;
  wire \NM/n69 ;
  wire \NM/n7 ;
  wire \NM/n70 ;
  wire \NM/n71 ;
  wire \NM/n72 ;
  wire \NM/n73 ;
  wire \NM/n74 ;
  wire \NM/n75 ;
  wire \NM/n76 ;
  wire \NM/n77 ;
  wire \NM/n78 ;
  wire \NM/n79 ;
  wire \NM/n8 ;
  wire \NM/n80 ;
  wire \NM/n81 ;
  wire \NM/n82 ;
  wire \NM/n83 ;
  wire \NM/n84 ;
  wire \NM/n85 ;
  wire \NM/n86 ;
  wire \NM/n87 ;
  wire \NM/n88 ;
  wire \NM/n89 ;
  wire \NM/n9 ;
  wire \NM/n90 ;
  wire \NM/n91 ;
  wire \NM/n92 ;
  wire \NM/n93 ;
  wire \NM/n94 ;
  wire \NM/n95 ;
  wire \NM/n96 ;
  wire \NM/n97 ;
  wire \NM/n98 ;
  wire \NM/n99 ;
  wire \NM/sel0_b1/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B13_al_b40_B14_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B12_al_b39_or_B13_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B13_al_b40_B14_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B12_al_b39_or_B13_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B13_al_b40_B14_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B10_al_b37_B11_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B12_al_b39_or_B13_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B13_al_b40_B14_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B10_al_b37_B11_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B12_al_b39_or_B13_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B13_al_b40_B14_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B9_al_b36_or_B10__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B10_al_b37_B11_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B12_al_b39_or_B13_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B13_al_b40_B14_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B9_al_b36_or_B10__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_or_B6_al_b33_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B10_al_b37_B11_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B12_al_b39_or_B13_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B13_al_b40_B14_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B7_al_b34_B8_al_b_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B9_al_b36_or_B10__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_or_B6_al_b33_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B10_al_b37_B11_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B12_al_b39_or_B13_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B13_al_b40_B14_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B6_al_b33_or_B7_a_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B7_al_b34_B8_al_b_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B9_al_b36_or_B10__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_or_B6_al_b33_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B10_al_b37_B11_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B12_al_b39_or_B13_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B13_al_b40_B14_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B6_al_b33_or_B7_a_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B7_al_b34_B8_al_b_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B9_al_b36_or_B10__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_or_B6_al_b33_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_or_or_B0_al_b27_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b2/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b2/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B10_al_b37_B11_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B12_al_b39_or_B13_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B13_al_b40_B14_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B4_al_b31_B5_al_b_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B6_al_b33_or_B7_a_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B7_al_b34_B8_al_b_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B9_al_b36_or_B10__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_or_B6_al_b33_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_or_or_B0_al_b27_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B10_al_b37_B11_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B12_al_b39_or_B13_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B13_al_b40_B14_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B3_al_b30_or_B4_a_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B4_al_b31_B5_al_b_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B6_al_b33_or_B7_a_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B7_al_b34_B8_al_b_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B9_al_b36_or_B10__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_or_B6_al_b33_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_or_or_B0_al_b27_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B10_al_b37_B11_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B12_al_b39_or_B13_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B13_al_b40_B14_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B3_al_b30_or_B4_a_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B4_al_b31_B5_al_b_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B6_al_b33_or_B7_a_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B7_al_b34_B8_al_b_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B9_al_b36_or_B10__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_B0_al_b27_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_B12_al_b39_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_B6_al_b33_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_or_B0_al_b27_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b3/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b3/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b3/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b4/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b4/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b4/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b4/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b5/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b5/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b5/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b5/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b5/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b6/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b6/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b6/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b6/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b6/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b6/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_B15_al_b42_or_B16_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_B16_al_b43_B17_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_B18_al_b45_or_B19_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_B19_al_b46_B20_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_B21_al_b48_B22_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_B23_al_b50_B24_al_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_or_B18_al_b45_or__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_or_B21_al_b48_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_or_or_B12_al_b39__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel1_b0_sel_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel1_b1_sel_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel1_b2_sel_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel1_b3_sel_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel1_b4_sel_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \RO01/w1 ;  // ../RTL/core/fpu_utils.v(13)
  wire \RO01/w2 ;  // ../RTL/core/fpu_utils.v(13)
  wire \RO01/w3 ;  // ../RTL/core/fpu_utils.v(13)
  wire \RO01/w4 ;  // ../RTL/core/fpu_utils.v(13)
  wire \RO01/w5 ;  // ../RTL/core/fpu_utils.v(13)
  wire \RO01/w6 ;  // ../RTL/core/fpu_utils.v(13)
  wire \exp_diff[4]_neg ;
  wire isE1GreaterThanE2;  // ../RTL/core/fpu.v(116)
  wire n10;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n11;
  wire n110;
  wire n110_neg;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n164;
  wire n165;
  wire n171;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n243;
  wire n244;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n265;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n5;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n6;
  wire n60;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n7;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n8;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n9;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire \new_E[5]_neg ;
  wire \new_E[6]_neg ;
  wire \new_E[7]_neg ;
  wire real_oper;  // ../RTL/core/fpu.v(93)
  wire reduced_or_E1;  // ../RTL/core/fpu.v(94)
  wire u194_sel_is_0_o;
  wire w1;  // ../RTL/core/fpu.v(98)
  wire w2;  // ../RTL/core/fpu.v(98)
  wire w3;  // ../RTL/core/fpu.v(98)

  assign result[23] = \ADD03/ADD01/p0_neg ;
  not \ADD01/ADD01/p0_inv  (\ADD01/ADD01/p0_neg , \ADD01/ADD01/p0 );
  and \ADD01/ADD01/u0  (\ADD01/ADD01/g0 , n1[23], complemented_E2[0]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD01/ADD01/u1  (\ADD01/ADD01/g1 , n1[24], complemented_E2[1]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD01/ADD01/u10  (\ADD01/ADD01/n1 , \ADD01/ADD01/p1 , \ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD01/ADD01/u11  (\ADD01/ADD01/n2 , \ADD01/ADD01/g1 , \ADD01/ADD01/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD01/ADD01/u12  (\ADD01/ADD01/n3 , \ADD01/ADD01/p1 , \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD01/ADD01/u14  (\ADD01/ADD01/c1 , \ADD01/ADD01/n2 , \ADD01/ADD01/n3 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD01/ADD01/u15  (\ADD01/ADD01/n5 , \ADD01/ADD01/p2 , \ADD01/ADD01/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD01/ADD01/u16  (\ADD01/ADD01/n6 , \ADD01/ADD01/g2 , \ADD01/ADD01/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD01/u17  (\ADD01/ADD01/n7 , \ADD01/ADD01/p2 , \ADD01/ADD01/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD01/u18  (\ADD01/ADD01/n8 , \ADD01/ADD01/n7 , \ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD01/ADD01/u19  (\ADD01/ADD01/n9 , \ADD01/ADD01/n6 , \ADD01/ADD01/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD01/u2  (\ADD01/ADD01/g2 , n1[25], complemented_E2[2]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD01/ADD01/u20  (temp_exp_diff[3], \ADD01/ADD01/p3 , \ADD01/ADD01/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD01/ADD01/u21  (\ADD01/ADD01/n10 , \ADD01/ADD01/n7 , \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD01/ADD01/u23  (\ADD01/ADD01/c2 , \ADD01/ADD01/n9 , \ADD01/ADD01/n10 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD01/u24  (\ADD01/ADD01/n12 , \ADD01/ADD01/p3 , \ADD01/ADD01/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD01/u25  (\ADD01/ADD01/n13 , \ADD01/ADD01/g3 , \ADD01/ADD01/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD01/u26  (\ADD01/ADD01/n14 , \ADD01/ADD01/p3 , \ADD01/ADD01/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD01/u27  (\ADD01/ADD01/n15 , \ADD01/ADD01/n14 , \ADD01/ADD01/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD01/u28  (\ADD01/ADD01/n16 , \ADD01/ADD01/n13 , \ADD01/ADD01/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD01/ADD01/u29  (temp_exp_diff[2], \ADD01/ADD01/p2 , \ADD01/ADD01/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD01/ADD01/u3  (\ADD01/ADD01/g3 , n1[26], complemented_E2[3]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD01/ADD01/u30  (\ADD01/ADD01/n17 , \ADD01/ADD01/n14 , \ADD01/ADD01/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD01/u31  (\ADD01/ADD01/n18 , \ADD01/ADD01/n17 , \ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD01/u32  (\ADD01/ADD01/n19 , \ADD01/ADD01/n16 , \ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD01/ADD01/u33  (temp_exp_diff[1], \ADD01/ADD01/p1 , \ADD01/ADD01/c0 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD01/ADD01/u35  (\ADD01/ADD01/n20 , \ADD01/ADD01/n17 , \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD01/u37  (\ADD01/ctemp , \ADD01/ADD01/n19 , \ADD01/ADD01/n20 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD01/ADD01/u4  (\ADD01/ADD01/p0 , n1[23], complemented_E2[0]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD01/ADD01/u5  (\ADD01/ADD01/p1 , n1[24], complemented_E2[1]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD01/ADD01/u6  (\ADD01/ADD01/p2 , n1[25], complemented_E2[2]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD01/ADD01/u7  (\ADD01/ADD01/p3 , n1[26], complemented_E2[3]);  // ../RTL/core/fpu_utils.v(62)
  or \ADD01/ADD01/u9  (\ADD01/ADD01/c0 , \ADD01/ADD01/g0 , \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD01/ADD02/u0  (\ADD01/ADD02/g0 , n1[27], complemented_E2[4]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD01/ADD02/u1  (\ADD01/ADD02/g1 , n1[28], complemented_E2[5]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD01/ADD02/u10  (\ADD01/ADD02/n1 , \ADD01/ADD02/p1 , \ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD01/ADD02/u11  (\ADD01/ADD02/n2 , \ADD01/ADD02/g1 , \ADD01/ADD02/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD01/ADD02/u12  (\ADD01/ADD02/n3 , \ADD01/ADD02/p1 , \ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD01/ADD02/u13  (\ADD01/ADD02/n4 , \ADD01/ADD02/n3 , \ADD01/ctemp );  // ../RTL/core/fpu_utils.v(64)
  or \ADD01/ADD02/u14  (\ADD01/ADD02/c1 , \ADD01/ADD02/n2 , \ADD01/ADD02/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD01/ADD02/u15  (\ADD01/ADD02/n5 , \ADD01/ADD02/p2 , \ADD01/ADD02/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD01/ADD02/u16  (\ADD01/ADD02/n6 , \ADD01/ADD02/g2 , \ADD01/ADD02/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD02/u17  (\ADD01/ADD02/n7 , \ADD01/ADD02/p2 , \ADD01/ADD02/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD02/u18  (\ADD01/ADD02/n8 , \ADD01/ADD02/n7 , \ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD01/ADD02/u19  (\ADD01/ADD02/n9 , \ADD01/ADD02/n6 , \ADD01/ADD02/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD02/u2  (\ADD01/ADD02/g2 , n1[29], complemented_E2[6]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD01/ADD02/u20  (temp_exp_diff[7], \ADD01/ADD02/p3 , \ADD01/ADD02/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD01/ADD02/u21  (\ADD01/ADD02/n10 , \ADD01/ADD02/n7 , \ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD02/u22  (\ADD01/ADD02/n11 , \ADD01/ADD02/n10 , \ADD01/ctemp );  // ../RTL/core/fpu_utils.v(65)
  or \ADD01/ADD02/u23  (\ADD01/ADD02/c2 , \ADD01/ADD02/n9 , \ADD01/ADD02/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD02/u24  (\ADD01/ADD02/n12 , \ADD01/ADD02/p3 , \ADD01/ADD02/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD02/u25  (\ADD01/ADD02/n13 , \ADD01/ADD02/g3 , \ADD01/ADD02/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD02/u26  (\ADD01/ADD02/n14 , \ADD01/ADD02/p3 , \ADD01/ADD02/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD02/u27  (\ADD01/ADD02/n15 , \ADD01/ADD02/n14 , \ADD01/ADD02/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD02/u28  (\ADD01/ADD02/n16 , \ADD01/ADD02/n13 , \ADD01/ADD02/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD01/ADD02/u29  (temp_exp_diff[6], \ADD01/ADD02/p2 , \ADD01/ADD02/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD01/ADD02/u3  (\ADD01/ADD02/g3 , n1[30], complemented_E2[7]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD01/ADD02/u30  (\ADD01/ADD02/n17 , \ADD01/ADD02/n14 , \ADD01/ADD02/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD02/u31  (\ADD01/ADD02/n18 , \ADD01/ADD02/n17 , \ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD02/u32  (\ADD01/ADD02/n19 , \ADD01/ADD02/n16 , \ADD01/ADD02/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD01/ADD02/u33  (temp_exp_diff[5], \ADD01/ADD02/p1 , \ADD01/ADD02/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD01/ADD02/u34  (temp_exp_diff[4], \ADD01/ADD02/p0 , \ADD01/ctemp );  // ../RTL/core/fpu_utils.v(71)
  and \ADD01/ADD02/u35  (\ADD01/ADD02/n20 , \ADD01/ADD02/n17 , \ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD02/u36  (\ADD01/ADD02/n21 , \ADD01/ADD02/n20 , \ADD01/ctemp );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD02/u37  (isE1GreaterThanE2, \ADD01/ADD02/n19 , \ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD01/ADD02/u4  (\ADD01/ADD02/p0 , n1[27], complemented_E2[4]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD01/ADD02/u5  (\ADD01/ADD02/p1 , n1[28], complemented_E2[5]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD01/ADD02/u6  (\ADD01/ADD02/p2 , n1[29], complemented_E2[6]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD01/ADD02/u7  (\ADD01/ADD02/p3 , n1[30], complemented_E2[7]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD01/ADD02/u8  (\ADD01/ADD02/n0 , \ADD01/ADD02/p0 , \ADD01/ctemp );  // ../RTL/core/fpu_utils.v(63)
  or \ADD01/ADD02/u9  (\ADD01/ADD02/c0 , \ADD01/ADD02/g0 , \ADD01/ADD02/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD02/ADD01/ADD01/u0  (\ADD02/ADD01/ADD01/g0 , M1[0], new_M2[0]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD02/ADD01/ADD01/u1  (\ADD02/ADD01/ADD01/g1 , M1[1], new_M2[1]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD02/ADD01/ADD01/u10  (\ADD02/ADD01/ADD01/n1 , \ADD02/ADD01/ADD01/p1 , \ADD02/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD01/ADD01/u11  (\ADD02/ADD01/ADD01/n2 , \ADD02/ADD01/ADD01/g1 , \ADD02/ADD01/ADD01/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD01/ADD01/u12  (\ADD02/ADD01/ADD01/n3 , \ADD02/ADD01/ADD01/p1 , \ADD02/ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD01/ADD01/u13  (\ADD02/ADD01/ADD01/n4 , \ADD02/ADD01/ADD01/n3 , real_oper);  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD01/ADD01/u14  (\ADD02/ADD01/ADD01/c1 , \ADD02/ADD01/ADD01/n2 , \ADD02/ADD01/ADD01/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD01/ADD01/u15  (\ADD02/ADD01/ADD01/n5 , \ADD02/ADD01/ADD01/p2 , \ADD02/ADD01/ADD01/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD01/ADD01/u16  (\ADD02/ADD01/ADD01/n6 , \ADD02/ADD01/ADD01/g2 , \ADD02/ADD01/ADD01/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD01/u17  (\ADD02/ADD01/ADD01/n7 , \ADD02/ADD01/ADD01/p2 , \ADD02/ADD01/ADD01/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD01/u18  (\ADD02/ADD01/ADD01/n8 , \ADD02/ADD01/ADD01/n7 , \ADD02/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD01/ADD01/u19  (\ADD02/ADD01/ADD01/n9 , \ADD02/ADD01/ADD01/n6 , \ADD02/ADD01/ADD01/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD01/u2  (\ADD02/ADD01/ADD01/g2 , M1[2], new_M2[2]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD02/ADD01/ADD01/u20  (M_result[3], \ADD02/ADD01/ADD01/p3 , \ADD02/ADD01/ADD01/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD01/ADD01/u21  (\ADD02/ADD01/ADD01/n10 , \ADD02/ADD01/ADD01/n7 , \ADD02/ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD01/u22  (\ADD02/ADD01/ADD01/n11 , \ADD02/ADD01/ADD01/n10 , real_oper);  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD01/ADD01/u23  (\ADD02/ADD01/ADD01/c2 , \ADD02/ADD01/ADD01/n9 , \ADD02/ADD01/ADD01/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD01/u24  (\ADD02/ADD01/ADD01/n12 , \ADD02/ADD01/ADD01/p3 , \ADD02/ADD01/ADD01/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD01/u25  (\ADD02/ADD01/ADD01/n13 , \ADD02/ADD01/ADD01/g3 , \ADD02/ADD01/ADD01/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD01/u26  (\ADD02/ADD01/ADD01/n14 , \ADD02/ADD01/ADD01/p3 , \ADD02/ADD01/ADD01/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD01/u27  (\ADD02/ADD01/ADD01/n15 , \ADD02/ADD01/ADD01/n14 , \ADD02/ADD01/ADD01/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD01/u28  (\ADD02/ADD01/ADD01/n16 , \ADD02/ADD01/ADD01/n13 , \ADD02/ADD01/ADD01/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD01/ADD01/u29  (M_result[2], \ADD02/ADD01/ADD01/p2 , \ADD02/ADD01/ADD01/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD01/ADD01/u3  (\ADD02/ADD01/ADD01/g3 , M1[3], new_M2[3]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD02/ADD01/ADD01/u30  (\ADD02/ADD01/ADD01/n17 , \ADD02/ADD01/ADD01/n14 , \ADD02/ADD01/ADD01/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD01/u31  (\ADD02/ADD01/ADD01/n18 , \ADD02/ADD01/ADD01/n17 , \ADD02/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD01/u32  (\ADD02/ADD01/ADD01/n19 , \ADD02/ADD01/ADD01/n16 , \ADD02/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD01/ADD01/u33  (M_result[1], \ADD02/ADD01/ADD01/p1 , \ADD02/ADD01/ADD01/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD02/ADD01/ADD01/u34  (M_result[0], \ADD02/ADD01/ADD01/p0 , real_oper);  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD01/ADD01/u35  (\ADD02/ADD01/ADD01/n20 , \ADD02/ADD01/ADD01/n17 , \ADD02/ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD01/u36  (\ADD02/ADD01/ADD01/n21 , \ADD02/ADD01/ADD01/n20 , real_oper);  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD01/u37  (\ADD02/ADD01/ctemp , \ADD02/ADD01/ADD01/n19 , \ADD02/ADD01/ADD01/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD01/ADD01/u4  (\ADD02/ADD01/ADD01/p0 , M1[0], new_M2[0]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD02/ADD01/ADD01/u5  (\ADD02/ADD01/ADD01/p1 , M1[1], new_M2[1]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD02/ADD01/ADD01/u6  (\ADD02/ADD01/ADD01/p2 , M1[2], new_M2[2]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD02/ADD01/ADD01/u7  (\ADD02/ADD01/ADD01/p3 , M1[3], new_M2[3]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD02/ADD01/ADD01/u8  (\ADD02/ADD01/ADD01/n0 , \ADD02/ADD01/ADD01/p0 , real_oper);  // ../RTL/core/fpu_utils.v(63)
  or \ADD02/ADD01/ADD01/u9  (\ADD02/ADD01/ADD01/c0 , \ADD02/ADD01/ADD01/g0 , \ADD02/ADD01/ADD01/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD02/ADD01/ADD02/u0  (\ADD02/ADD01/ADD02/g0 , M1[4], new_M2[4]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD02/ADD01/ADD02/u1  (\ADD02/ADD01/ADD02/g1 , M1[5], new_M2[5]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD02/ADD01/ADD02/u10  (\ADD02/ADD01/ADD02/n1 , \ADD02/ADD01/ADD02/p1 , \ADD02/ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD01/ADD02/u11  (\ADD02/ADD01/ADD02/n2 , \ADD02/ADD01/ADD02/g1 , \ADD02/ADD01/ADD02/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD01/ADD02/u12  (\ADD02/ADD01/ADD02/n3 , \ADD02/ADD01/ADD02/p1 , \ADD02/ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD01/ADD02/u13  (\ADD02/ADD01/ADD02/n4 , \ADD02/ADD01/ADD02/n3 , \ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD01/ADD02/u14  (\ADD02/ADD01/ADD02/c1 , \ADD02/ADD01/ADD02/n2 , \ADD02/ADD01/ADD02/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD01/ADD02/u15  (\ADD02/ADD01/ADD02/n5 , \ADD02/ADD01/ADD02/p2 , \ADD02/ADD01/ADD02/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD01/ADD02/u16  (\ADD02/ADD01/ADD02/n6 , \ADD02/ADD01/ADD02/g2 , \ADD02/ADD01/ADD02/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD02/u17  (\ADD02/ADD01/ADD02/n7 , \ADD02/ADD01/ADD02/p2 , \ADD02/ADD01/ADD02/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD02/u18  (\ADD02/ADD01/ADD02/n8 , \ADD02/ADD01/ADD02/n7 , \ADD02/ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD01/ADD02/u19  (\ADD02/ADD01/ADD02/n9 , \ADD02/ADD01/ADD02/n6 , \ADD02/ADD01/ADD02/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD02/u2  (\ADD02/ADD01/ADD02/g2 , M1[6], new_M2[6]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD02/ADD01/ADD02/u20  (M_result[7], \ADD02/ADD01/ADD02/p3 , \ADD02/ADD01/ADD02/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD01/ADD02/u21  (\ADD02/ADD01/ADD02/n10 , \ADD02/ADD01/ADD02/n7 , \ADD02/ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD02/u22  (\ADD02/ADD01/ADD02/n11 , \ADD02/ADD01/ADD02/n10 , \ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD01/ADD02/u23  (\ADD02/ADD01/ADD02/c2 , \ADD02/ADD01/ADD02/n9 , \ADD02/ADD01/ADD02/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD02/u24  (\ADD02/ADD01/ADD02/n12 , \ADD02/ADD01/ADD02/p3 , \ADD02/ADD01/ADD02/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD02/u25  (\ADD02/ADD01/ADD02/n13 , \ADD02/ADD01/ADD02/g3 , \ADD02/ADD01/ADD02/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD02/u26  (\ADD02/ADD01/ADD02/n14 , \ADD02/ADD01/ADD02/p3 , \ADD02/ADD01/ADD02/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD02/u27  (\ADD02/ADD01/ADD02/n15 , \ADD02/ADD01/ADD02/n14 , \ADD02/ADD01/ADD02/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD02/u28  (\ADD02/ADD01/ADD02/n16 , \ADD02/ADD01/ADD02/n13 , \ADD02/ADD01/ADD02/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD01/ADD02/u29  (M_result[6], \ADD02/ADD01/ADD02/p2 , \ADD02/ADD01/ADD02/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD01/ADD02/u3  (\ADD02/ADD01/ADD02/g3 , M1[7], new_M2[7]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD02/ADD01/ADD02/u30  (\ADD02/ADD01/ADD02/n17 , \ADD02/ADD01/ADD02/n14 , \ADD02/ADD01/ADD02/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD02/u31  (\ADD02/ADD01/ADD02/n18 , \ADD02/ADD01/ADD02/n17 , \ADD02/ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD02/u32  (\ADD02/ADD01/ADD02/n19 , \ADD02/ADD01/ADD02/n16 , \ADD02/ADD01/ADD02/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD01/ADD02/u33  (M_result[5], \ADD02/ADD01/ADD02/p1 , \ADD02/ADD01/ADD02/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD02/ADD01/ADD02/u34  (M_result[4], \ADD02/ADD01/ADD02/p0 , \ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD01/ADD02/u35  (\ADD02/ADD01/ADD02/n20 , \ADD02/ADD01/ADD02/n17 , \ADD02/ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD02/u36  (\ADD02/ADD01/ADD02/n21 , \ADD02/ADD01/ADD02/n20 , \ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD02/u37  (\ADD02/ctemp1 , \ADD02/ADD01/ADD02/n19 , \ADD02/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD01/ADD02/u4  (\ADD02/ADD01/ADD02/p0 , M1[4], new_M2[4]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD02/ADD01/ADD02/u5  (\ADD02/ADD01/ADD02/p1 , M1[5], new_M2[5]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD02/ADD01/ADD02/u6  (\ADD02/ADD01/ADD02/p2 , M1[6], new_M2[6]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD02/ADD01/ADD02/u7  (\ADD02/ADD01/ADD02/p3 , M1[7], new_M2[7]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD02/ADD01/ADD02/u8  (\ADD02/ADD01/ADD02/n0 , \ADD02/ADD01/ADD02/p0 , \ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(63)
  or \ADD02/ADD01/ADD02/u9  (\ADD02/ADD01/ADD02/c0 , \ADD02/ADD01/ADD02/g0 , \ADD02/ADD01/ADD02/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD02/ADD02/ADD01/u0  (\ADD02/ADD02/ADD01/g0 , M1[8], new_M2[8]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD02/ADD02/ADD01/u1  (\ADD02/ADD02/ADD01/g1 , M1[9], new_M2[9]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD02/ADD02/ADD01/u10  (\ADD02/ADD02/ADD01/n1 , \ADD02/ADD02/ADD01/p1 , \ADD02/ADD02/ADD01/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD02/ADD01/u11  (\ADD02/ADD02/ADD01/n2 , \ADD02/ADD02/ADD01/g1 , \ADD02/ADD02/ADD01/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD02/ADD01/u12  (\ADD02/ADD02/ADD01/n3 , \ADD02/ADD02/ADD01/p1 , \ADD02/ADD02/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD02/ADD01/u13  (\ADD02/ADD02/ADD01/n4 , \ADD02/ADD02/ADD01/n3 , \ADD02/ctemp1 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD02/ADD01/u14  (\ADD02/ADD02/ADD01/c1 , \ADD02/ADD02/ADD01/n2 , \ADD02/ADD02/ADD01/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD02/ADD01/u15  (\ADD02/ADD02/ADD01/n5 , \ADD02/ADD02/ADD01/p2 , \ADD02/ADD02/ADD01/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD02/ADD01/u16  (\ADD02/ADD02/ADD01/n6 , \ADD02/ADD02/ADD01/g2 , \ADD02/ADD02/ADD01/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD01/u17  (\ADD02/ADD02/ADD01/n7 , \ADD02/ADD02/ADD01/p2 , \ADD02/ADD02/ADD01/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD01/u18  (\ADD02/ADD02/ADD01/n8 , \ADD02/ADD02/ADD01/n7 , \ADD02/ADD02/ADD01/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD02/ADD01/u19  (\ADD02/ADD02/ADD01/n9 , \ADD02/ADD02/ADD01/n6 , \ADD02/ADD02/ADD01/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD01/u2  (\ADD02/ADD02/ADD01/g2 , M1[10], new_M2[10]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD02/ADD02/ADD01/u20  (M_result[11], \ADD02/ADD02/ADD01/p3 , \ADD02/ADD02/ADD01/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD02/ADD01/u21  (\ADD02/ADD02/ADD01/n10 , \ADD02/ADD02/ADD01/n7 , \ADD02/ADD02/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD01/u22  (\ADD02/ADD02/ADD01/n11 , \ADD02/ADD02/ADD01/n10 , \ADD02/ctemp1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD02/ADD01/u23  (\ADD02/ADD02/ADD01/c2 , \ADD02/ADD02/ADD01/n9 , \ADD02/ADD02/ADD01/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD01/u24  (\ADD02/ADD02/ADD01/n12 , \ADD02/ADD02/ADD01/p3 , \ADD02/ADD02/ADD01/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD01/u25  (\ADD02/ADD02/ADD01/n13 , \ADD02/ADD02/ADD01/g3 , \ADD02/ADD02/ADD01/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD01/u26  (\ADD02/ADD02/ADD01/n14 , \ADD02/ADD02/ADD01/p3 , \ADD02/ADD02/ADD01/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD01/u27  (\ADD02/ADD02/ADD01/n15 , \ADD02/ADD02/ADD01/n14 , \ADD02/ADD02/ADD01/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD01/u28  (\ADD02/ADD02/ADD01/n16 , \ADD02/ADD02/ADD01/n13 , \ADD02/ADD02/ADD01/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD02/ADD01/u29  (M_result[10], \ADD02/ADD02/ADD01/p2 , \ADD02/ADD02/ADD01/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD02/ADD01/u3  (\ADD02/ADD02/ADD01/g3 , M1[11], new_M2[11]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD02/ADD02/ADD01/u30  (\ADD02/ADD02/ADD01/n17 , \ADD02/ADD02/ADD01/n14 , \ADD02/ADD02/ADD01/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD01/u31  (\ADD02/ADD02/ADD01/n18 , \ADD02/ADD02/ADD01/n17 , \ADD02/ADD02/ADD01/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD01/u32  (\ADD02/ADD02/ADD01/n19 , \ADD02/ADD02/ADD01/n16 , \ADD02/ADD02/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD02/ADD01/u33  (M_result[9], \ADD02/ADD02/ADD01/p1 , \ADD02/ADD02/ADD01/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD02/ADD02/ADD01/u34  (M_result[8], \ADD02/ADD02/ADD01/p0 , \ADD02/ctemp1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD02/ADD01/u35  (\ADD02/ADD02/ADD01/n20 , \ADD02/ADD02/ADD01/n17 , \ADD02/ADD02/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD01/u36  (\ADD02/ADD02/ADD01/n21 , \ADD02/ADD02/ADD01/n20 , \ADD02/ctemp1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD01/u37  (\ADD02/ADD02/ctemp , \ADD02/ADD02/ADD01/n19 , \ADD02/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD02/ADD01/u4  (\ADD02/ADD02/ADD01/p0 , M1[8], new_M2[8]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD02/ADD02/ADD01/u5  (\ADD02/ADD02/ADD01/p1 , M1[9], new_M2[9]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD02/ADD02/ADD01/u6  (\ADD02/ADD02/ADD01/p2 , M1[10], new_M2[10]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD02/ADD02/ADD01/u7  (\ADD02/ADD02/ADD01/p3 , M1[11], new_M2[11]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD02/ADD02/ADD01/u8  (\ADD02/ADD02/ADD01/n0 , \ADD02/ADD02/ADD01/p0 , \ADD02/ctemp1 );  // ../RTL/core/fpu_utils.v(63)
  or \ADD02/ADD02/ADD01/u9  (\ADD02/ADD02/ADD01/c0 , \ADD02/ADD02/ADD01/g0 , \ADD02/ADD02/ADD01/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD02/ADD02/ADD02/u0  (\ADD02/ADD02/ADD02/g0 , M1[12], new_M2[12]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD02/ADD02/ADD02/u1  (\ADD02/ADD02/ADD02/g1 , M1[13], new_M2[13]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD02/ADD02/ADD02/u10  (\ADD02/ADD02/ADD02/n1 , \ADD02/ADD02/ADD02/p1 , \ADD02/ADD02/ADD02/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD02/ADD02/u11  (\ADD02/ADD02/ADD02/n2 , \ADD02/ADD02/ADD02/g1 , \ADD02/ADD02/ADD02/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD02/ADD02/u12  (\ADD02/ADD02/ADD02/n3 , \ADD02/ADD02/ADD02/p1 , \ADD02/ADD02/ADD02/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD02/ADD02/u13  (\ADD02/ADD02/ADD02/n4 , \ADD02/ADD02/ADD02/n3 , \ADD02/ADD02/ctemp );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD02/ADD02/u14  (\ADD02/ADD02/ADD02/c1 , \ADD02/ADD02/ADD02/n2 , \ADD02/ADD02/ADD02/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD02/ADD02/u15  (\ADD02/ADD02/ADD02/n5 , \ADD02/ADD02/ADD02/p2 , \ADD02/ADD02/ADD02/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD02/ADD02/u16  (\ADD02/ADD02/ADD02/n6 , \ADD02/ADD02/ADD02/g2 , \ADD02/ADD02/ADD02/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD02/u17  (\ADD02/ADD02/ADD02/n7 , \ADD02/ADD02/ADD02/p2 , \ADD02/ADD02/ADD02/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD02/u18  (\ADD02/ADD02/ADD02/n8 , \ADD02/ADD02/ADD02/n7 , \ADD02/ADD02/ADD02/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD02/ADD02/u19  (\ADD02/ADD02/ADD02/n9 , \ADD02/ADD02/ADD02/n6 , \ADD02/ADD02/ADD02/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD02/u2  (\ADD02/ADD02/ADD02/g2 , M1[14], new_M2[14]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD02/ADD02/ADD02/u20  (M_result[15], \ADD02/ADD02/ADD02/p3 , \ADD02/ADD02/ADD02/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD02/ADD02/u21  (\ADD02/ADD02/ADD02/n10 , \ADD02/ADD02/ADD02/n7 , \ADD02/ADD02/ADD02/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD02/u22  (\ADD02/ADD02/ADD02/n11 , \ADD02/ADD02/ADD02/n10 , \ADD02/ADD02/ctemp );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD02/ADD02/u23  (\ADD02/ADD02/ADD02/c2 , \ADD02/ADD02/ADD02/n9 , \ADD02/ADD02/ADD02/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD02/u24  (\ADD02/ADD02/ADD02/n12 , \ADD02/ADD02/ADD02/p3 , \ADD02/ADD02/ADD02/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD02/u25  (\ADD02/ADD02/ADD02/n13 , \ADD02/ADD02/ADD02/g3 , \ADD02/ADD02/ADD02/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD02/u26  (\ADD02/ADD02/ADD02/n14 , \ADD02/ADD02/ADD02/p3 , \ADD02/ADD02/ADD02/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD02/u27  (\ADD02/ADD02/ADD02/n15 , \ADD02/ADD02/ADD02/n14 , \ADD02/ADD02/ADD02/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD02/u28  (\ADD02/ADD02/ADD02/n16 , \ADD02/ADD02/ADD02/n13 , \ADD02/ADD02/ADD02/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD02/ADD02/u29  (M_result[14], \ADD02/ADD02/ADD02/p2 , \ADD02/ADD02/ADD02/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD02/ADD02/u3  (\ADD02/ADD02/ADD02/g3 , M1[15], new_M2[15]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD02/ADD02/ADD02/u30  (\ADD02/ADD02/ADD02/n17 , \ADD02/ADD02/ADD02/n14 , \ADD02/ADD02/ADD02/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD02/u31  (\ADD02/ADD02/ADD02/n18 , \ADD02/ADD02/ADD02/n17 , \ADD02/ADD02/ADD02/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD02/u32  (\ADD02/ADD02/ADD02/n19 , \ADD02/ADD02/ADD02/n16 , \ADD02/ADD02/ADD02/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD02/ADD02/u33  (M_result[13], \ADD02/ADD02/ADD02/p1 , \ADD02/ADD02/ADD02/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD02/ADD02/ADD02/u34  (M_result[12], \ADD02/ADD02/ADD02/p0 , \ADD02/ADD02/ctemp );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD02/ADD02/u35  (\ADD02/ADD02/ADD02/n20 , \ADD02/ADD02/ADD02/n17 , \ADD02/ADD02/ADD02/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD02/u36  (\ADD02/ADD02/ADD02/n21 , \ADD02/ADD02/ADD02/n20 , \ADD02/ADD02/ctemp );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD02/u37  (\ADD02/ctemp2 , \ADD02/ADD02/ADD02/n19 , \ADD02/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD02/ADD02/u4  (\ADD02/ADD02/ADD02/p0 , M1[12], new_M2[12]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD02/ADD02/ADD02/u5  (\ADD02/ADD02/ADD02/p1 , M1[13], new_M2[13]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD02/ADD02/ADD02/u6  (\ADD02/ADD02/ADD02/p2 , M1[14], new_M2[14]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD02/ADD02/ADD02/u7  (\ADD02/ADD02/ADD02/p3 , M1[15], new_M2[15]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD02/ADD02/ADD02/u8  (\ADD02/ADD02/ADD02/n0 , \ADD02/ADD02/ADD02/p0 , \ADD02/ADD02/ctemp );  // ../RTL/core/fpu_utils.v(63)
  or \ADD02/ADD02/ADD02/u9  (\ADD02/ADD02/ADD02/c0 , \ADD02/ADD02/ADD02/g0 , \ADD02/ADD02/ADD02/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD02/ADD03/ADD01/u0  (\ADD02/ADD03/ADD01/g0 , M1[16], new_M2[16]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD02/ADD03/ADD01/u1  (\ADD02/ADD03/ADD01/g1 , M1[17], new_M2[17]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD02/ADD03/ADD01/u10  (\ADD02/ADD03/ADD01/n1 , \ADD02/ADD03/ADD01/p1 , \ADD02/ADD03/ADD01/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD03/ADD01/u11  (\ADD02/ADD03/ADD01/n2 , \ADD02/ADD03/ADD01/g1 , \ADD02/ADD03/ADD01/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD03/ADD01/u12  (\ADD02/ADD03/ADD01/n3 , \ADD02/ADD03/ADD01/p1 , \ADD02/ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD03/ADD01/u13  (\ADD02/ADD03/ADD01/n4 , \ADD02/ADD03/ADD01/n3 , \ADD02/ctemp2 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD03/ADD01/u14  (\ADD02/ADD03/ADD01/c1 , \ADD02/ADD03/ADD01/n2 , \ADD02/ADD03/ADD01/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD03/ADD01/u15  (\ADD02/ADD03/ADD01/n5 , \ADD02/ADD03/ADD01/p2 , \ADD02/ADD03/ADD01/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD03/ADD01/u16  (\ADD02/ADD03/ADD01/n6 , \ADD02/ADD03/ADD01/g2 , \ADD02/ADD03/ADD01/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD01/u17  (\ADD02/ADD03/ADD01/n7 , \ADD02/ADD03/ADD01/p2 , \ADD02/ADD03/ADD01/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD01/u18  (\ADD02/ADD03/ADD01/n8 , \ADD02/ADD03/ADD01/n7 , \ADD02/ADD03/ADD01/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD03/ADD01/u19  (\ADD02/ADD03/ADD01/n9 , \ADD02/ADD03/ADD01/n6 , \ADD02/ADD03/ADD01/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD01/u2  (\ADD02/ADD03/ADD01/g2 , M1[18], new_M2[18]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD02/ADD03/ADD01/u20  (M_result[19], \ADD02/ADD03/ADD01/p3 , \ADD02/ADD03/ADD01/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD03/ADD01/u21  (\ADD02/ADD03/ADD01/n10 , \ADD02/ADD03/ADD01/n7 , \ADD02/ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD01/u22  (\ADD02/ADD03/ADD01/n11 , \ADD02/ADD03/ADD01/n10 , \ADD02/ctemp2 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD03/ADD01/u23  (\ADD02/ADD03/ADD01/c2 , \ADD02/ADD03/ADD01/n9 , \ADD02/ADD03/ADD01/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD01/u24  (\ADD02/ADD03/ADD01/n12 , \ADD02/ADD03/ADD01/p3 , \ADD02/ADD03/ADD01/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD01/u25  (\ADD02/ADD03/ADD01/n13 , \ADD02/ADD03/ADD01/g3 , \ADD02/ADD03/ADD01/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD01/u26  (\ADD02/ADD03/ADD01/n14 , \ADD02/ADD03/ADD01/p3 , \ADD02/ADD03/ADD01/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD01/u27  (\ADD02/ADD03/ADD01/n15 , \ADD02/ADD03/ADD01/n14 , \ADD02/ADD03/ADD01/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD01/u28  (\ADD02/ADD03/ADD01/n16 , \ADD02/ADD03/ADD01/n13 , \ADD02/ADD03/ADD01/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD03/ADD01/u29  (M_result[18], \ADD02/ADD03/ADD01/p2 , \ADD02/ADD03/ADD01/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD03/ADD01/u3  (\ADD02/ADD03/ADD01/g3 , M1[19], new_M2[19]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD02/ADD03/ADD01/u30  (\ADD02/ADD03/ADD01/n17 , \ADD02/ADD03/ADD01/n14 , \ADD02/ADD03/ADD01/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD01/u31  (\ADD02/ADD03/ADD01/n18 , \ADD02/ADD03/ADD01/n17 , \ADD02/ADD03/ADD01/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD01/u32  (\ADD02/ADD03/ADD01/n19 , \ADD02/ADD03/ADD01/n16 , \ADD02/ADD03/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD03/ADD01/u33  (M_result[17], \ADD02/ADD03/ADD01/p1 , \ADD02/ADD03/ADD01/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD02/ADD03/ADD01/u34  (M_result[16], \ADD02/ADD03/ADD01/p0 , \ADD02/ctemp2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD03/ADD01/u35  (\ADD02/ADD03/ADD01/n20 , \ADD02/ADD03/ADD01/n17 , \ADD02/ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD01/u36  (\ADD02/ADD03/ADD01/n21 , \ADD02/ADD03/ADD01/n20 , \ADD02/ctemp2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD01/u37  (\ADD02/ADD03/ctemp , \ADD02/ADD03/ADD01/n19 , \ADD02/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD03/ADD01/u4  (\ADD02/ADD03/ADD01/p0 , M1[16], new_M2[16]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD02/ADD03/ADD01/u5  (\ADD02/ADD03/ADD01/p1 , M1[17], new_M2[17]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD02/ADD03/ADD01/u6  (\ADD02/ADD03/ADD01/p2 , M1[18], new_M2[18]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD02/ADD03/ADD01/u7  (\ADD02/ADD03/ADD01/p3 , M1[19], new_M2[19]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD02/ADD03/ADD01/u8  (\ADD02/ADD03/ADD01/n0 , \ADD02/ADD03/ADD01/p0 , \ADD02/ctemp2 );  // ../RTL/core/fpu_utils.v(63)
  or \ADD02/ADD03/ADD01/u9  (\ADD02/ADD03/ADD01/c0 , \ADD02/ADD03/ADD01/g0 , \ADD02/ADD03/ADD01/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD02/ADD03/ADD02/u0  (\ADD02/ADD03/ADD02/g0 , M1[20], new_M2[20]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD02/ADD03/ADD02/u1  (\ADD02/ADD03/ADD02/g1 , M1[21], new_M2[21]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD02/ADD03/ADD02/u10  (\ADD02/ADD03/ADD02/n1 , \ADD02/ADD03/ADD02/p1 , \ADD02/ADD03/ADD02/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD03/ADD02/u11  (\ADD02/ADD03/ADD02/n2 , \ADD02/ADD03/ADD02/g1 , \ADD02/ADD03/ADD02/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD03/ADD02/u12  (\ADD02/ADD03/ADD02/n3 , \ADD02/ADD03/ADD02/p1 , \ADD02/ADD03/ADD02/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD03/ADD02/u13  (\ADD02/ADD03/ADD02/n4 , \ADD02/ADD03/ADD02/n3 , \ADD02/ADD03/ctemp );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD03/ADD02/u14  (\ADD02/ADD03/ADD02/c1 , \ADD02/ADD03/ADD02/n2 , \ADD02/ADD03/ADD02/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD03/ADD02/u15  (\ADD02/ADD03/ADD02/n5 , \ADD02/ADD03/ADD02/p2 , \ADD02/ADD03/ADD02/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD03/ADD02/u16  (\ADD02/ADD03/ADD02/n6 , \ADD02/ADD03/ADD02/g2 , \ADD02/ADD03/ADD02/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD02/u17  (\ADD02/ADD03/ADD02/n7 , \ADD02/ADD03/ADD02/p2 , \ADD02/ADD03/ADD02/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD02/u18  (\ADD02/ADD03/ADD02/n8 , \ADD02/ADD03/ADD02/n7 , \ADD02/ADD03/ADD02/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD03/ADD02/u19  (\ADD02/ADD03/ADD02/n9 , \ADD02/ADD03/ADD02/n6 , \ADD02/ADD03/ADD02/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD02/u2  (\ADD02/ADD03/ADD02/g2 , M1[22], new_M2[22]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD02/ADD03/ADD02/u20  (M_result[23], \ADD02/ADD03/ADD02/p3 , \ADD02/ADD03/ADD02/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD03/ADD02/u21  (\ADD02/ADD03/ADD02/n10 , \ADD02/ADD03/ADD02/n7 , \ADD02/ADD03/ADD02/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD02/u22  (\ADD02/ADD03/ADD02/n11 , \ADD02/ADD03/ADD02/n10 , \ADD02/ADD03/ctemp );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD03/ADD02/u23  (\ADD02/ADD03/ADD02/c2 , \ADD02/ADD03/ADD02/n9 , \ADD02/ADD03/ADD02/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD02/u24  (\ADD02/ADD03/ADD02/n12 , \ADD02/ADD03/ADD02/p3 , \ADD02/ADD03/ADD02/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD02/u25  (\ADD02/ADD03/ADD02/n13 , \ADD02/ADD03/ADD02/g3 , \ADD02/ADD03/ADD02/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD02/u26  (\ADD02/ADD03/ADD02/n14 , \ADD02/ADD03/ADD02/p3 , \ADD02/ADD03/ADD02/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD02/u27  (\ADD02/ADD03/ADD02/n15 , \ADD02/ADD03/ADD02/n14 , \ADD02/ADD03/ADD02/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD02/u28  (\ADD02/ADD03/ADD02/n16 , \ADD02/ADD03/ADD02/n13 , \ADD02/ADD03/ADD02/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD03/ADD02/u29  (M_result[22], \ADD02/ADD03/ADD02/p2 , \ADD02/ADD03/ADD02/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD03/ADD02/u3  (\ADD02/ADD03/ADD02/g3 , M1[23], new_M2[23]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD02/ADD03/ADD02/u30  (\ADD02/ADD03/ADD02/n17 , \ADD02/ADD03/ADD02/n14 , \ADD02/ADD03/ADD02/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD02/u31  (\ADD02/ADD03/ADD02/n18 , \ADD02/ADD03/ADD02/n17 , \ADD02/ADD03/ADD02/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD02/u32  (\ADD02/ADD03/ADD02/n19 , \ADD02/ADD03/ADD02/n16 , \ADD02/ADD03/ADD02/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD03/ADD02/u33  (M_result[21], \ADD02/ADD03/ADD02/p1 , \ADD02/ADD03/ADD02/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD02/ADD03/ADD02/u34  (M_result[20], \ADD02/ADD03/ADD02/p0 , \ADD02/ADD03/ctemp );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD03/ADD02/u35  (\ADD02/ADD03/ADD02/n20 , \ADD02/ADD03/ADD02/n17 , \ADD02/ADD03/ADD02/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD02/u36  (\ADD02/ADD03/ADD02/n21 , \ADD02/ADD03/ADD02/n20 , \ADD02/ADD03/ctemp );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD02/u37  (M_carry, \ADD02/ADD03/ADD02/n19 , \ADD02/ADD03/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD03/ADD02/u4  (\ADD02/ADD03/ADD02/p0 , M1[20], new_M2[20]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD02/ADD03/ADD02/u5  (\ADD02/ADD03/ADD02/p1 , M1[21], new_M2[21]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD02/ADD03/ADD02/u6  (\ADD02/ADD03/ADD02/p2 , M1[22], new_M2[22]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD02/ADD03/ADD02/u7  (\ADD02/ADD03/ADD02/p3 , M1[23], new_M2[23]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD02/ADD03/ADD02/u8  (\ADD02/ADD03/ADD02/n0 , \ADD02/ADD03/ADD02/p0 , \ADD02/ADD03/ctemp );  // ../RTL/core/fpu_utils.v(63)
  or \ADD02/ADD03/ADD02/u9  (\ADD02/ADD03/ADD02/c0 , \ADD02/ADD03/ADD02/g0 , \ADD02/ADD03/ADD02/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD0212/ADD01/u10  (\ADD0212/ADD01/n1 , E[1], E[0]);  // ../RTL/core/fpu_utils.v(64)
  and \ADD0212/ADD01/u17  (\ADD0212/ADD01/n7 , E[2], E[1]);  // ../RTL/core/fpu_utils.v(65)
  and \ADD0212/ADD01/u18  (\ADD0212/ADD01/n8 , \ADD0212/ADD01/n7 , E[0]);  // ../RTL/core/fpu_utils.v(65)
  xor \ADD0212/ADD01/u20  (One_Added_E[3], E[3], \ADD0212/ADD01/n8 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD0212/ADD01/u26  (\ADD0212/ADD01/n14 , E[3], E[2]);  // ../RTL/core/fpu_utils.v(66)
  xor \ADD0212/ADD01/u29  (One_Added_E[2], E[2], \ADD0212/ADD01/n1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD0212/ADD01/u30  (\ADD0212/ADD01/n17 , \ADD0212/ADD01/n14 , E[1]);  // ../RTL/core/fpu_utils.v(66)
  and \ADD0212/ADD01/u31  (\ADD0212/ADD01/n18 , \ADD0212/ADD01/n17 , E[0]);  // ../RTL/core/fpu_utils.v(66)
  xor \ADD0212/ADD01/u33  (One_Added_E[1], E[1], E[0]);  // ../RTL/core/fpu_utils.v(71)
  and \ADD0212/ADD02/u12  (\ADD0212/ADD02/n3 , E[5], E[4]);  // ../RTL/core/fpu_utils.v(64)
  and \ADD0212/ADD02/u13  (\ADD0212/ADD02/n4 , \ADD0212/ADD02/n3 , \ADD0212/ADD01/n18 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD0212/ADD02/u17  (\ADD0212/ADD02/n7 , E[6], E[5]);  // ../RTL/core/fpu_utils.v(65)
  xor \ADD0212/ADD02/u20  (One_Added_E[7], E[7], \ADD0212/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD0212/ADD02/u21  (\ADD0212/ADD02/n10 , \ADD0212/ADD02/n7 , E[4]);  // ../RTL/core/fpu_utils.v(65)
  and \ADD0212/ADD02/u22  (\ADD0212/ADD02/n11 , \ADD0212/ADD02/n10 , \ADD0212/ADD01/n18 );  // ../RTL/core/fpu_utils.v(65)
  xor \ADD0212/ADD02/u29  (One_Added_E[6], E[6], \ADD0212/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD0212/ADD02/u33  (One_Added_E[5], E[5], \ADD0212/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD0212/ADD02/u34  (One_Added_E[4], E[4], \ADD0212/ADD01/n18 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD0212/ADD02/u8  (\ADD0212/ADD02/n0 , E[4], \ADD0212/ADD01/n18 );  // ../RTL/core/fpu_utils.v(63)
  not \ADD03/ADD01/p0_inv  (\ADD03/ADD01/p0_neg , \ADD03/ADD01/p0 );
  and \ADD03/ADD01/u0  (\ADD03/ADD01/g0 , new_E[0], complemented_shift_E[0]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD03/ADD01/u1  (\ADD03/ADD01/g1 , new_E[1], complemented_shift_E[1]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD03/ADD01/u10  (\ADD03/ADD01/n1 , \ADD03/ADD01/p1 , \ADD03/ADD01/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD03/ADD01/u11  (\ADD03/ADD01/n2 , \ADD03/ADD01/g1 , \ADD03/ADD01/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD03/ADD01/u12  (\ADD03/ADD01/n3 , \ADD03/ADD01/p1 , \ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD03/ADD01/u14  (\ADD03/ADD01/c1 , \ADD03/ADD01/n2 , \ADD03/ADD01/n3 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD03/ADD01/u15  (\ADD03/ADD01/n5 , \ADD03/ADD01/p2 , \ADD03/ADD01/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD03/ADD01/u16  (\ADD03/ADD01/n6 , \ADD03/ADD01/g2 , \ADD03/ADD01/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD01/u17  (\ADD03/ADD01/n7 , \ADD03/ADD01/p2 , \ADD03/ADD01/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD01/u18  (\ADD03/ADD01/n8 , \ADD03/ADD01/n7 , \ADD03/ADD01/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD03/ADD01/u19  (\ADD03/ADD01/n9 , \ADD03/ADD01/n6 , \ADD03/ADD01/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD01/u2  (\ADD03/ADD01/g2 , new_E[2], complemented_shift_E[2]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD03/ADD01/u20  (result[26], \ADD03/ADD01/p3 , \ADD03/ADD01/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD03/ADD01/u21  (\ADD03/ADD01/n10 , \ADD03/ADD01/n7 , \ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD03/ADD01/u23  (\ADD03/ADD01/c2 , \ADD03/ADD01/n9 , \ADD03/ADD01/n10 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD01/u24  (\ADD03/ADD01/n12 , \ADD03/ADD01/p3 , \ADD03/ADD01/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD03/ADD01/u25  (\ADD03/ADD01/n13 , \ADD03/ADD01/g3 , \ADD03/ADD01/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD03/ADD01/u26  (\ADD03/ADD01/n14 , \ADD03/ADD01/p3 , \ADD03/ADD01/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD03/ADD01/u27  (\ADD03/ADD01/n15 , \ADD03/ADD01/n14 , \ADD03/ADD01/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD03/ADD01/u28  (\ADD03/ADD01/n16 , \ADD03/ADD01/n13 , \ADD03/ADD01/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD03/ADD01/u29  (result[25], \ADD03/ADD01/p2 , \ADD03/ADD01/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD03/ADD01/u3  (\ADD03/ADD01/g3 , new_E[3], complemented_shift_E[3]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD03/ADD01/u30  (\ADD03/ADD01/n17 , \ADD03/ADD01/n14 , \ADD03/ADD01/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD03/ADD01/u31  (\ADD03/ADD01/n18 , \ADD03/ADD01/n17 , \ADD03/ADD01/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD03/ADD01/u32  (\ADD03/ADD01/n19 , \ADD03/ADD01/n16 , \ADD03/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD03/ADD01/u33  (result[24], \ADD03/ADD01/p1 , \ADD03/ADD01/c0 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD03/ADD01/u35  (\ADD03/ADD01/n20 , \ADD03/ADD01/n17 , \ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD03/ADD01/u37  (\ADD03/ctemp , \ADD03/ADD01/n19 , \ADD03/ADD01/n20 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD03/ADD01/u4  (\ADD03/ADD01/p0 , new_E[0], complemented_shift_E[0]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD03/ADD01/u5  (\ADD03/ADD01/p1 , new_E[1], complemented_shift_E[1]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD03/ADD01/u6  (\ADD03/ADD01/p2 , new_E[2], complemented_shift_E[2]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD03/ADD01/u7  (\ADD03/ADD01/p3 , new_E[3], complemented_shift_E[3]);  // ../RTL/core/fpu_utils.v(62)
  or \ADD03/ADD01/u9  (\ADD03/ADD01/c0 , \ADD03/ADD01/g0 , \ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD03/ADD02/u0  (\ADD03/ADD02/g0 , new_E[4], complemented_shift_E[4]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD03/ADD02/u10  (\ADD03/ADD02/n1 , \new_E[5]_neg , \ADD03/ADD02/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD03/ADD02/u11  (\ADD03/ADD02/n2 , new_E[5], \ADD03/ADD02/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD03/ADD02/u12  (\ADD03/ADD02/n3 , \new_E[5]_neg , \ADD03/ADD02/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD03/ADD02/u13  (\ADD03/ADD02/n4 , \ADD03/ADD02/n3 , \ADD03/ctemp );  // ../RTL/core/fpu_utils.v(64)
  or \ADD03/ADD02/u14  (\ADD03/ADD02/c1 , \ADD03/ADD02/n2 , \ADD03/ADD02/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD03/ADD02/u15  (\ADD03/ADD02/n5 , \new_E[6]_neg , new_E[5]);  // ../RTL/core/fpu_utils.v(65)
  or \ADD03/ADD02/u16  (\ADD03/ADD02/n6 , new_E[6], \ADD03/ADD02/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD02/u17  (\ADD03/ADD02/n7 , \new_E[6]_neg , \new_E[5]_neg );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD02/u18  (\ADD03/ADD02/n8 , \ADD03/ADD02/n7 , \ADD03/ADD02/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD03/ADD02/u19  (\ADD03/ADD02/n9 , \ADD03/ADD02/n6 , \ADD03/ADD02/n8 );  // ../RTL/core/fpu_utils.v(65)
  xor \ADD03/ADD02/u20  (result[30], \new_E[7]_neg , \ADD03/ADD02/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD03/ADD02/u21  (\ADD03/ADD02/n10 , \ADD03/ADD02/n7 , \ADD03/ADD02/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD02/u22  (\ADD03/ADD02/n11 , \ADD03/ADD02/n10 , \ADD03/ctemp );  // ../RTL/core/fpu_utils.v(65)
  or \ADD03/ADD02/u23  (\ADD03/ADD02/c2 , \ADD03/ADD02/n9 , \ADD03/ADD02/n11 );  // ../RTL/core/fpu_utils.v(65)
  xor \ADD03/ADD02/u29  (result[29], \new_E[6]_neg , \ADD03/ADD02/c1 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD03/ADD02/u33  (result[28], \new_E[5]_neg , \ADD03/ADD02/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD03/ADD02/u34  (result[27], \ADD03/ADD02/p0 , \ADD03/ctemp );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD03/ADD02/u4  (\ADD03/ADD02/p0 , new_E[4], complemented_shift_E[4]);  // ../RTL/core/fpu_utils.v(59)
  and \ADD03/ADD02/u8  (\ADD03/ADD02/n0 , \ADD03/ADD02/p0 , \ADD03/ctemp );  // ../RTL/core/fpu_utils.v(63)
  or \ADD03/ADD02/u9  (\ADD03/ADD02/c0 , \ADD03/ADD02/g0 , \ADD03/ADD02/n0 );  // ../RTL/core/fpu_utils.v(63)
  not \C01/u0  (complemented_E2[3], n2[26]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u1  (complemented_E2[2], n2[25]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u2  (complemented_E2[1], n2[24]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u3  (complemented_E2[0], n2[23]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u4  (complemented_E2[7], n2[30]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u5  (complemented_E2[6], n2[29]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u6  (complemented_E2[5], n2[28]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u7  (complemented_E2[4], n2[27]);  // ../RTL/core/fpu_utils.v(44)
  and \C023/ADD01/ADD01/u10  (\C023/ADD01/ADD01/n1 , \C023/outtemp [1], \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \C023/ADD01/ADD01/u17  (\C023/ADD01/ADD01/n7 , \C023/outtemp [2], \C023/outtemp [1]);  // ../RTL/core/fpu_utils.v(65)
  and \C023/ADD01/ADD01/u18  (\C023/ADD01/ADD01/n8 , \C023/ADD01/ADD01/n7 , \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  xor \C023/ADD01/ADD01/u20  (complemented_temp_exp_diff[3], \C023/outtemp [3], \C023/ADD01/ADD01/n8 );  // ../RTL/core/fpu_utils.v(71)
  and \C023/ADD01/ADD01/u26  (\C023/ADD01/ADD01/n14 , \C023/outtemp [3], \C023/outtemp [2]);  // ../RTL/core/fpu_utils.v(66)
  xor \C023/ADD01/ADD01/u29  (complemented_temp_exp_diff[2], \C023/outtemp [2], \C023/ADD01/ADD01/n1 );  // ../RTL/core/fpu_utils.v(71)
  and \C023/ADD01/ADD01/u30  (\C023/ADD01/ADD01/n17 , \C023/ADD01/ADD01/n14 , \C023/outtemp [1]);  // ../RTL/core/fpu_utils.v(66)
  and \C023/ADD01/ADD01/u31  (\C023/ADD01/ADD01/n18 , \C023/ADD01/ADD01/n17 , \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  xor \C023/ADD01/ADD01/u33  (complemented_temp_exp_diff[1], \C023/outtemp [1], \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(71)
  and \C023/ADD01/ADD02/u12  (\C023/ADD01/ADD02/n3 , \C023/outtemp [5], \C023/outtemp [4]);  // ../RTL/core/fpu_utils.v(64)
  and \C023/ADD01/ADD02/u13  (\C023/ADD01/ADD02/n4 , \C023/ADD01/ADD02/n3 , \C023/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(64)
  and \C023/ADD01/ADD02/u17  (\C023/ADD01/ADD02/n7 , \C023/outtemp [6], \C023/outtemp [5]);  // ../RTL/core/fpu_utils.v(65)
  xor \C023/ADD01/ADD02/u20  (complemented_temp_exp_diff[7], \C023/outtemp [7], \C023/ADD01/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \C023/ADD01/ADD02/u21  (\C023/ADD01/ADD02/n10 , \C023/ADD01/ADD02/n7 , \C023/outtemp [4]);  // ../RTL/core/fpu_utils.v(65)
  and \C023/ADD01/ADD02/u22  (\C023/ADD01/ADD02/n11 , \C023/ADD01/ADD02/n10 , \C023/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(65)
  xor \C023/ADD01/ADD02/u29  (complemented_temp_exp_diff[6], \C023/outtemp [6], \C023/ADD01/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  xor \C023/ADD01/ADD02/u33  (complemented_temp_exp_diff[5], \C023/outtemp [5], \C023/ADD01/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \C023/ADD01/ADD02/u34  (complemented_temp_exp_diff[4], \C023/outtemp [4], \C023/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(71)
  and \C023/ADD01/ADD02/u8  (\C023/ADD01/ADD02/n0 , \C023/outtemp [4], \C023/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(63)
  not \C023/C01/u0  (\C023/outtemp [3], temp_exp_diff[3]);  // ../RTL/core/fpu_utils.v(44)
  not \C023/C01/u1  (\C023/outtemp [2], temp_exp_diff[2]);  // ../RTL/core/fpu_utils.v(44)
  not \C023/C01/u2  (\C023/outtemp [1], temp_exp_diff[1]);  // ../RTL/core/fpu_utils.v(44)
  not \C023/C01/u4  (\C023/outtemp [7], temp_exp_diff[7]);  // ../RTL/core/fpu_utils.v(44)
  not \C023/C01/u5  (\C023/outtemp [6], temp_exp_diff[6]);  // ../RTL/core/fpu_utils.v(44)
  not \C023/C01/u6  (\C023/outtemp [5], temp_exp_diff[5]);  // ../RTL/core/fpu_utils.v(44)
  not \C023/C01/u7  (\C023/outtemp [4], temp_exp_diff[4]);  // ../RTL/core/fpu_utils.v(44)
  and \C03/ADD01/ADD01/ADD01/u10  (\C03/ADD01/ADD01/ADD01/n1 , \C03/outtemp [1], \C03/outtemp [0]);  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD01/ADD01/u17  (\C03/ADD01/ADD01/ADD01/n7 , \C03/outtemp [2], \C03/outtemp [1]);  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD01/ADD01/u18  (\C03/ADD01/ADD01/ADD01/n8 , \C03/ADD01/ADD01/ADD01/n7 , \C03/outtemp [0]);  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD01/ADD01/u20  (complemented_M_result[3], \C03/outtemp [3], \C03/ADD01/ADD01/ADD01/n8 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD01/ADD01/u26  (\C03/ADD01/ADD01/ADD01/n14 , \C03/outtemp [3], \C03/outtemp [2]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD01/ADD01/u29  (complemented_M_result[2], \C03/outtemp [2], \C03/ADD01/ADD01/ADD01/n1 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD01/ADD01/u30  (\C03/ADD01/ADD01/ADD01/n17 , \C03/ADD01/ADD01/ADD01/n14 , \C03/outtemp [1]);  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD01/ADD01/u31  (\C03/ADD01/ADD01/ADD01/n18 , \C03/ADD01/ADD01/ADD01/n17 , \C03/outtemp [0]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD01/ADD01/u33  (complemented_M_result[1], \C03/outtemp [1], \C03/outtemp [0]);  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD01/ADD02/u12  (\C03/ADD01/ADD01/ADD02/n3 , \C03/outtemp [5], \C03/outtemp [4]);  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD01/ADD02/u13  (\C03/ADD01/ADD01/ADD02/n4 , \C03/ADD01/ADD01/ADD02/n3 , \C03/ADD01/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD01/ADD02/u17  (\C03/ADD01/ADD01/ADD02/n7 , \C03/outtemp [6], \C03/outtemp [5]);  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD01/ADD02/u20  (complemented_M_result[7], \C03/outtemp [7], \C03/ADD01/ADD01/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD01/ADD02/u21  (\C03/ADD01/ADD01/ADD02/n10 , \C03/ADD01/ADD01/ADD02/n7 , \C03/outtemp [4]);  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD01/ADD02/u22  (\C03/ADD01/ADD01/ADD02/n11 , \C03/ADD01/ADD01/ADD02/n10 , \C03/ADD01/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD01/ADD02/u26  (\C03/ADD01/ADD01/ADD02/n14 , \C03/outtemp [7], \C03/outtemp [6]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD01/ADD02/u29  (complemented_M_result[6], \C03/outtemp [6], \C03/ADD01/ADD01/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD01/ADD02/u30  (\C03/ADD01/ADD01/ADD02/n17 , \C03/ADD01/ADD01/ADD02/n14 , \C03/outtemp [5]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD01/ADD02/u33  (complemented_M_result[5], \C03/outtemp [5], \C03/ADD01/ADD01/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \C03/ADD01/ADD01/ADD02/u34  (complemented_M_result[4], \C03/outtemp [4], \C03/ADD01/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD01/ADD02/u35  (\C03/ADD01/ADD01/ADD02/n20 , \C03/ADD01/ADD01/ADD02/n17 , \C03/outtemp [4]);  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD01/ADD02/u36  (\C03/ADD01/ADD01/ADD02/n21 , \C03/ADD01/ADD01/ADD02/n20 , \C03/ADD01/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD01/ADD02/u8  (\C03/ADD01/ADD01/ADD02/n0 , \C03/outtemp [4], \C03/ADD01/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(63)
  and \C03/ADD01/ADD02/ADD01/u12  (\C03/ADD01/ADD02/ADD01/n3 , \C03/outtemp [9], \C03/outtemp [8]);  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD02/ADD01/u13  (\C03/ADD01/ADD02/ADD01/n4 , \C03/ADD01/ADD02/ADD01/n3 , \C03/ADD01/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD02/ADD01/u17  (\C03/ADD01/ADD02/ADD01/n7 , \C03/outtemp [10], \C03/outtemp [9]);  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD02/ADD01/u20  (complemented_M_result[11], \C03/outtemp [11], \C03/ADD01/ADD02/ADD01/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD02/ADD01/u21  (\C03/ADD01/ADD02/ADD01/n10 , \C03/ADD01/ADD02/ADD01/n7 , \C03/outtemp [8]);  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD02/ADD01/u22  (\C03/ADD01/ADD02/ADD01/n11 , \C03/ADD01/ADD02/ADD01/n10 , \C03/ADD01/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD02/ADD01/u26  (\C03/ADD01/ADD02/ADD01/n14 , \C03/outtemp [11], \C03/outtemp [10]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD02/ADD01/u29  (complemented_M_result[10], \C03/outtemp [10], \C03/ADD01/ADD02/ADD01/n4 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD02/ADD01/u30  (\C03/ADD01/ADD02/ADD01/n17 , \C03/ADD01/ADD02/ADD01/n14 , \C03/outtemp [9]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD02/ADD01/u33  (complemented_M_result[9], \C03/outtemp [9], \C03/ADD01/ADD02/ADD01/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \C03/ADD01/ADD02/ADD01/u34  (complemented_M_result[8], \C03/outtemp [8], \C03/ADD01/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD02/ADD01/u35  (\C03/ADD01/ADD02/ADD01/n20 , \C03/ADD01/ADD02/ADD01/n17 , \C03/outtemp [8]);  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD02/ADD01/u36  (\C03/ADD01/ADD02/ADD01/n21 , \C03/ADD01/ADD02/ADD01/n20 , \C03/ADD01/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD02/ADD01/u8  (\C03/ADD01/ADD02/ADD01/n0 , \C03/outtemp [8], \C03/ADD01/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(63)
  and \C03/ADD01/ADD02/ADD02/u12  (\C03/ADD01/ADD02/ADD02/n3 , \C03/outtemp [13], \C03/outtemp [12]);  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD02/ADD02/u13  (\C03/ADD01/ADD02/ADD02/n4 , \C03/ADD01/ADD02/ADD02/n3 , \C03/ADD01/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD02/ADD02/u17  (\C03/ADD01/ADD02/ADD02/n7 , \C03/outtemp [14], \C03/outtemp [13]);  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD02/ADD02/u20  (complemented_M_result[15], \C03/outtemp [15], \C03/ADD01/ADD02/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD02/ADD02/u21  (\C03/ADD01/ADD02/ADD02/n10 , \C03/ADD01/ADD02/ADD02/n7 , \C03/outtemp [12]);  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD02/ADD02/u22  (\C03/ADD01/ADD02/ADD02/n11 , \C03/ADD01/ADD02/ADD02/n10 , \C03/ADD01/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD02/ADD02/u26  (\C03/ADD01/ADD02/ADD02/n14 , \C03/outtemp [15], \C03/outtemp [14]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD02/ADD02/u29  (complemented_M_result[14], \C03/outtemp [14], \C03/ADD01/ADD02/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD02/ADD02/u30  (\C03/ADD01/ADD02/ADD02/n17 , \C03/ADD01/ADD02/ADD02/n14 , \C03/outtemp [13]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD02/ADD02/u33  (complemented_M_result[13], \C03/outtemp [13], \C03/ADD01/ADD02/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \C03/ADD01/ADD02/ADD02/u34  (complemented_M_result[12], \C03/outtemp [12], \C03/ADD01/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD02/ADD02/u35  (\C03/ADD01/ADD02/ADD02/n20 , \C03/ADD01/ADD02/ADD02/n17 , \C03/outtemp [12]);  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD02/ADD02/u36  (\C03/ADD01/ADD02/ADD02/n21 , \C03/ADD01/ADD02/ADD02/n20 , \C03/ADD01/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD02/ADD02/u8  (\C03/ADD01/ADD02/ADD02/n0 , \C03/outtemp [12], \C03/ADD01/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(63)
  and \C03/ADD01/ADD03/ADD01/u12  (\C03/ADD01/ADD03/ADD01/n3 , \C03/outtemp [17], \C03/outtemp [16]);  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD03/ADD01/u13  (\C03/ADD01/ADD03/ADD01/n4 , \C03/ADD01/ADD03/ADD01/n3 , \C03/ADD01/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD03/ADD01/u17  (\C03/ADD01/ADD03/ADD01/n7 , \C03/outtemp [18], \C03/outtemp [17]);  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD03/ADD01/u20  (complemented_M_result[19], \C03/outtemp [19], \C03/ADD01/ADD03/ADD01/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD03/ADD01/u21  (\C03/ADD01/ADD03/ADD01/n10 , \C03/ADD01/ADD03/ADD01/n7 , \C03/outtemp [16]);  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD03/ADD01/u22  (\C03/ADD01/ADD03/ADD01/n11 , \C03/ADD01/ADD03/ADD01/n10 , \C03/ADD01/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD03/ADD01/u26  (\C03/ADD01/ADD03/ADD01/n14 , \C03/outtemp [19], \C03/outtemp [18]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD03/ADD01/u29  (complemented_M_result[18], \C03/outtemp [18], \C03/ADD01/ADD03/ADD01/n4 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD03/ADD01/u30  (\C03/ADD01/ADD03/ADD01/n17 , \C03/ADD01/ADD03/ADD01/n14 , \C03/outtemp [17]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD03/ADD01/u33  (complemented_M_result[17], \C03/outtemp [17], \C03/ADD01/ADD03/ADD01/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \C03/ADD01/ADD03/ADD01/u34  (complemented_M_result[16], \C03/outtemp [16], \C03/ADD01/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD03/ADD01/u35  (\C03/ADD01/ADD03/ADD01/n20 , \C03/ADD01/ADD03/ADD01/n17 , \C03/outtemp [16]);  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD03/ADD01/u36  (\C03/ADD01/ADD03/ADD01/n21 , \C03/ADD01/ADD03/ADD01/n20 , \C03/ADD01/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD03/ADD01/u8  (\C03/ADD01/ADD03/ADD01/n0 , \C03/outtemp [16], \C03/ADD01/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(63)
  and \C03/ADD01/ADD03/ADD02/u12  (\C03/ADD01/ADD03/ADD02/n3 , \C03/outtemp [21], \C03/outtemp [20]);  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD03/ADD02/u13  (\C03/ADD01/ADD03/ADD02/n4 , \C03/ADD01/ADD03/ADD02/n3 , \C03/ADD01/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD03/ADD02/u17  (\C03/ADD01/ADD03/ADD02/n7 , \C03/outtemp [22], \C03/outtemp [21]);  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD03/ADD02/u20  (complemented_M_result[23], \C03/outtemp [23], \C03/ADD01/ADD03/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD03/ADD02/u21  (\C03/ADD01/ADD03/ADD02/n10 , \C03/ADD01/ADD03/ADD02/n7 , \C03/outtemp [20]);  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD03/ADD02/u22  (\C03/ADD01/ADD03/ADD02/n11 , \C03/ADD01/ADD03/ADD02/n10 , \C03/ADD01/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD03/ADD02/u29  (complemented_M_result[22], \C03/outtemp [22], \C03/ADD01/ADD03/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  xor \C03/ADD01/ADD03/ADD02/u33  (complemented_M_result[21], \C03/outtemp [21], \C03/ADD01/ADD03/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \C03/ADD01/ADD03/ADD02/u34  (complemented_M_result[20], \C03/outtemp [20], \C03/ADD01/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD03/ADD02/u8  (\C03/ADD01/ADD03/ADD02/n0 , \C03/outtemp [20], \C03/ADD01/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(63)
  not \C03/C01/C01/u0  (\C03/outtemp [3], M_result[3]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u1  (\C03/outtemp [2], M_result[2]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u2  (\C03/outtemp [1], M_result[1]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u3  (\C03/outtemp [0], M_result[0]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u4  (\C03/outtemp [7], M_result[7]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u5  (\C03/outtemp [6], M_result[6]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u6  (\C03/outtemp [5], M_result[5]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u7  (\C03/outtemp [4], M_result[4]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u0  (\C03/outtemp [11], M_result[11]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u1  (\C03/outtemp [10], M_result[10]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u2  (\C03/outtemp [9], M_result[9]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u3  (\C03/outtemp [8], M_result[8]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u4  (\C03/outtemp [15], M_result[15]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u5  (\C03/outtemp [14], M_result[14]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u6  (\C03/outtemp [13], M_result[13]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u7  (\C03/outtemp [12], M_result[12]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u0  (\C03/outtemp [19], M_result[19]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u1  (\C03/outtemp [18], M_result[18]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u2  (\C03/outtemp [17], M_result[17]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u3  (\C03/outtemp [16], M_result[16]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u4  (\C03/outtemp [23], M_result[23]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u5  (\C03/outtemp [22], M_result[22]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u6  (\C03/outtemp [21], M_result[21]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u7  (\C03/outtemp [20], M_result[20]);  // ../RTL/core/fpu_utils.v(44)
  not \C04/u0  (complemented_shift_E[3], shift_E[3]);  // ../RTL/core/fpu_utils.v(44)
  not \C04/u1  (complemented_shift_E[2], shift_E[2]);  // ../RTL/core/fpu_utils.v(44)
  not \C04/u2  (complemented_shift_E[1], shift_E[1]);  // ../RTL/core/fpu_utils.v(44)
  not \C04/u3  (complemented_shift_E[0], shift_E[0]);  // ../RTL/core/fpu_utils.v(44)
  not \C04/u7  (complemented_shift_E[4], shift_E[4]);  // ../RTL/core/fpu_utils.v(44)
  AL_MUX \M011/M02/u3  (
    .i0(complemented_temp_exp_diff[1]),
    .i1(temp_exp_diff[1]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[1]));
  AL_MUX \M011/M03/u3  (
    .i0(complemented_temp_exp_diff[2]),
    .i1(temp_exp_diff[2]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[2]));
  AL_MUX \M011/M04/u3  (
    .i0(complemented_temp_exp_diff[3]),
    .i1(temp_exp_diff[3]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[3]));
  AL_MUX \M011/M05/u3  (
    .i0(complemented_temp_exp_diff[4]),
    .i1(temp_exp_diff[4]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[4]));
  AL_MUX \M011/M06/u3  (
    .i0(complemented_temp_exp_diff[5]),
    .i1(temp_exp_diff[5]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[5]));
  AL_MUX \M011/M07/u3  (
    .i0(complemented_temp_exp_diff[6]),
    .i1(temp_exp_diff[6]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[6]));
  AL_MUX \M011/M08/u3  (
    .i0(complemented_temp_exp_diff[7]),
    .i1(temp_exp_diff[7]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[7]));
  AL_MUX \M03/M01/u3  (
    .i0(n2[23]),
    .i1(n1[23]),
    .sel(isE1GreaterThanE2),
    .o(E[0]));
  AL_MUX \M03/M02/u3  (
    .i0(n2[24]),
    .i1(n1[24]),
    .sel(isE1GreaterThanE2),
    .o(E[1]));
  AL_MUX \M03/M03/u3  (
    .i0(n2[25]),
    .i1(n1[25]),
    .sel(isE1GreaterThanE2),
    .o(E[2]));
  AL_MUX \M03/M04/u3  (
    .i0(n2[26]),
    .i1(n1[26]),
    .sel(isE1GreaterThanE2),
    .o(E[3]));
  AL_MUX \M03/M05/u3  (
    .i0(n2[27]),
    .i1(n1[27]),
    .sel(isE1GreaterThanE2),
    .o(E[4]));
  AL_MUX \M03/M06/u3  (
    .i0(n2[28]),
    .i1(n1[28]),
    .sel(isE1GreaterThanE2),
    .o(E[5]));
  AL_MUX \M03/M07/u3  (
    .i0(n2[29]),
    .i1(n1[29]),
    .sel(isE1GreaterThanE2),
    .o(E[6]));
  AL_MUX \M03/M08/u3  (
    .i0(n2[30]),
    .i1(n1[30]),
    .sel(isE1GreaterThanE2),
    .o(E[7]));
  not \M031/M01/u0  (\M031/M01/invSL , \NM/n2 );  // ../RTL/core/fpu_utils.v(106)
  AL_MUX \M031/M01/u3  (
    .i0(\NM/n2 ),
    .i1(\M031/M01/invSL ),
    .sel(E[0]),
    .o(new_E[0]));
  AL_MUX \M031/M02/u3  (
    .i0(E[1]),
    .i1(One_Added_E[1]),
    .sel(\NM/n2 ),
    .o(new_E[1]));
  AL_MUX \M031/M03/u3  (
    .i0(E[2]),
    .i1(One_Added_E[2]),
    .sel(\NM/n2 ),
    .o(new_E[2]));
  AL_MUX \M031/M04/u3  (
    .i0(E[3]),
    .i1(One_Added_E[3]),
    .sel(\NM/n2 ),
    .o(new_E[3]));
  AL_MUX \M031/M05/u3  (
    .i0(E[4]),
    .i1(One_Added_E[4]),
    .sel(\NM/n2 ),
    .o(new_E[4]));
  AL_MUX \M031/M06/u3  (
    .i0(E[5]),
    .i1(One_Added_E[5]),
    .sel(\NM/n2 ),
    .o(new_E[5]));
  AL_MUX \M031/M07/u3  (
    .i0(E[6]),
    .i1(One_Added_E[6]),
    .sel(\NM/n2 ),
    .o(new_E[6]));
  AL_MUX \M031/M08/u3  (
    .i0(E[7]),
    .i1(One_Added_E[7]),
    .sel(\NM/n2 ),
    .o(new_E[7]));
  not \M04/M01/M01/u0  (\M04/M01/M01/invSL , real_oper);  // ../RTL/core/fpu_utils.v(106)
  AL_MUX \M04/M01/M01/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[0]),
    .o(new_M2[0]));
  AL_MUX \M04/M01/M02/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[1]),
    .o(new_M2[1]));
  AL_MUX \M04/M01/M03/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[2]),
    .o(new_M2[2]));
  AL_MUX \M04/M01/M04/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[3]),
    .o(new_M2[3]));
  AL_MUX \M04/M01/M05/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[4]),
    .o(new_M2[4]));
  AL_MUX \M04/M01/M06/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[5]),
    .o(new_M2[5]));
  AL_MUX \M04/M01/M07/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[6]),
    .o(new_M2[6]));
  AL_MUX \M04/M01/M08/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[7]),
    .o(new_M2[7]));
  AL_MUX \M04/M02/M01/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[8]),
    .o(new_M2[8]));
  AL_MUX \M04/M02/M02/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[9]),
    .o(new_M2[9]));
  AL_MUX \M04/M02/M03/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[10]),
    .o(new_M2[10]));
  AL_MUX \M04/M02/M04/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[11]),
    .o(new_M2[11]));
  AL_MUX \M04/M02/M05/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[12]),
    .o(new_M2[12]));
  AL_MUX \M04/M02/M06/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[13]),
    .o(new_M2[13]));
  AL_MUX \M04/M02/M07/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[14]),
    .o(new_M2[14]));
  AL_MUX \M04/M02/M08/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[15]),
    .o(new_M2[15]));
  AL_MUX \M04/M03/M01/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[16]),
    .o(new_M2[16]));
  AL_MUX \M04/M03/M02/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[17]),
    .o(new_M2[17]));
  AL_MUX \M04/M03/M03/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[18]),
    .o(new_M2[18]));
  AL_MUX \M04/M03/M04/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[19]),
    .o(new_M2[19]));
  AL_MUX \M04/M03/M05/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[20]),
    .o(new_M2[20]));
  AL_MUX \M04/M03/M06/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[21]),
    .o(new_M2[21]));
  AL_MUX \M04/M03/M07/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[22]),
    .o(new_M2[22]));
  AL_MUX \M04/M03/M08/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[23]),
    .o(new_M2[23]));
  AL_MUX \M05/M01/M02/u3  (
    .i0(M_result[1]),
    .i1(complemented_M_result[1]),
    .sel(n196),
    .o(M_result2[1]));
  AL_MUX \M05/M01/M03/u3  (
    .i0(M_result[2]),
    .i1(complemented_M_result[2]),
    .sel(n196),
    .o(M_result2[2]));
  AL_MUX \M05/M01/M04/u3  (
    .i0(M_result[3]),
    .i1(complemented_M_result[3]),
    .sel(n196),
    .o(M_result2[3]));
  AL_MUX \M05/M01/M05/u3  (
    .i0(M_result[4]),
    .i1(complemented_M_result[4]),
    .sel(n196),
    .o(M_result2[4]));
  AL_MUX \M05/M01/M06/u3  (
    .i0(M_result[5]),
    .i1(complemented_M_result[5]),
    .sel(n196),
    .o(M_result2[5]));
  AL_MUX \M05/M01/M07/u3  (
    .i0(M_result[6]),
    .i1(complemented_M_result[6]),
    .sel(n196),
    .o(M_result2[6]));
  AL_MUX \M05/M01/M08/u3  (
    .i0(M_result[7]),
    .i1(complemented_M_result[7]),
    .sel(n196),
    .o(M_result2[7]));
  AL_MUX \M05/M02/M01/u3  (
    .i0(M_result[8]),
    .i1(complemented_M_result[8]),
    .sel(n196),
    .o(M_result2[8]));
  AL_MUX \M05/M02/M02/u3  (
    .i0(M_result[9]),
    .i1(complemented_M_result[9]),
    .sel(n196),
    .o(M_result2[9]));
  AL_MUX \M05/M02/M03/u3  (
    .i0(M_result[10]),
    .i1(complemented_M_result[10]),
    .sel(n196),
    .o(M_result2[10]));
  AL_MUX \M05/M02/M04/u3  (
    .i0(M_result[11]),
    .i1(complemented_M_result[11]),
    .sel(n196),
    .o(M_result2[11]));
  AL_MUX \M05/M02/M05/u3  (
    .i0(M_result[12]),
    .i1(complemented_M_result[12]),
    .sel(n196),
    .o(M_result2[12]));
  AL_MUX \M05/M02/M06/u3  (
    .i0(M_result[13]),
    .i1(complemented_M_result[13]),
    .sel(n196),
    .o(M_result2[13]));
  AL_MUX \M05/M02/M07/u3  (
    .i0(M_result[14]),
    .i1(complemented_M_result[14]),
    .sel(n196),
    .o(M_result2[14]));
  AL_MUX \M05/M02/M08/u3  (
    .i0(M_result[15]),
    .i1(complemented_M_result[15]),
    .sel(n196),
    .o(M_result2[15]));
  AL_MUX \M05/M03/M01/u3  (
    .i0(M_result[16]),
    .i1(complemented_M_result[16]),
    .sel(n196),
    .o(M_result2[16]));
  AL_MUX \M05/M03/M02/u3  (
    .i0(M_result[17]),
    .i1(complemented_M_result[17]),
    .sel(n196),
    .o(M_result2[17]));
  AL_MUX \M05/M03/M03/u3  (
    .i0(M_result[18]),
    .i1(complemented_M_result[18]),
    .sel(n196),
    .o(M_result2[18]));
  AL_MUX \M05/M03/M04/u3  (
    .i0(M_result[19]),
    .i1(complemented_M_result[19]),
    .sel(n196),
    .o(M_result2[19]));
  AL_MUX \M05/M03/M05/u3  (
    .i0(M_result[20]),
    .i1(complemented_M_result[20]),
    .sel(n196),
    .o(M_result2[20]));
  AL_MUX \M05/M03/M06/u3  (
    .i0(M_result[21]),
    .i1(complemented_M_result[21]),
    .sel(n196),
    .o(M_result2[21]));
  AL_MUX \M05/M03/M07/u3  (
    .i0(M_result[22]),
    .i1(complemented_M_result[22]),
    .sel(n196),
    .o(M_result2[22]));
  AL_MUX \M05/M03/M08/u3  (
    .i0(M_result[23]),
    .i1(complemented_M_result[23]),
    .sel(n196),
    .o(M_result2[23]));
  add_pu23_pu23_o23_1 \NM/add0  (
    .i0(M_result2[23:1]),
    .i1({22'b0000000000000000000000,M_result[0]}),
    .o(\NM/n4 ));  // ../RTL/core/fpu_utils.v(158)
  eq_w24_1 \NM/eq0  (
    .i0({M_result2[23:1],M_result[0]}),
    .i1(24'b000000000000000000000001),
    .o(\NM/n51 ));  // ../RTL/core/fpu_utils.v(301)
  binary_mux_s1_w1 \NM/mux0_b0  (
    .i0(\NM/n122 [0]),
    .i1(\NM/n4 [0]),
    .sel(\NM/n2 ),
    .o(result[0]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b1  (
    .i0(\NM/sel0_b1/or_B23_al_b50_B24_al_o ),
    .i1(\NM/n4 [1]),
    .sel(\NM/n2 ),
    .o(result[1]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b10  (
    .i0(\NM/sel0_b10/or_or_or_B12_al_b39__o ),
    .i1(\NM/n4 [10]),
    .sel(\NM/n2 ),
    .o(result[10]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b11  (
    .i0(\NM/sel0_b11/or_or_or_B12_al_b39__o ),
    .i1(\NM/n4 [11]),
    .sel(\NM/n2 ),
    .o(result[11]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b12  (
    .i0(\NM/sel0_b12/or_or_or_B12_al_b39__o ),
    .i1(\NM/n4 [12]),
    .sel(\NM/n2 ),
    .o(result[12]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b13  (
    .i0(\NM/n122 [13]),
    .i1(\NM/n4 [13]),
    .sel(\NM/n2 ),
    .o(result[13]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b14  (
    .i0(\NM/n122 [14]),
    .i1(\NM/n4 [14]),
    .sel(\NM/n2 ),
    .o(result[14]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b15  (
    .i0(\NM/n122 [15]),
    .i1(\NM/n4 [15]),
    .sel(\NM/n2 ),
    .o(result[15]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b16  (
    .i0(\NM/n122 [16]),
    .i1(\NM/n4 [16]),
    .sel(\NM/n2 ),
    .o(result[16]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b17  (
    .i0(\NM/n122 [17]),
    .i1(\NM/n4 [17]),
    .sel(\NM/n2 ),
    .o(result[17]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b18  (
    .i0(\NM/n122 [18]),
    .i1(\NM/n4 [18]),
    .sel(\NM/n2 ),
    .o(result[18]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b19  (
    .i0(\NM/n122 [19]),
    .i1(\NM/n4 [19]),
    .sel(\NM/n2 ),
    .o(result[19]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b2  (
    .i0(\NM/sel0_b2/or_or_B21_al_b48_B22_o ),
    .i1(\NM/n4 [2]),
    .sel(\NM/n2 ),
    .o(result[2]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b20  (
    .i0(\NM/n122 [20]),
    .i1(\NM/n4 [20]),
    .sel(\NM/n2 ),
    .o(result[20]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b21  (
    .i0(\NM/n122 [21]),
    .i1(\NM/n4 [21]),
    .sel(\NM/n2 ),
    .o(result[21]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b22  (
    .i0(\NM/n122 [22]),
    .i1(\NM/n4 [22]),
    .sel(\NM/n2 ),
    .o(result[22]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b3  (
    .i0(\NM/sel0_b3/or_or_B21_al_b48_B22_o ),
    .i1(\NM/n4 [3]),
    .sel(\NM/n2 ),
    .o(result[3]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b4  (
    .i0(\NM/sel0_b4/or_or_B18_al_b45_or__o ),
    .i1(\NM/n4 [4]),
    .sel(\NM/n2 ),
    .o(result[4]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b5  (
    .i0(\NM/sel0_b5/or_or_B18_al_b45_or__o ),
    .i1(\NM/n4 [5]),
    .sel(\NM/n2 ),
    .o(result[5]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b6  (
    .i0(\NM/sel0_b6/or_or_B18_al_b45_or__o ),
    .i1(\NM/n4 [6]),
    .sel(\NM/n2 ),
    .o(result[6]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b7  (
    .i0(\NM/sel0_b7/or_or_or_B12_al_b39__o ),
    .i1(\NM/n4 [7]),
    .sel(\NM/n2 ),
    .o(result[7]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b8  (
    .i0(\NM/sel0_b8/or_or_or_B12_al_b39__o ),
    .i1(\NM/n4 [8]),
    .sel(\NM/n2 ),
    .o(result[8]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b9  (
    .i0(\NM/sel0_b9/or_or_or_B12_al_b39__o ),
    .i1(\NM/n4 [9]),
    .sel(\NM/n2 ),
    .o(result[9]));  // ../RTL/core/fpu_utils.v(156)
  AL_MUX \NM/mux1_b0  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\NM/mux1_b0_sel_is_2_o ),
    .o(shift_E[0]));
  and \NM/mux1_b0_sel_is_2  (\NM/mux1_b0_sel_is_2_o , \M031/M01/invSL , \NM/sel1_b0_sel_o );
  AL_MUX \NM/mux1_b1  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\NM/mux1_b1_sel_is_2_o ),
    .o(shift_E[1]));
  and \NM/mux1_b1_sel_is_2  (\NM/mux1_b1_sel_is_2_o , \M031/M01/invSL , \NM/sel1_b1_sel_o );
  AL_MUX \NM/mux1_b2  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\NM/mux1_b2_sel_is_2_o ),
    .o(shift_E[2]));
  and \NM/mux1_b2_sel_is_2  (\NM/mux1_b2_sel_is_2_o , \M031/M01/invSL , \NM/sel1_b2_sel_o );
  AL_MUX \NM/mux1_b3  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\NM/mux1_b3_sel_is_2_o ),
    .o(shift_E[3]));
  and \NM/mux1_b3_sel_is_2  (\NM/mux1_b3_sel_is_2_o , \M031/M01/invSL , \NM/sel1_b3_sel_o );
  AL_MUX \NM/mux1_b4  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\NM/mux1_b4_sel_is_2_o ),
    .o(shift_E[4]));
  and \NM/mux1_b4_sel_is_2  (\NM/mux1_b4_sel_is_2_o , \M031/M01/invSL , \NM/sel1_b4_sel_o );
  AL_MUX \NM/sel0_b0  (
    .i0(1'b0),
    .i1(M_result[0]),
    .sel(M_result2[23]),
    .o(\NM/n122 [0]));  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b1/and_b0_23_al_u23  (\NM/sel0_b1/B23_al_b50 , M_result[0], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b1/and_b0_24_al_u24  (\NM/sel0_b1/B24_al_b51 , M_result2[1], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b1/or_B23_al_b50_B24_al  (\NM/sel0_b1/or_B23_al_b50_B24_al_o , \NM/sel0_b1/B23_al_b50 , \NM/sel0_b1/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_14_al_u14  (\NM/sel0_b10/B14_al_b41 , M_result[0], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_15_al_u15  (\NM/sel0_b10/B15_al_b42 , M_result2[1], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_16_al_u16  (\NM/sel0_b10/B16_al_b43 , M_result2[2], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_17_al_u17  (\NM/sel0_b10/B17_al_b44 , M_result2[3], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_18_al_u18  (\NM/sel0_b10/B18_al_b45 , M_result2[4], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_19_al_u19  (\NM/sel0_b10/B19_al_b46 , M_result2[5], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_20_al_u20  (\NM/sel0_b10/B20_al_b47 , M_result2[6], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_21_al_u21  (\NM/sel0_b10/B21_al_b48 , M_result2[7], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_22_al_u22  (\NM/sel0_b10/B22_al_b49 , M_result2[8], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_23_al_u23  (\NM/sel0_b10/B23_al_b50 , M_result2[9], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_24_al_u24  (\NM/sel0_b10/B24_al_b51 , M_result2[10], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_B15_al_b42_or_B16  (\NM/sel0_b10/or_B15_al_b42_or_B16_o , \NM/sel0_b10/B15_al_b42 , \NM/sel0_b10/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_B16_al_b43_B17_al  (\NM/sel0_b10/or_B16_al_b43_B17_al_o , \NM/sel0_b10/B16_al_b43 , \NM/sel0_b10/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_B18_al_b45_or_B19  (\NM/sel0_b10/or_B18_al_b45_or_B19_o , \NM/sel0_b10/B18_al_b45 , \NM/sel0_b10/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_B19_al_b46_B20_al  (\NM/sel0_b10/or_B19_al_b46_B20_al_o , \NM/sel0_b10/B19_al_b46 , \NM/sel0_b10/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_B21_al_b48_B22_al  (\NM/sel0_b10/or_B21_al_b48_B22_al_o , \NM/sel0_b10/B21_al_b48 , \NM/sel0_b10/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_B23_al_b50_B24_al  (\NM/sel0_b10/or_B23_al_b50_B24_al_o , \NM/sel0_b10/B23_al_b50 , \NM/sel0_b10/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_or_B12_al_b39_or_  (\NM/sel0_b10/or_or_B12_al_b39_or__o , \NM/sel0_b10/B14_al_b41 , \NM/sel0_b10/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_or_B18_al_b45_or_  (\NM/sel0_b10/or_or_B18_al_b45_or__o , \NM/sel0_b10/or_B18_al_b45_or_B19_o , \NM/sel0_b10/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_or_B21_al_b48_B22  (\NM/sel0_b10/or_or_B21_al_b48_B22_o , \NM/sel0_b10/or_B21_al_b48_B22_al_o , \NM/sel0_b10/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_or_or_B12_al_b39_  (\NM/sel0_b10/or_or_or_B12_al_b39__o , \NM/sel0_b10/or_or_B12_al_b39_or__o , \NM/sel0_b10/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_13_al_u13  (\NM/sel0_b11/B13_al_b40 , M_result[0], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_14_al_u14  (\NM/sel0_b11/B14_al_b41 , M_result2[1], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_15_al_u15  (\NM/sel0_b11/B15_al_b42 , M_result2[2], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_16_al_u16  (\NM/sel0_b11/B16_al_b43 , M_result2[3], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_17_al_u17  (\NM/sel0_b11/B17_al_b44 , M_result2[4], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_18_al_u18  (\NM/sel0_b11/B18_al_b45 , M_result2[5], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_19_al_u19  (\NM/sel0_b11/B19_al_b46 , M_result2[6], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_20_al_u20  (\NM/sel0_b11/B20_al_b47 , M_result2[7], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_21_al_u21  (\NM/sel0_b11/B21_al_b48 , M_result2[8], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_22_al_u22  (\NM/sel0_b11/B22_al_b49 , M_result2[9], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_23_al_u23  (\NM/sel0_b11/B23_al_b50 , M_result2[10], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_24_al_u24  (\NM/sel0_b11/B24_al_b51 , M_result2[11], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B13_al_b40_B14_al  (\NM/sel0_b11/or_B13_al_b40_B14_al_o , \NM/sel0_b11/B13_al_b40 , \NM/sel0_b11/B14_al_b41 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B15_al_b42_or_B16  (\NM/sel0_b11/or_B15_al_b42_or_B16_o , \NM/sel0_b11/B15_al_b42 , \NM/sel0_b11/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B16_al_b43_B17_al  (\NM/sel0_b11/or_B16_al_b43_B17_al_o , \NM/sel0_b11/B16_al_b43 , \NM/sel0_b11/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B18_al_b45_or_B19  (\NM/sel0_b11/or_B18_al_b45_or_B19_o , \NM/sel0_b11/B18_al_b45 , \NM/sel0_b11/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B19_al_b46_B20_al  (\NM/sel0_b11/or_B19_al_b46_B20_al_o , \NM/sel0_b11/B19_al_b46 , \NM/sel0_b11/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B21_al_b48_B22_al  (\NM/sel0_b11/or_B21_al_b48_B22_al_o , \NM/sel0_b11/B21_al_b48 , \NM/sel0_b11/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B23_al_b50_B24_al  (\NM/sel0_b11/or_B23_al_b50_B24_al_o , \NM/sel0_b11/B23_al_b50 , \NM/sel0_b11/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_or_B12_al_b39_or_  (\NM/sel0_b11/or_or_B12_al_b39_or__o , \NM/sel0_b11/or_B13_al_b40_B14_al_o , \NM/sel0_b11/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_or_B18_al_b45_or_  (\NM/sel0_b11/or_or_B18_al_b45_or__o , \NM/sel0_b11/or_B18_al_b45_or_B19_o , \NM/sel0_b11/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_or_B21_al_b48_B22  (\NM/sel0_b11/or_or_B21_al_b48_B22_o , \NM/sel0_b11/or_B21_al_b48_B22_al_o , \NM/sel0_b11/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_or_or_B12_al_b39_  (\NM/sel0_b11/or_or_or_B12_al_b39__o , \NM/sel0_b11/or_or_B12_al_b39_or__o , \NM/sel0_b11/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_12_al_u12  (\NM/sel0_b12/B12_al_b39 , M_result[0], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_13_al_u13  (\NM/sel0_b12/B13_al_b40 , M_result2[1], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_14_al_u14  (\NM/sel0_b12/B14_al_b41 , M_result2[2], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_15_al_u15  (\NM/sel0_b12/B15_al_b42 , M_result2[3], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_16_al_u16  (\NM/sel0_b12/B16_al_b43 , M_result2[4], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_17_al_u17  (\NM/sel0_b12/B17_al_b44 , M_result2[5], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_18_al_u18  (\NM/sel0_b12/B18_al_b45 , M_result2[6], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_19_al_u19  (\NM/sel0_b12/B19_al_b46 , M_result2[7], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_20_al_u20  (\NM/sel0_b12/B20_al_b47 , M_result2[8], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_21_al_u21  (\NM/sel0_b12/B21_al_b48 , M_result2[9], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_22_al_u22  (\NM/sel0_b12/B22_al_b49 , M_result2[10], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_23_al_u23  (\NM/sel0_b12/B23_al_b50 , M_result2[11], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_24_al_u24  (\NM/sel0_b12/B24_al_b51 , M_result2[12], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B12_al_b39_or_B13  (\NM/sel0_b12/or_B12_al_b39_or_B13_o , \NM/sel0_b12/B12_al_b39 , \NM/sel0_b12/or_B13_al_b40_B14_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B13_al_b40_B14_al  (\NM/sel0_b12/or_B13_al_b40_B14_al_o , \NM/sel0_b12/B13_al_b40 , \NM/sel0_b12/B14_al_b41 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B15_al_b42_or_B16  (\NM/sel0_b12/or_B15_al_b42_or_B16_o , \NM/sel0_b12/B15_al_b42 , \NM/sel0_b12/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B16_al_b43_B17_al  (\NM/sel0_b12/or_B16_al_b43_B17_al_o , \NM/sel0_b12/B16_al_b43 , \NM/sel0_b12/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B18_al_b45_or_B19  (\NM/sel0_b12/or_B18_al_b45_or_B19_o , \NM/sel0_b12/B18_al_b45 , \NM/sel0_b12/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B19_al_b46_B20_al  (\NM/sel0_b12/or_B19_al_b46_B20_al_o , \NM/sel0_b12/B19_al_b46 , \NM/sel0_b12/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B21_al_b48_B22_al  (\NM/sel0_b12/or_B21_al_b48_B22_al_o , \NM/sel0_b12/B21_al_b48 , \NM/sel0_b12/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B23_al_b50_B24_al  (\NM/sel0_b12/or_B23_al_b50_B24_al_o , \NM/sel0_b12/B23_al_b50 , \NM/sel0_b12/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_or_B12_al_b39_or_  (\NM/sel0_b12/or_or_B12_al_b39_or__o , \NM/sel0_b12/or_B12_al_b39_or_B13_o , \NM/sel0_b12/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_or_B18_al_b45_or_  (\NM/sel0_b12/or_or_B18_al_b45_or__o , \NM/sel0_b12/or_B18_al_b45_or_B19_o , \NM/sel0_b12/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_or_B21_al_b48_B22  (\NM/sel0_b12/or_or_B21_al_b48_B22_o , \NM/sel0_b12/or_B21_al_b48_B22_al_o , \NM/sel0_b12/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_or_or_B12_al_b39_  (\NM/sel0_b12/or_or_or_B12_al_b39__o , \NM/sel0_b12/or_or_B12_al_b39_or__o , \NM/sel0_b12/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_11_al_u11  (\NM/sel0_b13/B11_al_b38 , M_result[0], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_12_al_u12  (\NM/sel0_b13/B12_al_b39 , M_result2[1], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_13_al_u13  (\NM/sel0_b13/B13_al_b40 , M_result2[2], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_14_al_u14  (\NM/sel0_b13/B14_al_b41 , M_result2[3], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_15_al_u15  (\NM/sel0_b13/B15_al_b42 , M_result2[4], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_16_al_u16  (\NM/sel0_b13/B16_al_b43 , M_result2[5], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_17_al_u17  (\NM/sel0_b13/B17_al_b44 , M_result2[6], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_18_al_u18  (\NM/sel0_b13/B18_al_b45 , M_result2[7], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_19_al_u19  (\NM/sel0_b13/B19_al_b46 , M_result2[8], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_20_al_u20  (\NM/sel0_b13/B20_al_b47 , M_result2[9], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_21_al_u21  (\NM/sel0_b13/B21_al_b48 , M_result2[10], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_22_al_u22  (\NM/sel0_b13/B22_al_b49 , M_result2[11], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_23_al_u23  (\NM/sel0_b13/B23_al_b50 , M_result2[12], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_24_al_u24  (\NM/sel0_b13/B24_al_b51 , M_result2[13], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B12_al_b39_or_B13  (\NM/sel0_b13/or_B12_al_b39_or_B13_o , \NM/sel0_b13/B12_al_b39 , \NM/sel0_b13/or_B13_al_b40_B14_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B13_al_b40_B14_al  (\NM/sel0_b13/or_B13_al_b40_B14_al_o , \NM/sel0_b13/B13_al_b40 , \NM/sel0_b13/B14_al_b41 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B15_al_b42_or_B16  (\NM/sel0_b13/or_B15_al_b42_or_B16_o , \NM/sel0_b13/B15_al_b42 , \NM/sel0_b13/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B16_al_b43_B17_al  (\NM/sel0_b13/or_B16_al_b43_B17_al_o , \NM/sel0_b13/B16_al_b43 , \NM/sel0_b13/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B18_al_b45_or_B19  (\NM/sel0_b13/or_B18_al_b45_or_B19_o , \NM/sel0_b13/B18_al_b45 , \NM/sel0_b13/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B19_al_b46_B20_al  (\NM/sel0_b13/or_B19_al_b46_B20_al_o , \NM/sel0_b13/B19_al_b46 , \NM/sel0_b13/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B21_al_b48_B22_al  (\NM/sel0_b13/or_B21_al_b48_B22_al_o , \NM/sel0_b13/B21_al_b48 , \NM/sel0_b13/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B23_al_b50_B24_al  (\NM/sel0_b13/or_B23_al_b50_B24_al_o , \NM/sel0_b13/B23_al_b50 , \NM/sel0_b13/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_or_B12_al_b39_or_  (\NM/sel0_b13/or_or_B12_al_b39_or__o , \NM/sel0_b13/or_B12_al_b39_or_B13_o , \NM/sel0_b13/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_or_B18_al_b45_or_  (\NM/sel0_b13/or_or_B18_al_b45_or__o , \NM/sel0_b13/or_B18_al_b45_or_B19_o , \NM/sel0_b13/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_or_B21_al_b48_B22  (\NM/sel0_b13/or_or_B21_al_b48_B22_o , \NM/sel0_b13/or_B21_al_b48_B22_al_o , \NM/sel0_b13/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_or_or_B12_al_b39_  (\NM/sel0_b13/or_or_or_B12_al_b39__o , \NM/sel0_b13/or_or_B12_al_b39_or__o , \NM/sel0_b13/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_or_or_or_B0_al_b2  (\NM/n122 [13], \NM/sel0_b13/B11_al_b38 , \NM/sel0_b13/or_or_or_B12_al_b39__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_10_al_u10  (\NM/sel0_b14/B10_al_b37 , M_result[0], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_11_al_u11  (\NM/sel0_b14/B11_al_b38 , M_result2[1], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_12_al_u12  (\NM/sel0_b14/B12_al_b39 , M_result2[2], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_13_al_u13  (\NM/sel0_b14/B13_al_b40 , M_result2[3], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_14_al_u14  (\NM/sel0_b14/B14_al_b41 , M_result2[4], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_15_al_u15  (\NM/sel0_b14/B15_al_b42 , M_result2[5], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_16_al_u16  (\NM/sel0_b14/B16_al_b43 , M_result2[6], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_17_al_u17  (\NM/sel0_b14/B17_al_b44 , M_result2[7], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_18_al_u18  (\NM/sel0_b14/B18_al_b45 , M_result2[8], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_19_al_u19  (\NM/sel0_b14/B19_al_b46 , M_result2[9], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_20_al_u20  (\NM/sel0_b14/B20_al_b47 , M_result2[10], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_21_al_u21  (\NM/sel0_b14/B21_al_b48 , M_result2[11], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_22_al_u22  (\NM/sel0_b14/B22_al_b49 , M_result2[12], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_23_al_u23  (\NM/sel0_b14/B23_al_b50 , M_result2[13], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_24_al_u24  (\NM/sel0_b14/B24_al_b51 , M_result2[14], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B10_al_b37_B11_al  (\NM/sel0_b14/or_B10_al_b37_B11_al_o , \NM/sel0_b14/B10_al_b37 , \NM/sel0_b14/B11_al_b38 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B12_al_b39_or_B13  (\NM/sel0_b14/or_B12_al_b39_or_B13_o , \NM/sel0_b14/B12_al_b39 , \NM/sel0_b14/or_B13_al_b40_B14_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B13_al_b40_B14_al  (\NM/sel0_b14/or_B13_al_b40_B14_al_o , \NM/sel0_b14/B13_al_b40 , \NM/sel0_b14/B14_al_b41 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B15_al_b42_or_B16  (\NM/sel0_b14/or_B15_al_b42_or_B16_o , \NM/sel0_b14/B15_al_b42 , \NM/sel0_b14/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B16_al_b43_B17_al  (\NM/sel0_b14/or_B16_al_b43_B17_al_o , \NM/sel0_b14/B16_al_b43 , \NM/sel0_b14/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B18_al_b45_or_B19  (\NM/sel0_b14/or_B18_al_b45_or_B19_o , \NM/sel0_b14/B18_al_b45 , \NM/sel0_b14/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B19_al_b46_B20_al  (\NM/sel0_b14/or_B19_al_b46_B20_al_o , \NM/sel0_b14/B19_al_b46 , \NM/sel0_b14/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B21_al_b48_B22_al  (\NM/sel0_b14/or_B21_al_b48_B22_al_o , \NM/sel0_b14/B21_al_b48 , \NM/sel0_b14/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B23_al_b50_B24_al  (\NM/sel0_b14/or_B23_al_b50_B24_al_o , \NM/sel0_b14/B23_al_b50 , \NM/sel0_b14/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_or_B12_al_b39_or_  (\NM/sel0_b14/or_or_B12_al_b39_or__o , \NM/sel0_b14/or_B12_al_b39_or_B13_o , \NM/sel0_b14/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_or_B18_al_b45_or_  (\NM/sel0_b14/or_or_B18_al_b45_or__o , \NM/sel0_b14/or_B18_al_b45_or_B19_o , \NM/sel0_b14/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_or_B21_al_b48_B22  (\NM/sel0_b14/or_or_B21_al_b48_B22_o , \NM/sel0_b14/or_B21_al_b48_B22_al_o , \NM/sel0_b14/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_or_or_B12_al_b39_  (\NM/sel0_b14/or_or_or_B12_al_b39__o , \NM/sel0_b14/or_or_B12_al_b39_or__o , \NM/sel0_b14/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_or_or_or_B0_al_b2  (\NM/n122 [14], \NM/sel0_b14/or_B10_al_b37_B11_al_o , \NM/sel0_b14/or_or_or_B12_al_b39__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_10_al_u10  (\NM/sel0_b15/B10_al_b37 , M_result2[1], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_11_al_u11  (\NM/sel0_b15/B11_al_b38 , M_result2[2], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_12_al_u12  (\NM/sel0_b15/B12_al_b39 , M_result2[3], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_13_al_u13  (\NM/sel0_b15/B13_al_b40 , M_result2[4], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_14_al_u14  (\NM/sel0_b15/B14_al_b41 , M_result2[5], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_15_al_u15  (\NM/sel0_b15/B15_al_b42 , M_result2[6], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_16_al_u16  (\NM/sel0_b15/B16_al_b43 , M_result2[7], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_17_al_u17  (\NM/sel0_b15/B17_al_b44 , M_result2[8], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_18_al_u18  (\NM/sel0_b15/B18_al_b45 , M_result2[9], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_19_al_u19  (\NM/sel0_b15/B19_al_b46 , M_result2[10], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_20_al_u20  (\NM/sel0_b15/B20_al_b47 , M_result2[11], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_21_al_u21  (\NM/sel0_b15/B21_al_b48 , M_result2[12], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_22_al_u22  (\NM/sel0_b15/B22_al_b49 , M_result2[13], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_23_al_u23  (\NM/sel0_b15/B23_al_b50 , M_result2[14], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_24_al_u24  (\NM/sel0_b15/B24_al_b51 , M_result2[15], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_9_al_u9  (\NM/sel0_b15/B9_al_b36 , M_result[0], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B10_al_b37_B11_al  (\NM/sel0_b15/or_B10_al_b37_B11_al_o , \NM/sel0_b15/B10_al_b37 , \NM/sel0_b15/B11_al_b38 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B12_al_b39_or_B13  (\NM/sel0_b15/or_B12_al_b39_or_B13_o , \NM/sel0_b15/B12_al_b39 , \NM/sel0_b15/or_B13_al_b40_B14_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B13_al_b40_B14_al  (\NM/sel0_b15/or_B13_al_b40_B14_al_o , \NM/sel0_b15/B13_al_b40 , \NM/sel0_b15/B14_al_b41 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B15_al_b42_or_B16  (\NM/sel0_b15/or_B15_al_b42_or_B16_o , \NM/sel0_b15/B15_al_b42 , \NM/sel0_b15/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B16_al_b43_B17_al  (\NM/sel0_b15/or_B16_al_b43_B17_al_o , \NM/sel0_b15/B16_al_b43 , \NM/sel0_b15/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B18_al_b45_or_B19  (\NM/sel0_b15/or_B18_al_b45_or_B19_o , \NM/sel0_b15/B18_al_b45 , \NM/sel0_b15/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B19_al_b46_B20_al  (\NM/sel0_b15/or_B19_al_b46_B20_al_o , \NM/sel0_b15/B19_al_b46 , \NM/sel0_b15/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B21_al_b48_B22_al  (\NM/sel0_b15/or_B21_al_b48_B22_al_o , \NM/sel0_b15/B21_al_b48 , \NM/sel0_b15/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B23_al_b50_B24_al  (\NM/sel0_b15/or_B23_al_b50_B24_al_o , \NM/sel0_b15/B23_al_b50 , \NM/sel0_b15/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B9_al_b36_or_B10_  (\NM/sel0_b15/or_B9_al_b36_or_B10__o , \NM/sel0_b15/B9_al_b36 , \NM/sel0_b15/or_B10_al_b37_B11_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_or_B12_al_b39_or_  (\NM/sel0_b15/or_or_B12_al_b39_or__o , \NM/sel0_b15/or_B12_al_b39_or_B13_o , \NM/sel0_b15/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_or_B18_al_b45_or_  (\NM/sel0_b15/or_or_B18_al_b45_or__o , \NM/sel0_b15/or_B18_al_b45_or_B19_o , \NM/sel0_b15/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_or_B21_al_b48_B22  (\NM/sel0_b15/or_or_B21_al_b48_B22_o , \NM/sel0_b15/or_B21_al_b48_B22_al_o , \NM/sel0_b15/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_or_or_B12_al_b39_  (\NM/sel0_b15/or_or_or_B12_al_b39__o , \NM/sel0_b15/or_or_B12_al_b39_or__o , \NM/sel0_b15/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_or_or_or_B0_al_b2  (\NM/n122 [15], \NM/sel0_b15/or_B9_al_b36_or_B10__o , \NM/sel0_b15/or_or_or_B12_al_b39__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_10_al_u10  (\NM/sel0_b16/B10_al_b37 , M_result2[2], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_11_al_u11  (\NM/sel0_b16/B11_al_b38 , M_result2[3], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_12_al_u12  (\NM/sel0_b16/B12_al_b39 , M_result2[4], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_13_al_u13  (\NM/sel0_b16/B13_al_b40 , M_result2[5], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_14_al_u14  (\NM/sel0_b16/B14_al_b41 , M_result2[6], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_15_al_u15  (\NM/sel0_b16/B15_al_b42 , M_result2[7], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_16_al_u16  (\NM/sel0_b16/B16_al_b43 , M_result2[8], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_17_al_u17  (\NM/sel0_b16/B17_al_b44 , M_result2[9], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_18_al_u18  (\NM/sel0_b16/B18_al_b45 , M_result2[10], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_19_al_u19  (\NM/sel0_b16/B19_al_b46 , M_result2[11], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_20_al_u20  (\NM/sel0_b16/B20_al_b47 , M_result2[12], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_21_al_u21  (\NM/sel0_b16/B21_al_b48 , M_result2[13], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_22_al_u22  (\NM/sel0_b16/B22_al_b49 , M_result2[14], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_23_al_u23  (\NM/sel0_b16/B23_al_b50 , M_result2[15], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_24_al_u24  (\NM/sel0_b16/B24_al_b51 , M_result2[16], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_8_al_u8  (\NM/sel0_b16/B8_al_b35 , M_result[0], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_9_al_u9  (\NM/sel0_b16/B9_al_b36 , M_result2[1], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B10_al_b37_B11_al  (\NM/sel0_b16/or_B10_al_b37_B11_al_o , \NM/sel0_b16/B10_al_b37 , \NM/sel0_b16/B11_al_b38 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B12_al_b39_or_B13  (\NM/sel0_b16/or_B12_al_b39_or_B13_o , \NM/sel0_b16/B12_al_b39 , \NM/sel0_b16/or_B13_al_b40_B14_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B13_al_b40_B14_al  (\NM/sel0_b16/or_B13_al_b40_B14_al_o , \NM/sel0_b16/B13_al_b40 , \NM/sel0_b16/B14_al_b41 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B15_al_b42_or_B16  (\NM/sel0_b16/or_B15_al_b42_or_B16_o , \NM/sel0_b16/B15_al_b42 , \NM/sel0_b16/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B16_al_b43_B17_al  (\NM/sel0_b16/or_B16_al_b43_B17_al_o , \NM/sel0_b16/B16_al_b43 , \NM/sel0_b16/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B18_al_b45_or_B19  (\NM/sel0_b16/or_B18_al_b45_or_B19_o , \NM/sel0_b16/B18_al_b45 , \NM/sel0_b16/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B19_al_b46_B20_al  (\NM/sel0_b16/or_B19_al_b46_B20_al_o , \NM/sel0_b16/B19_al_b46 , \NM/sel0_b16/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B21_al_b48_B22_al  (\NM/sel0_b16/or_B21_al_b48_B22_al_o , \NM/sel0_b16/B21_al_b48 , \NM/sel0_b16/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B23_al_b50_B24_al  (\NM/sel0_b16/or_B23_al_b50_B24_al_o , \NM/sel0_b16/B23_al_b50 , \NM/sel0_b16/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B9_al_b36_or_B10_  (\NM/sel0_b16/or_B9_al_b36_or_B10__o , \NM/sel0_b16/B9_al_b36 , \NM/sel0_b16/or_B10_al_b37_B11_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_or_B12_al_b39_or_  (\NM/sel0_b16/or_or_B12_al_b39_or__o , \NM/sel0_b16/or_B12_al_b39_or_B13_o , \NM/sel0_b16/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_or_B18_al_b45_or_  (\NM/sel0_b16/or_or_B18_al_b45_or__o , \NM/sel0_b16/or_B18_al_b45_or_B19_o , \NM/sel0_b16/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_or_B21_al_b48_B22  (\NM/sel0_b16/or_or_B21_al_b48_B22_o , \NM/sel0_b16/or_B21_al_b48_B22_al_o , \NM/sel0_b16/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_or_B6_al_b33_or_B  (\NM/sel0_b16/or_or_B6_al_b33_or_B_o , \NM/sel0_b16/B8_al_b35 , \NM/sel0_b16/or_B9_al_b36_or_B10__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_or_or_B12_al_b39_  (\NM/sel0_b16/or_or_or_B12_al_b39__o , \NM/sel0_b16/or_or_B12_al_b39_or__o , \NM/sel0_b16/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_or_or_or_B0_al_b2  (\NM/n122 [16], \NM/sel0_b16/or_or_B6_al_b33_or_B_o , \NM/sel0_b16/or_or_or_B12_al_b39__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_10_al_u10  (\NM/sel0_b17/B10_al_b37 , M_result2[3], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_11_al_u11  (\NM/sel0_b17/B11_al_b38 , M_result2[4], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_12_al_u12  (\NM/sel0_b17/B12_al_b39 , M_result2[5], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_13_al_u13  (\NM/sel0_b17/B13_al_b40 , M_result2[6], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_14_al_u14  (\NM/sel0_b17/B14_al_b41 , M_result2[7], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_15_al_u15  (\NM/sel0_b17/B15_al_b42 , M_result2[8], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_16_al_u16  (\NM/sel0_b17/B16_al_b43 , M_result2[9], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_17_al_u17  (\NM/sel0_b17/B17_al_b44 , M_result2[10], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_18_al_u18  (\NM/sel0_b17/B18_al_b45 , M_result2[11], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_19_al_u19  (\NM/sel0_b17/B19_al_b46 , M_result2[12], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_20_al_u20  (\NM/sel0_b17/B20_al_b47 , M_result2[13], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_21_al_u21  (\NM/sel0_b17/B21_al_b48 , M_result2[14], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_22_al_u22  (\NM/sel0_b17/B22_al_b49 , M_result2[15], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_23_al_u23  (\NM/sel0_b17/B23_al_b50 , M_result2[16], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_24_al_u24  (\NM/sel0_b17/B24_al_b51 , M_result2[17], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_7_al_u7  (\NM/sel0_b17/B7_al_b34 , M_result[0], \NM/n101 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_8_al_u8  (\NM/sel0_b17/B8_al_b35 , M_result2[1], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_9_al_u9  (\NM/sel0_b17/B9_al_b36 , M_result2[2], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B10_al_b37_B11_al  (\NM/sel0_b17/or_B10_al_b37_B11_al_o , \NM/sel0_b17/B10_al_b37 , \NM/sel0_b17/B11_al_b38 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B12_al_b39_or_B13  (\NM/sel0_b17/or_B12_al_b39_or_B13_o , \NM/sel0_b17/B12_al_b39 , \NM/sel0_b17/or_B13_al_b40_B14_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B13_al_b40_B14_al  (\NM/sel0_b17/or_B13_al_b40_B14_al_o , \NM/sel0_b17/B13_al_b40 , \NM/sel0_b17/B14_al_b41 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B15_al_b42_or_B16  (\NM/sel0_b17/or_B15_al_b42_or_B16_o , \NM/sel0_b17/B15_al_b42 , \NM/sel0_b17/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B16_al_b43_B17_al  (\NM/sel0_b17/or_B16_al_b43_B17_al_o , \NM/sel0_b17/B16_al_b43 , \NM/sel0_b17/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B18_al_b45_or_B19  (\NM/sel0_b17/or_B18_al_b45_or_B19_o , \NM/sel0_b17/B18_al_b45 , \NM/sel0_b17/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B19_al_b46_B20_al  (\NM/sel0_b17/or_B19_al_b46_B20_al_o , \NM/sel0_b17/B19_al_b46 , \NM/sel0_b17/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B21_al_b48_B22_al  (\NM/sel0_b17/or_B21_al_b48_B22_al_o , \NM/sel0_b17/B21_al_b48 , \NM/sel0_b17/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B23_al_b50_B24_al  (\NM/sel0_b17/or_B23_al_b50_B24_al_o , \NM/sel0_b17/B23_al_b50 , \NM/sel0_b17/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B7_al_b34_B8_al_b  (\NM/sel0_b17/or_B7_al_b34_B8_al_b_o , \NM/sel0_b17/B7_al_b34 , \NM/sel0_b17/B8_al_b35 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B9_al_b36_or_B10_  (\NM/sel0_b17/or_B9_al_b36_or_B10__o , \NM/sel0_b17/B9_al_b36 , \NM/sel0_b17/or_B10_al_b37_B11_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_or_B12_al_b39_or_  (\NM/sel0_b17/or_or_B12_al_b39_or__o , \NM/sel0_b17/or_B12_al_b39_or_B13_o , \NM/sel0_b17/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_or_B18_al_b45_or_  (\NM/sel0_b17/or_or_B18_al_b45_or__o , \NM/sel0_b17/or_B18_al_b45_or_B19_o , \NM/sel0_b17/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_or_B21_al_b48_B22  (\NM/sel0_b17/or_or_B21_al_b48_B22_o , \NM/sel0_b17/or_B21_al_b48_B22_al_o , \NM/sel0_b17/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_or_B6_al_b33_or_B  (\NM/sel0_b17/or_or_B6_al_b33_or_B_o , \NM/sel0_b17/or_B7_al_b34_B8_al_b_o , \NM/sel0_b17/or_B9_al_b36_or_B10__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_or_or_B12_al_b39_  (\NM/sel0_b17/or_or_or_B12_al_b39__o , \NM/sel0_b17/or_or_B12_al_b39_or__o , \NM/sel0_b17/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_or_or_or_B0_al_b2  (\NM/n122 [17], \NM/sel0_b17/or_or_B6_al_b33_or_B_o , \NM/sel0_b17/or_or_or_B12_al_b39__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_10_al_u10  (\NM/sel0_b18/B10_al_b37 , M_result2[4], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_11_al_u11  (\NM/sel0_b18/B11_al_b38 , M_result2[5], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_12_al_u12  (\NM/sel0_b18/B12_al_b39 , M_result2[6], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_13_al_u13  (\NM/sel0_b18/B13_al_b40 , M_result2[7], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_14_al_u14  (\NM/sel0_b18/B14_al_b41 , M_result2[8], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_15_al_u15  (\NM/sel0_b18/B15_al_b42 , M_result2[9], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_16_al_u16  (\NM/sel0_b18/B16_al_b43 , M_result2[10], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_17_al_u17  (\NM/sel0_b18/B17_al_b44 , M_result2[11], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_18_al_u18  (\NM/sel0_b18/B18_al_b45 , M_result2[12], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_19_al_u19  (\NM/sel0_b18/B19_al_b46 , M_result2[13], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_20_al_u20  (\NM/sel0_b18/B20_al_b47 , M_result2[14], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_21_al_u21  (\NM/sel0_b18/B21_al_b48 , M_result2[15], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_22_al_u22  (\NM/sel0_b18/B22_al_b49 , M_result2[16], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_23_al_u23  (\NM/sel0_b18/B23_al_b50 , M_result2[17], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_24_al_u24  (\NM/sel0_b18/B24_al_b51 , M_result2[18], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_6_al_u6  (\NM/sel0_b18/B6_al_b33 , M_result[0], \NM/n104 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_7_al_u7  (\NM/sel0_b18/B7_al_b34 , M_result2[1], \NM/n101 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_8_al_u8  (\NM/sel0_b18/B8_al_b35 , M_result2[2], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_9_al_u9  (\NM/sel0_b18/B9_al_b36 , M_result2[3], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B10_al_b37_B11_al  (\NM/sel0_b18/or_B10_al_b37_B11_al_o , \NM/sel0_b18/B10_al_b37 , \NM/sel0_b18/B11_al_b38 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B12_al_b39_or_B13  (\NM/sel0_b18/or_B12_al_b39_or_B13_o , \NM/sel0_b18/B12_al_b39 , \NM/sel0_b18/or_B13_al_b40_B14_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B13_al_b40_B14_al  (\NM/sel0_b18/or_B13_al_b40_B14_al_o , \NM/sel0_b18/B13_al_b40 , \NM/sel0_b18/B14_al_b41 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B15_al_b42_or_B16  (\NM/sel0_b18/or_B15_al_b42_or_B16_o , \NM/sel0_b18/B15_al_b42 , \NM/sel0_b18/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B16_al_b43_B17_al  (\NM/sel0_b18/or_B16_al_b43_B17_al_o , \NM/sel0_b18/B16_al_b43 , \NM/sel0_b18/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B18_al_b45_or_B19  (\NM/sel0_b18/or_B18_al_b45_or_B19_o , \NM/sel0_b18/B18_al_b45 , \NM/sel0_b18/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B19_al_b46_B20_al  (\NM/sel0_b18/or_B19_al_b46_B20_al_o , \NM/sel0_b18/B19_al_b46 , \NM/sel0_b18/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B21_al_b48_B22_al  (\NM/sel0_b18/or_B21_al_b48_B22_al_o , \NM/sel0_b18/B21_al_b48 , \NM/sel0_b18/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B23_al_b50_B24_al  (\NM/sel0_b18/or_B23_al_b50_B24_al_o , \NM/sel0_b18/B23_al_b50 , \NM/sel0_b18/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B6_al_b33_or_B7_a  (\NM/sel0_b18/or_B6_al_b33_or_B7_a_o , \NM/sel0_b18/B6_al_b33 , \NM/sel0_b18/or_B7_al_b34_B8_al_b_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B7_al_b34_B8_al_b  (\NM/sel0_b18/or_B7_al_b34_B8_al_b_o , \NM/sel0_b18/B7_al_b34 , \NM/sel0_b18/B8_al_b35 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B9_al_b36_or_B10_  (\NM/sel0_b18/or_B9_al_b36_or_B10__o , \NM/sel0_b18/B9_al_b36 , \NM/sel0_b18/or_B10_al_b37_B11_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_or_B12_al_b39_or_  (\NM/sel0_b18/or_or_B12_al_b39_or__o , \NM/sel0_b18/or_B12_al_b39_or_B13_o , \NM/sel0_b18/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_or_B18_al_b45_or_  (\NM/sel0_b18/or_or_B18_al_b45_or__o , \NM/sel0_b18/or_B18_al_b45_or_B19_o , \NM/sel0_b18/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_or_B21_al_b48_B22  (\NM/sel0_b18/or_or_B21_al_b48_B22_o , \NM/sel0_b18/or_B21_al_b48_B22_al_o , \NM/sel0_b18/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_or_B6_al_b33_or_B  (\NM/sel0_b18/or_or_B6_al_b33_or_B_o , \NM/sel0_b18/or_B6_al_b33_or_B7_a_o , \NM/sel0_b18/or_B9_al_b36_or_B10__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_or_or_B12_al_b39_  (\NM/sel0_b18/or_or_or_B12_al_b39__o , \NM/sel0_b18/or_or_B12_al_b39_or__o , \NM/sel0_b18/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_or_or_or_B0_al_b2  (\NM/n122 [18], \NM/sel0_b18/or_or_B6_al_b33_or_B_o , \NM/sel0_b18/or_or_or_B12_al_b39__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_10_al_u10  (\NM/sel0_b19/B10_al_b37 , M_result2[5], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_11_al_u11  (\NM/sel0_b19/B11_al_b38 , M_result2[6], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_12_al_u12  (\NM/sel0_b19/B12_al_b39 , M_result2[7], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_13_al_u13  (\NM/sel0_b19/B13_al_b40 , M_result2[8], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_14_al_u14  (\NM/sel0_b19/B14_al_b41 , M_result2[9], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_15_al_u15  (\NM/sel0_b19/B15_al_b42 , M_result2[10], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_16_al_u16  (\NM/sel0_b19/B16_al_b43 , M_result2[11], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_17_al_u17  (\NM/sel0_b19/B17_al_b44 , M_result2[12], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_18_al_u18  (\NM/sel0_b19/B18_al_b45 , M_result2[13], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_19_al_u19  (\NM/sel0_b19/B19_al_b46 , M_result2[14], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_20_al_u20  (\NM/sel0_b19/B20_al_b47 , M_result2[15], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_21_al_u21  (\NM/sel0_b19/B21_al_b48 , M_result2[16], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_22_al_u22  (\NM/sel0_b19/B22_al_b49 , M_result2[17], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_23_al_u23  (\NM/sel0_b19/B23_al_b50 , M_result2[18], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_24_al_u24  (\NM/sel0_b19/B24_al_b51 , M_result2[19], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_5_al_u5  (\NM/sel0_b19/B5_al_b32 , M_result[0], \NM/n107 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_6_al_u6  (\NM/sel0_b19/B6_al_b33 , M_result2[1], \NM/n104 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_7_al_u7  (\NM/sel0_b19/B7_al_b34 , M_result2[2], \NM/n101 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_8_al_u8  (\NM/sel0_b19/B8_al_b35 , M_result2[3], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_9_al_u9  (\NM/sel0_b19/B9_al_b36 , M_result2[4], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B10_al_b37_B11_al  (\NM/sel0_b19/or_B10_al_b37_B11_al_o , \NM/sel0_b19/B10_al_b37 , \NM/sel0_b19/B11_al_b38 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B12_al_b39_or_B13  (\NM/sel0_b19/or_B12_al_b39_or_B13_o , \NM/sel0_b19/B12_al_b39 , \NM/sel0_b19/or_B13_al_b40_B14_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B13_al_b40_B14_al  (\NM/sel0_b19/or_B13_al_b40_B14_al_o , \NM/sel0_b19/B13_al_b40 , \NM/sel0_b19/B14_al_b41 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B15_al_b42_or_B16  (\NM/sel0_b19/or_B15_al_b42_or_B16_o , \NM/sel0_b19/B15_al_b42 , \NM/sel0_b19/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B16_al_b43_B17_al  (\NM/sel0_b19/or_B16_al_b43_B17_al_o , \NM/sel0_b19/B16_al_b43 , \NM/sel0_b19/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B18_al_b45_or_B19  (\NM/sel0_b19/or_B18_al_b45_or_B19_o , \NM/sel0_b19/B18_al_b45 , \NM/sel0_b19/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B19_al_b46_B20_al  (\NM/sel0_b19/or_B19_al_b46_B20_al_o , \NM/sel0_b19/B19_al_b46 , \NM/sel0_b19/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B21_al_b48_B22_al  (\NM/sel0_b19/or_B21_al_b48_B22_al_o , \NM/sel0_b19/B21_al_b48 , \NM/sel0_b19/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B23_al_b50_B24_al  (\NM/sel0_b19/or_B23_al_b50_B24_al_o , \NM/sel0_b19/B23_al_b50 , \NM/sel0_b19/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B6_al_b33_or_B7_a  (\NM/sel0_b19/or_B6_al_b33_or_B7_a_o , \NM/sel0_b19/B6_al_b33 , \NM/sel0_b19/or_B7_al_b34_B8_al_b_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B7_al_b34_B8_al_b  (\NM/sel0_b19/or_B7_al_b34_B8_al_b_o , \NM/sel0_b19/B7_al_b34 , \NM/sel0_b19/B8_al_b35 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B9_al_b36_or_B10_  (\NM/sel0_b19/or_B9_al_b36_or_B10__o , \NM/sel0_b19/B9_al_b36 , \NM/sel0_b19/or_B10_al_b37_B11_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_B12_al_b39_or_  (\NM/sel0_b19/or_or_B12_al_b39_or__o , \NM/sel0_b19/or_B12_al_b39_or_B13_o , \NM/sel0_b19/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_B18_al_b45_or_  (\NM/sel0_b19/or_or_B18_al_b45_or__o , \NM/sel0_b19/or_B18_al_b45_or_B19_o , \NM/sel0_b19/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_B21_al_b48_B22  (\NM/sel0_b19/or_or_B21_al_b48_B22_o , \NM/sel0_b19/or_B21_al_b48_B22_al_o , \NM/sel0_b19/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_B6_al_b33_or_B  (\NM/sel0_b19/or_or_B6_al_b33_or_B_o , \NM/sel0_b19/or_B6_al_b33_or_B7_a_o , \NM/sel0_b19/or_B9_al_b36_or_B10__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_or_B0_al_b27_o  (\NM/sel0_b19/or_or_or_B0_al_b27_o_o , \NM/sel0_b19/B5_al_b32 , \NM/sel0_b19/or_or_B6_al_b33_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_or_B12_al_b39_  (\NM/sel0_b19/or_or_or_B12_al_b39__o , \NM/sel0_b19/or_or_B12_al_b39_or__o , \NM/sel0_b19/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_or_or_B0_al_b2  (\NM/n122 [19], \NM/sel0_b19/or_or_or_B0_al_b27_o_o , \NM/sel0_b19/or_or_or_B12_al_b39__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b2/and_b0_22_al_u22  (\NM/sel0_b2/B22_al_b49 , M_result[0], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b2/and_b0_23_al_u23  (\NM/sel0_b2/B23_al_b50 , M_result2[1], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b2/and_b0_24_al_u24  (\NM/sel0_b2/B24_al_b51 , M_result2[2], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b2/or_B23_al_b50_B24_al  (\NM/sel0_b2/or_B23_al_b50_B24_al_o , \NM/sel0_b2/B23_al_b50 , \NM/sel0_b2/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b2/or_or_B21_al_b48_B22  (\NM/sel0_b2/or_or_B21_al_b48_B22_o , \NM/sel0_b2/B22_al_b49 , \NM/sel0_b2/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_10_al_u10  (\NM/sel0_b20/B10_al_b37 , M_result2[6], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_11_al_u11  (\NM/sel0_b20/B11_al_b38 , M_result2[7], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_12_al_u12  (\NM/sel0_b20/B12_al_b39 , M_result2[8], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_13_al_u13  (\NM/sel0_b20/B13_al_b40 , M_result2[9], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_14_al_u14  (\NM/sel0_b20/B14_al_b41 , M_result2[10], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_15_al_u15  (\NM/sel0_b20/B15_al_b42 , M_result2[11], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_16_al_u16  (\NM/sel0_b20/B16_al_b43 , M_result2[12], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_17_al_u17  (\NM/sel0_b20/B17_al_b44 , M_result2[13], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_18_al_u18  (\NM/sel0_b20/B18_al_b45 , M_result2[14], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_19_al_u19  (\NM/sel0_b20/B19_al_b46 , M_result2[15], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_20_al_u20  (\NM/sel0_b20/B20_al_b47 , M_result2[16], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_21_al_u21  (\NM/sel0_b20/B21_al_b48 , M_result2[17], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_22_al_u22  (\NM/sel0_b20/B22_al_b49 , M_result2[18], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_23_al_u23  (\NM/sel0_b20/B23_al_b50 , M_result2[19], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_24_al_u24  (\NM/sel0_b20/B24_al_b51 , M_result2[20], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_4_al_u4  (\NM/sel0_b20/B4_al_b31 , M_result[0], \NM/n110 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_5_al_u5  (\NM/sel0_b20/B5_al_b32 , M_result2[1], \NM/n107 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_6_al_u6  (\NM/sel0_b20/B6_al_b33 , M_result2[2], \NM/n104 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_7_al_u7  (\NM/sel0_b20/B7_al_b34 , M_result2[3], \NM/n101 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_8_al_u8  (\NM/sel0_b20/B8_al_b35 , M_result2[4], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_9_al_u9  (\NM/sel0_b20/B9_al_b36 , M_result2[5], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B10_al_b37_B11_al  (\NM/sel0_b20/or_B10_al_b37_B11_al_o , \NM/sel0_b20/B10_al_b37 , \NM/sel0_b20/B11_al_b38 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B12_al_b39_or_B13  (\NM/sel0_b20/or_B12_al_b39_or_B13_o , \NM/sel0_b20/B12_al_b39 , \NM/sel0_b20/or_B13_al_b40_B14_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B13_al_b40_B14_al  (\NM/sel0_b20/or_B13_al_b40_B14_al_o , \NM/sel0_b20/B13_al_b40 , \NM/sel0_b20/B14_al_b41 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B15_al_b42_or_B16  (\NM/sel0_b20/or_B15_al_b42_or_B16_o , \NM/sel0_b20/B15_al_b42 , \NM/sel0_b20/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B16_al_b43_B17_al  (\NM/sel0_b20/or_B16_al_b43_B17_al_o , \NM/sel0_b20/B16_al_b43 , \NM/sel0_b20/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B18_al_b45_or_B19  (\NM/sel0_b20/or_B18_al_b45_or_B19_o , \NM/sel0_b20/B18_al_b45 , \NM/sel0_b20/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B19_al_b46_B20_al  (\NM/sel0_b20/or_B19_al_b46_B20_al_o , \NM/sel0_b20/B19_al_b46 , \NM/sel0_b20/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B21_al_b48_B22_al  (\NM/sel0_b20/or_B21_al_b48_B22_al_o , \NM/sel0_b20/B21_al_b48 , \NM/sel0_b20/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B23_al_b50_B24_al  (\NM/sel0_b20/or_B23_al_b50_B24_al_o , \NM/sel0_b20/B23_al_b50 , \NM/sel0_b20/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B4_al_b31_B5_al_b  (\NM/sel0_b20/or_B4_al_b31_B5_al_b_o , \NM/sel0_b20/B4_al_b31 , \NM/sel0_b20/B5_al_b32 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B6_al_b33_or_B7_a  (\NM/sel0_b20/or_B6_al_b33_or_B7_a_o , \NM/sel0_b20/B6_al_b33 , \NM/sel0_b20/or_B7_al_b34_B8_al_b_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B7_al_b34_B8_al_b  (\NM/sel0_b20/or_B7_al_b34_B8_al_b_o , \NM/sel0_b20/B7_al_b34 , \NM/sel0_b20/B8_al_b35 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B9_al_b36_or_B10_  (\NM/sel0_b20/or_B9_al_b36_or_B10__o , \NM/sel0_b20/B9_al_b36 , \NM/sel0_b20/or_B10_al_b37_B11_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_B12_al_b39_or_  (\NM/sel0_b20/or_or_B12_al_b39_or__o , \NM/sel0_b20/or_B12_al_b39_or_B13_o , \NM/sel0_b20/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_B18_al_b45_or_  (\NM/sel0_b20/or_or_B18_al_b45_or__o , \NM/sel0_b20/or_B18_al_b45_or_B19_o , \NM/sel0_b20/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_B21_al_b48_B22  (\NM/sel0_b20/or_or_B21_al_b48_B22_o , \NM/sel0_b20/or_B21_al_b48_B22_al_o , \NM/sel0_b20/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_B6_al_b33_or_B  (\NM/sel0_b20/or_or_B6_al_b33_or_B_o , \NM/sel0_b20/or_B6_al_b33_or_B7_a_o , \NM/sel0_b20/or_B9_al_b36_or_B10__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_or_B0_al_b27_o  (\NM/sel0_b20/or_or_or_B0_al_b27_o_o , \NM/sel0_b20/or_B4_al_b31_B5_al_b_o , \NM/sel0_b20/or_or_B6_al_b33_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_or_B12_al_b39_  (\NM/sel0_b20/or_or_or_B12_al_b39__o , \NM/sel0_b20/or_or_B12_al_b39_or__o , \NM/sel0_b20/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_or_or_B0_al_b2  (\NM/n122 [20], \NM/sel0_b20/or_or_or_B0_al_b27_o_o , \NM/sel0_b20/or_or_or_B12_al_b39__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_10_al_u10  (\NM/sel0_b21/B10_al_b37 , M_result2[7], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_11_al_u11  (\NM/sel0_b21/B11_al_b38 , M_result2[8], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_12_al_u12  (\NM/sel0_b21/B12_al_b39 , M_result2[9], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_13_al_u13  (\NM/sel0_b21/B13_al_b40 , M_result2[10], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_14_al_u14  (\NM/sel0_b21/B14_al_b41 , M_result2[11], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_15_al_u15  (\NM/sel0_b21/B15_al_b42 , M_result2[12], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_16_al_u16  (\NM/sel0_b21/B16_al_b43 , M_result2[13], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_17_al_u17  (\NM/sel0_b21/B17_al_b44 , M_result2[14], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_18_al_u18  (\NM/sel0_b21/B18_al_b45 , M_result2[15], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_19_al_u19  (\NM/sel0_b21/B19_al_b46 , M_result2[16], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_20_al_u20  (\NM/sel0_b21/B20_al_b47 , M_result2[17], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_21_al_u21  (\NM/sel0_b21/B21_al_b48 , M_result2[18], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_22_al_u22  (\NM/sel0_b21/B22_al_b49 , M_result2[19], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_23_al_u23  (\NM/sel0_b21/B23_al_b50 , M_result2[20], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_24_al_u24  (\NM/sel0_b21/B24_al_b51 , M_result2[21], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_3_al_u3  (\NM/sel0_b21/B3_al_b30 , M_result[0], \NM/n113 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_4_al_u4  (\NM/sel0_b21/B4_al_b31 , M_result2[1], \NM/n110 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_5_al_u5  (\NM/sel0_b21/B5_al_b32 , M_result2[2], \NM/n107 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_6_al_u6  (\NM/sel0_b21/B6_al_b33 , M_result2[3], \NM/n104 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_7_al_u7  (\NM/sel0_b21/B7_al_b34 , M_result2[4], \NM/n101 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_8_al_u8  (\NM/sel0_b21/B8_al_b35 , M_result2[5], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_9_al_u9  (\NM/sel0_b21/B9_al_b36 , M_result2[6], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B10_al_b37_B11_al  (\NM/sel0_b21/or_B10_al_b37_B11_al_o , \NM/sel0_b21/B10_al_b37 , \NM/sel0_b21/B11_al_b38 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B12_al_b39_or_B13  (\NM/sel0_b21/or_B12_al_b39_or_B13_o , \NM/sel0_b21/B12_al_b39 , \NM/sel0_b21/or_B13_al_b40_B14_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B13_al_b40_B14_al  (\NM/sel0_b21/or_B13_al_b40_B14_al_o , \NM/sel0_b21/B13_al_b40 , \NM/sel0_b21/B14_al_b41 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B15_al_b42_or_B16  (\NM/sel0_b21/or_B15_al_b42_or_B16_o , \NM/sel0_b21/B15_al_b42 , \NM/sel0_b21/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B16_al_b43_B17_al  (\NM/sel0_b21/or_B16_al_b43_B17_al_o , \NM/sel0_b21/B16_al_b43 , \NM/sel0_b21/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B18_al_b45_or_B19  (\NM/sel0_b21/or_B18_al_b45_or_B19_o , \NM/sel0_b21/B18_al_b45 , \NM/sel0_b21/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B19_al_b46_B20_al  (\NM/sel0_b21/or_B19_al_b46_B20_al_o , \NM/sel0_b21/B19_al_b46 , \NM/sel0_b21/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B21_al_b48_B22_al  (\NM/sel0_b21/or_B21_al_b48_B22_al_o , \NM/sel0_b21/B21_al_b48 , \NM/sel0_b21/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B23_al_b50_B24_al  (\NM/sel0_b21/or_B23_al_b50_B24_al_o , \NM/sel0_b21/B23_al_b50 , \NM/sel0_b21/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B3_al_b30_or_B4_a  (\NM/sel0_b21/or_B3_al_b30_or_B4_a_o , \NM/sel0_b21/B3_al_b30 , \NM/sel0_b21/or_B4_al_b31_B5_al_b_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B4_al_b31_B5_al_b  (\NM/sel0_b21/or_B4_al_b31_B5_al_b_o , \NM/sel0_b21/B4_al_b31 , \NM/sel0_b21/B5_al_b32 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B6_al_b33_or_B7_a  (\NM/sel0_b21/or_B6_al_b33_or_B7_a_o , \NM/sel0_b21/B6_al_b33 , \NM/sel0_b21/or_B7_al_b34_B8_al_b_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B7_al_b34_B8_al_b  (\NM/sel0_b21/or_B7_al_b34_B8_al_b_o , \NM/sel0_b21/B7_al_b34 , \NM/sel0_b21/B8_al_b35 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B9_al_b36_or_B10_  (\NM/sel0_b21/or_B9_al_b36_or_B10__o , \NM/sel0_b21/B9_al_b36 , \NM/sel0_b21/or_B10_al_b37_B11_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_B12_al_b39_or_  (\NM/sel0_b21/or_or_B12_al_b39_or__o , \NM/sel0_b21/or_B12_al_b39_or_B13_o , \NM/sel0_b21/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_B18_al_b45_or_  (\NM/sel0_b21/or_or_B18_al_b45_or__o , \NM/sel0_b21/or_B18_al_b45_or_B19_o , \NM/sel0_b21/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_B21_al_b48_B22  (\NM/sel0_b21/or_or_B21_al_b48_B22_o , \NM/sel0_b21/or_B21_al_b48_B22_al_o , \NM/sel0_b21/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_B6_al_b33_or_B  (\NM/sel0_b21/or_or_B6_al_b33_or_B_o , \NM/sel0_b21/or_B6_al_b33_or_B7_a_o , \NM/sel0_b21/or_B9_al_b36_or_B10__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_or_B0_al_b27_o  (\NM/sel0_b21/or_or_or_B0_al_b27_o_o , \NM/sel0_b21/or_B3_al_b30_or_B4_a_o , \NM/sel0_b21/or_or_B6_al_b33_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_or_B12_al_b39_  (\NM/sel0_b21/or_or_or_B12_al_b39__o , \NM/sel0_b21/or_or_B12_al_b39_or__o , \NM/sel0_b21/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_or_or_B0_al_b2  (\NM/n122 [21], \NM/sel0_b21/or_or_or_B0_al_b27_o_o , \NM/sel0_b21/or_or_or_B12_al_b39__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_10_al_u10  (\NM/sel0_b22/B10_al_b37 , M_result2[8], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_11_al_u11  (\NM/sel0_b22/B11_al_b38 , M_result2[9], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_12_al_u12  (\NM/sel0_b22/B12_al_b39 , M_result2[10], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_13_al_u13  (\NM/sel0_b22/B13_al_b40 , M_result2[11], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_14_al_u14  (\NM/sel0_b22/B14_al_b41 , M_result2[12], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_15_al_u15  (\NM/sel0_b22/B15_al_b42 , M_result2[13], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_16_al_u16  (\NM/sel0_b22/B16_al_b43 , M_result2[14], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_17_al_u17  (\NM/sel0_b22/B17_al_b44 , M_result2[15], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_18_al_u18  (\NM/sel0_b22/B18_al_b45 , M_result2[16], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_19_al_u19  (\NM/sel0_b22/B19_al_b46 , M_result2[17], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_20_al_u20  (\NM/sel0_b22/B20_al_b47 , M_result2[18], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_21_al_u21  (\NM/sel0_b22/B21_al_b48 , M_result2[19], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_22_al_u22  (\NM/sel0_b22/B22_al_b49 , M_result2[20], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_23_al_u23  (\NM/sel0_b22/B23_al_b50 , M_result2[21], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_24_al_u24  (\NM/sel0_b22/B24_al_b51 , M_result2[22], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_2_al_u2  (\NM/sel0_b22/B2_al_b29 , M_result[0], \NM/n116 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_3_al_u3  (\NM/sel0_b22/B3_al_b30 , M_result2[1], \NM/n113 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_4_al_u4  (\NM/sel0_b22/B4_al_b31 , M_result2[2], \NM/n110 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_5_al_u5  (\NM/sel0_b22/B5_al_b32 , M_result2[3], \NM/n107 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_6_al_u6  (\NM/sel0_b22/B6_al_b33 , M_result2[4], \NM/n104 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_7_al_u7  (\NM/sel0_b22/B7_al_b34 , M_result2[5], \NM/n101 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_8_al_u8  (\NM/sel0_b22/B8_al_b35 , M_result2[6], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_9_al_u9  (\NM/sel0_b22/B9_al_b36 , M_result2[7], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B10_al_b37_B11_al  (\NM/sel0_b22/or_B10_al_b37_B11_al_o , \NM/sel0_b22/B10_al_b37 , \NM/sel0_b22/B11_al_b38 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B12_al_b39_or_B13  (\NM/sel0_b22/or_B12_al_b39_or_B13_o , \NM/sel0_b22/B12_al_b39 , \NM/sel0_b22/or_B13_al_b40_B14_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B13_al_b40_B14_al  (\NM/sel0_b22/or_B13_al_b40_B14_al_o , \NM/sel0_b22/B13_al_b40 , \NM/sel0_b22/B14_al_b41 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B15_al_b42_or_B16  (\NM/sel0_b22/or_B15_al_b42_or_B16_o , \NM/sel0_b22/B15_al_b42 , \NM/sel0_b22/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B16_al_b43_B17_al  (\NM/sel0_b22/or_B16_al_b43_B17_al_o , \NM/sel0_b22/B16_al_b43 , \NM/sel0_b22/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B18_al_b45_or_B19  (\NM/sel0_b22/or_B18_al_b45_or_B19_o , \NM/sel0_b22/B18_al_b45 , \NM/sel0_b22/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B19_al_b46_B20_al  (\NM/sel0_b22/or_B19_al_b46_B20_al_o , \NM/sel0_b22/B19_al_b46 , \NM/sel0_b22/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B21_al_b48_B22_al  (\NM/sel0_b22/or_B21_al_b48_B22_al_o , \NM/sel0_b22/B21_al_b48 , \NM/sel0_b22/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B23_al_b50_B24_al  (\NM/sel0_b22/or_B23_al_b50_B24_al_o , \NM/sel0_b22/B23_al_b50 , \NM/sel0_b22/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B3_al_b30_or_B4_a  (\NM/sel0_b22/or_B3_al_b30_or_B4_a_o , \NM/sel0_b22/B3_al_b30 , \NM/sel0_b22/or_B4_al_b31_B5_al_b_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B4_al_b31_B5_al_b  (\NM/sel0_b22/or_B4_al_b31_B5_al_b_o , \NM/sel0_b22/B4_al_b31 , \NM/sel0_b22/B5_al_b32 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B6_al_b33_or_B7_a  (\NM/sel0_b22/or_B6_al_b33_or_B7_a_o , \NM/sel0_b22/B6_al_b33 , \NM/sel0_b22/or_B7_al_b34_B8_al_b_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B7_al_b34_B8_al_b  (\NM/sel0_b22/or_B7_al_b34_B8_al_b_o , \NM/sel0_b22/B7_al_b34 , \NM/sel0_b22/B8_al_b35 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B9_al_b36_or_B10_  (\NM/sel0_b22/or_B9_al_b36_or_B10__o , \NM/sel0_b22/B9_al_b36 , \NM/sel0_b22/or_B10_al_b37_B11_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_B0_al_b27_or_B  (\NM/sel0_b22/or_or_B0_al_b27_or_B_o , \NM/sel0_b22/B2_al_b29 , \NM/sel0_b22/or_B3_al_b30_or_B4_a_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_B12_al_b39_or_  (\NM/sel0_b22/or_or_B12_al_b39_or__o , \NM/sel0_b22/or_B12_al_b39_or_B13_o , \NM/sel0_b22/or_B15_al_b42_or_B16_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_B18_al_b45_or_  (\NM/sel0_b22/or_or_B18_al_b45_or__o , \NM/sel0_b22/or_B18_al_b45_or_B19_o , \NM/sel0_b22/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_B21_al_b48_B22  (\NM/sel0_b22/or_or_B21_al_b48_B22_o , \NM/sel0_b22/or_B21_al_b48_B22_al_o , \NM/sel0_b22/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_B6_al_b33_or_B  (\NM/sel0_b22/or_or_B6_al_b33_or_B_o , \NM/sel0_b22/or_B6_al_b33_or_B7_a_o , \NM/sel0_b22/or_B9_al_b36_or_B10__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_or_B0_al_b27_o  (\NM/sel0_b22/or_or_or_B0_al_b27_o_o , \NM/sel0_b22/or_or_B0_al_b27_or_B_o , \NM/sel0_b22/or_or_B6_al_b33_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_or_B12_al_b39_  (\NM/sel0_b22/or_or_or_B12_al_b39__o , \NM/sel0_b22/or_or_B12_al_b39_or__o , \NM/sel0_b22/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_or_or_B0_al_b2  (\NM/n122 [22], \NM/sel0_b22/or_or_or_B0_al_b27_o_o , \NM/sel0_b22/or_or_or_B12_al_b39__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b3/and_b0_21_al_u21  (\NM/sel0_b3/B21_al_b48 , M_result[0], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b3/and_b0_22_al_u22  (\NM/sel0_b3/B22_al_b49 , M_result2[1], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b3/and_b0_23_al_u23  (\NM/sel0_b3/B23_al_b50 , M_result2[2], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b3/and_b0_24_al_u24  (\NM/sel0_b3/B24_al_b51 , M_result2[3], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b3/or_B21_al_b48_B22_al  (\NM/sel0_b3/or_B21_al_b48_B22_al_o , \NM/sel0_b3/B21_al_b48 , \NM/sel0_b3/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b3/or_B23_al_b50_B24_al  (\NM/sel0_b3/or_B23_al_b50_B24_al_o , \NM/sel0_b3/B23_al_b50 , \NM/sel0_b3/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b3/or_or_B21_al_b48_B22  (\NM/sel0_b3/or_or_B21_al_b48_B22_o , \NM/sel0_b3/or_B21_al_b48_B22_al_o , \NM/sel0_b3/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b4/and_b0_20_al_u20  (\NM/sel0_b4/B20_al_b47 , M_result[0], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b4/and_b0_21_al_u21  (\NM/sel0_b4/B21_al_b48 , M_result2[1], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b4/and_b0_22_al_u22  (\NM/sel0_b4/B22_al_b49 , M_result2[2], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b4/and_b0_23_al_u23  (\NM/sel0_b4/B23_al_b50 , M_result2[3], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b4/and_b0_24_al_u24  (\NM/sel0_b4/B24_al_b51 , M_result2[4], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b4/or_B21_al_b48_B22_al  (\NM/sel0_b4/or_B21_al_b48_B22_al_o , \NM/sel0_b4/B21_al_b48 , \NM/sel0_b4/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b4/or_B23_al_b50_B24_al  (\NM/sel0_b4/or_B23_al_b50_B24_al_o , \NM/sel0_b4/B23_al_b50 , \NM/sel0_b4/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b4/or_or_B18_al_b45_or_  (\NM/sel0_b4/or_or_B18_al_b45_or__o , \NM/sel0_b4/B20_al_b47 , \NM/sel0_b4/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b4/or_or_B21_al_b48_B22  (\NM/sel0_b4/or_or_B21_al_b48_B22_o , \NM/sel0_b4/or_B21_al_b48_B22_al_o , \NM/sel0_b4/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b5/and_b0_19_al_u19  (\NM/sel0_b5/B19_al_b46 , M_result[0], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b5/and_b0_20_al_u20  (\NM/sel0_b5/B20_al_b47 , M_result2[1], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b5/and_b0_21_al_u21  (\NM/sel0_b5/B21_al_b48 , M_result2[2], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b5/and_b0_22_al_u22  (\NM/sel0_b5/B22_al_b49 , M_result2[3], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b5/and_b0_23_al_u23  (\NM/sel0_b5/B23_al_b50 , M_result2[4], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b5/and_b0_24_al_u24  (\NM/sel0_b5/B24_al_b51 , M_result2[5], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b5/or_B19_al_b46_B20_al  (\NM/sel0_b5/or_B19_al_b46_B20_al_o , \NM/sel0_b5/B19_al_b46 , \NM/sel0_b5/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b5/or_B21_al_b48_B22_al  (\NM/sel0_b5/or_B21_al_b48_B22_al_o , \NM/sel0_b5/B21_al_b48 , \NM/sel0_b5/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b5/or_B23_al_b50_B24_al  (\NM/sel0_b5/or_B23_al_b50_B24_al_o , \NM/sel0_b5/B23_al_b50 , \NM/sel0_b5/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b5/or_or_B18_al_b45_or_  (\NM/sel0_b5/or_or_B18_al_b45_or__o , \NM/sel0_b5/or_B19_al_b46_B20_al_o , \NM/sel0_b5/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b5/or_or_B21_al_b48_B22  (\NM/sel0_b5/or_or_B21_al_b48_B22_o , \NM/sel0_b5/or_B21_al_b48_B22_al_o , \NM/sel0_b5/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_18_al_u18  (\NM/sel0_b6/B18_al_b45 , M_result[0], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_19_al_u19  (\NM/sel0_b6/B19_al_b46 , M_result2[1], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_20_al_u20  (\NM/sel0_b6/B20_al_b47 , M_result2[2], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_21_al_u21  (\NM/sel0_b6/B21_al_b48 , M_result2[3], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_22_al_u22  (\NM/sel0_b6/B22_al_b49 , M_result2[4], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_23_al_u23  (\NM/sel0_b6/B23_al_b50 , M_result2[5], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_24_al_u24  (\NM/sel0_b6/B24_al_b51 , M_result2[6], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b6/or_B18_al_b45_or_B19  (\NM/sel0_b6/or_B18_al_b45_or_B19_o , \NM/sel0_b6/B18_al_b45 , \NM/sel0_b6/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b6/or_B19_al_b46_B20_al  (\NM/sel0_b6/or_B19_al_b46_B20_al_o , \NM/sel0_b6/B19_al_b46 , \NM/sel0_b6/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b6/or_B21_al_b48_B22_al  (\NM/sel0_b6/or_B21_al_b48_B22_al_o , \NM/sel0_b6/B21_al_b48 , \NM/sel0_b6/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b6/or_B23_al_b50_B24_al  (\NM/sel0_b6/or_B23_al_b50_B24_al_o , \NM/sel0_b6/B23_al_b50 , \NM/sel0_b6/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b6/or_or_B18_al_b45_or_  (\NM/sel0_b6/or_or_B18_al_b45_or__o , \NM/sel0_b6/or_B18_al_b45_or_B19_o , \NM/sel0_b6/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b6/or_or_B21_al_b48_B22  (\NM/sel0_b6/or_or_B21_al_b48_B22_o , \NM/sel0_b6/or_B21_al_b48_B22_al_o , \NM/sel0_b6/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_17_al_u17  (\NM/sel0_b7/B17_al_b44 , M_result[0], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_18_al_u18  (\NM/sel0_b7/B18_al_b45 , M_result2[1], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_19_al_u19  (\NM/sel0_b7/B19_al_b46 , M_result2[2], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_20_al_u20  (\NM/sel0_b7/B20_al_b47 , M_result2[3], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_21_al_u21  (\NM/sel0_b7/B21_al_b48 , M_result2[4], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_22_al_u22  (\NM/sel0_b7/B22_al_b49 , M_result2[5], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_23_al_u23  (\NM/sel0_b7/B23_al_b50 , M_result2[6], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_24_al_u24  (\NM/sel0_b7/B24_al_b51 , M_result2[7], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_B18_al_b45_or_B19  (\NM/sel0_b7/or_B18_al_b45_or_B19_o , \NM/sel0_b7/B18_al_b45 , \NM/sel0_b7/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_B19_al_b46_B20_al  (\NM/sel0_b7/or_B19_al_b46_B20_al_o , \NM/sel0_b7/B19_al_b46 , \NM/sel0_b7/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_B21_al_b48_B22_al  (\NM/sel0_b7/or_B21_al_b48_B22_al_o , \NM/sel0_b7/B21_al_b48 , \NM/sel0_b7/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_B23_al_b50_B24_al  (\NM/sel0_b7/or_B23_al_b50_B24_al_o , \NM/sel0_b7/B23_al_b50 , \NM/sel0_b7/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_or_B18_al_b45_or_  (\NM/sel0_b7/or_or_B18_al_b45_or__o , \NM/sel0_b7/or_B18_al_b45_or_B19_o , \NM/sel0_b7/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_or_B21_al_b48_B22  (\NM/sel0_b7/or_or_B21_al_b48_B22_o , \NM/sel0_b7/or_B21_al_b48_B22_al_o , \NM/sel0_b7/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_or_or_B12_al_b39_  (\NM/sel0_b7/or_or_or_B12_al_b39__o , \NM/sel0_b7/B17_al_b44 , \NM/sel0_b7/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_16_al_u16  (\NM/sel0_b8/B16_al_b43 , M_result[0], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_17_al_u17  (\NM/sel0_b8/B17_al_b44 , M_result2[1], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_18_al_u18  (\NM/sel0_b8/B18_al_b45 , M_result2[2], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_19_al_u19  (\NM/sel0_b8/B19_al_b46 , M_result2[3], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_20_al_u20  (\NM/sel0_b8/B20_al_b47 , M_result2[4], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_21_al_u21  (\NM/sel0_b8/B21_al_b48 , M_result2[5], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_22_al_u22  (\NM/sel0_b8/B22_al_b49 , M_result2[6], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_23_al_u23  (\NM/sel0_b8/B23_al_b50 , M_result2[7], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_24_al_u24  (\NM/sel0_b8/B24_al_b51 , M_result2[8], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_B16_al_b43_B17_al  (\NM/sel0_b8/or_B16_al_b43_B17_al_o , \NM/sel0_b8/B16_al_b43 , \NM/sel0_b8/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_B18_al_b45_or_B19  (\NM/sel0_b8/or_B18_al_b45_or_B19_o , \NM/sel0_b8/B18_al_b45 , \NM/sel0_b8/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_B19_al_b46_B20_al  (\NM/sel0_b8/or_B19_al_b46_B20_al_o , \NM/sel0_b8/B19_al_b46 , \NM/sel0_b8/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_B21_al_b48_B22_al  (\NM/sel0_b8/or_B21_al_b48_B22_al_o , \NM/sel0_b8/B21_al_b48 , \NM/sel0_b8/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_B23_al_b50_B24_al  (\NM/sel0_b8/or_B23_al_b50_B24_al_o , \NM/sel0_b8/B23_al_b50 , \NM/sel0_b8/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_or_B18_al_b45_or_  (\NM/sel0_b8/or_or_B18_al_b45_or__o , \NM/sel0_b8/or_B18_al_b45_or_B19_o , \NM/sel0_b8/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_or_B21_al_b48_B22  (\NM/sel0_b8/or_or_B21_al_b48_B22_o , \NM/sel0_b8/or_B21_al_b48_B22_al_o , \NM/sel0_b8/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_or_or_B12_al_b39_  (\NM/sel0_b8/or_or_or_B12_al_b39__o , \NM/sel0_b8/or_B16_al_b43_B17_al_o , \NM/sel0_b8/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_15_al_u15  (\NM/sel0_b9/B15_al_b42 , M_result[0], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_16_al_u16  (\NM/sel0_b9/B16_al_b43 , M_result2[1], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_17_al_u17  (\NM/sel0_b9/B17_al_b44 , M_result2[2], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_18_al_u18  (\NM/sel0_b9/B18_al_b45 , M_result2[3], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_19_al_u19  (\NM/sel0_b9/B19_al_b46 , M_result2[4], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_20_al_u20  (\NM/sel0_b9/B20_al_b47 , M_result2[5], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_21_al_u21  (\NM/sel0_b9/B21_al_b48 , M_result2[6], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_22_al_u22  (\NM/sel0_b9/B22_al_b49 , M_result2[7], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_23_al_u23  (\NM/sel0_b9/B23_al_b50 , M_result2[8], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_24_al_u24  (\NM/sel0_b9/B24_al_b51 , M_result2[9], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_B15_al_b42_or_B16  (\NM/sel0_b9/or_B15_al_b42_or_B16_o , \NM/sel0_b9/B15_al_b42 , \NM/sel0_b9/or_B16_al_b43_B17_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_B16_al_b43_B17_al  (\NM/sel0_b9/or_B16_al_b43_B17_al_o , \NM/sel0_b9/B16_al_b43 , \NM/sel0_b9/B17_al_b44 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_B18_al_b45_or_B19  (\NM/sel0_b9/or_B18_al_b45_or_B19_o , \NM/sel0_b9/B18_al_b45 , \NM/sel0_b9/or_B19_al_b46_B20_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_B19_al_b46_B20_al  (\NM/sel0_b9/or_B19_al_b46_B20_al_o , \NM/sel0_b9/B19_al_b46 , \NM/sel0_b9/B20_al_b47 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_B21_al_b48_B22_al  (\NM/sel0_b9/or_B21_al_b48_B22_al_o , \NM/sel0_b9/B21_al_b48 , \NM/sel0_b9/B22_al_b49 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_B23_al_b50_B24_al  (\NM/sel0_b9/or_B23_al_b50_B24_al_o , \NM/sel0_b9/B23_al_b50 , \NM/sel0_b9/B24_al_b51 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_or_B18_al_b45_or_  (\NM/sel0_b9/or_or_B18_al_b45_or__o , \NM/sel0_b9/or_B18_al_b45_or_B19_o , \NM/sel0_b9/or_or_B21_al_b48_B22_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_or_B21_al_b48_B22  (\NM/sel0_b9/or_or_B21_al_b48_B22_o , \NM/sel0_b9/or_B21_al_b48_B22_al_o , \NM/sel0_b9/or_B23_al_b50_B24_al_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_or_or_B12_al_b39_  (\NM/sel0_b9/or_or_or_B12_al_b39__o , \NM/sel0_b9/or_B15_al_b42_or_B16_o , \NM/sel0_b9/or_or_B18_al_b45_or__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel1_b0_sel  (\NM/sel1_b0_sel_o , \NM/n119 , \NM/n113 , \NM/n107 , \NM/n101 , \NM/n95 , \NM/n89 , \NM/n83 , \NM/n77 , \NM/n71 , \NM/n65 , \NM/n59 , \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel1_b1_sel  (\NM/sel1_b1_sel_o , \NM/n119 , \NM/n116 , \NM/n107 , \NM/n104 , \NM/n95 , \NM/n92 , \NM/n83 , \NM/n80 , \NM/n71 , \NM/n68 , \NM/n59 , \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel1_b2_sel  (\NM/sel1_b2_sel_o , \NM/n119 , \NM/n116 , \NM/n113 , \NM/n110 , \NM/n95 , \NM/n92 , \NM/n89 , \NM/n86 , \NM/n71 , \NM/n68 , \NM/n65 , \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel1_b3_sel  (\NM/sel1_b3_sel_o , \NM/n95 , \NM/n92 , \NM/n89 , \NM/n86 , \NM/n83 , \NM/n80 , \NM/n77 , \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel1_b4_sel  (\NM/sel1_b4_sel_o , \NM/n119 , \NM/n116 , \NM/n113 , \NM/n110 , \NM/n107 , \NM/n104 , \NM/n101 , \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u10  (\NM/n10 , M_result2[20]);  // ../RTL/core/fpu_utils.v(181)
  and \NM/u100  (\NM/n101 , \NM/n39 , \NM/n100 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u101  (\NM/n102 , \NM/n99 , \NM/n39 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u102  (\NM/n103 , \NM/n102 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u103  (\NM/n104 , \NM/n41 , \NM/n103 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u104  (\NM/n105 , \NM/n102 , \NM/n41 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u105  (\NM/n106 , \NM/n105 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u106  (\NM/n107 , \NM/n44 , \NM/n106 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u107  (\NM/n108 , \NM/n105 , \NM/n44 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u108  (\NM/n109 , \NM/n108 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u109  (\NM/n110 , \NM/n46 , \NM/n109 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u11  (\NM/n374 , M_result2[22], M_result2[23]);  // ../RTL/core/fpu_utils.v(175)
  or \NM/u110  (\NM/n111 , \NM/n108 , \NM/n46 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u111  (\NM/n112 , \NM/n111 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u112  (\NM/n113 , \NM/n48 , \NM/n112 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u113  (\NM/n114 , \NM/n111 , \NM/n48 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u114  (\NM/n115 , \NM/n114 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u115  (\NM/n116 , \NM/n50 , \NM/n115 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u116  (\NM/n117 , \NM/n114 , \NM/n50 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u117  (\NM/n118 , \NM/n117 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u118  (\NM/n119 , \NM/n51 , \NM/n118 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u12  (\NM/n12 , M_result2[19]);  // ../RTL/core/fpu_utils.v(187)
  or \NM/u121  (\NM/n124 , M_result2[18], M_result2[19]);  // ../RTL/core/fpu_utils.v(253)
  or \NM/u122  (\NM/n125 , M_result2[16], M_result2[17]);  // ../RTL/core/fpu_utils.v(253)
  or \NM/u123  (\NM/n126 , \NM/n130 , \NM/n127 );  // ../RTL/core/fpu_utils.v(253)
  or \NM/u126  (\NM/n318 , M_result2[4], M_result2[5]);  // ../RTL/core/fpu_utils.v(295)
  or \NM/u127  (\NM/n279 , M_result2[4], \NM/n281 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u128  (\NM/n179 , \NM/n182 , \NM/n180 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u129  (\NM/n127 , \NM/n129 , \NM/n128 );  // ../RTL/core/fpu_utils.v(253)
  or \NM/u13  (\NM/n371 , \NM/n10 , M_result2[21]);  // ../RTL/core/fpu_utils.v(181)
  or \NM/u130  (\NM/n180 , M_result2[21], \NM/n374 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u132  (\NM/n316 , M_result2[3], \NM/n318 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u133  (\NM/n278 , \NM/n283 , \NM/n279 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u134  (\NM/n182 , M_result2[19], M_result2[20]);  // ../RTL/core/fpu_utils.v(265)
  or \NM/u135  (\NM/n128 , M_result2[14], M_result2[15]);  // ../RTL/core/fpu_utils.v(253)
  or \NM/u136  (\NM/n183 , \NM/n185 , \NM/n184 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u137  (\NM/n184 , M_result2[17], M_result2[18]);  // ../RTL/core/fpu_utils.v(265)
  or \NM/u138  (\NM/n314 , \NM/n319 , \NM/n316 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u139  (\NM/n276 , M_result2[8], M_result2[9]);  // ../RTL/core/fpu_utils.v(289)
  not \NM/u14  (\NM/n14 , M_result2[18]);  // ../RTL/core/fpu_utils.v(193)
  or \NM/u140  (\NM/n185 , M_result2[15], M_result2[16]);  // ../RTL/core/fpu_utils.v(265)
  or \NM/u141  (\NM/n129 , M_result2[12], M_result2[13]);  // ../RTL/core/fpu_utils.v(253)
  or \NM/u142  (\NM/n186 , \NM/n191 , \NM/n187 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u143  (\NM/n187 , \NM/n190 , \NM/n188 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u144  (\NM/n313 , M_result2[7], M_result2[8]);  // ../RTL/core/fpu_utils.v(295)
  or \NM/u145  (\NM/n274 , M_result2[7], \NM/n276 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u146  (\NM/n188 , M_result2[12], \NM/n189 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u147  (\NM/n130 , \NM/n132 , \NM/n190 );  // ../RTL/core/fpu_utils.v(253)
  or \NM/u148  (\NM/n189 , M_result2[13], M_result2[14]);  // ../RTL/core/fpu_utils.v(265)
  or \NM/u149  (\NM/n190 , M_result2[10], M_result2[11]);  // ../RTL/core/fpu_utils.v(265)
  or \NM/u15  (\NM/n367 , \NM/n12 , M_result2[20]);  // ../RTL/core/fpu_utils.v(187)
  or \NM/u150  (\NM/n311 , M_result2[6], \NM/n313 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u151  (\NM/n273 , M_result2[11], M_result2[12]);  // ../RTL/core/fpu_utils.v(289)
  or \NM/u152  (\NM/n191 , \NM/n193 , \NM/n276 );  // ../RTL/core/fpu_utils.v(265)
  not \NM/u155  (\NM/n41 , \NM/n194 );  // ../RTL/core/fpu_utils.v(271)
  or \NM/u157  (\NM/n271 , M_result2[10], \NM/n273 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u158  (\NM/n194 , \NM/n222 , \NM/n195 );  // ../RTL/core/fpu_utils.v(271)
  not \NM/u159  (\NM/n37 , \NM/n133 );  // ../RTL/core/fpu_utils.v(259)
  not \NM/u16  (\NM/n16 , M_result2[17]);  // ../RTL/core/fpu_utils.v(199)
  or \NM/u160  (\NM/n195 , \NM/n202 , \NM/n179 );  // ../RTL/core/fpu_utils.v(271)
  or \NM/u162  (\NM/n308 , M_result2[9], \NM/n190 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u163  (\NM/n269 , \NM/n274 , \NM/n271 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u165  (\NM/n133 , \NM/n142 , \NM/n134 );  // ../RTL/core/fpu_utils.v(259)
  or \NM/u168  (\NM/n306 , \NM/n311 , \NM/n308 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u169  (\NM/n268 , \NM/n278 , \NM/n269 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u170  (\NM/n202 , \NM/n128 , \NM/n207 );  // ../RTL/core/fpu_utils.v(271)
  or \NM/u171  (\NM/n134 , \NM/n183 , \NM/n179 );  // ../RTL/core/fpu_utils.v(259)
  or \NM/u172  (\NM/n207 , M_result2[16], \NM/n184 );  // ../RTL/core/fpu_utils.v(271)
  or \NM/u174  (\NM/n304 , \NM/n314 , \NM/n306 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u178  (\NM/n222 , \NM/n247 , \NM/n227 );  // ../RTL/core/fpu_utils.v(271)
  or \NM/u179  (\NM/n227 , \NM/n242 , \NM/n232 );  // ../RTL/core/fpu_utils.v(271)
  not \NM/u18  (\NM/n18 , M_result2[16]);  // ../RTL/core/fpu_utils.v(205)
  or \NM/u182  (\NM/n232 , M_result2[11], \NM/n129 );  // ../RTL/core/fpu_utils.v(271)
  or \NM/u185  (\NM/n242 , M_result2[9], M_result2[10]);  // ../RTL/core/fpu_utils.v(271)
  or \NM/u187  (\NM/n263 , M_result2[15], \NM/n125 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u188  (\NM/n247 , \NM/n257 , \NM/n313 );  // ../RTL/core/fpu_utils.v(271)
  not \NM/u191  (\NM/n44 , \NM/n262 );  // ../RTL/core/fpu_utils.v(277)
  or \NM/u193  (\NM/n261 , \NM/n189 , \NM/n263 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u194  (\NM/n262 , \NM/n312 , \NM/n195 );  // ../RTL/core/fpu_utils.v(277)
  not \NM/u20  (\NM/n20 , M_result2[15]);  // ../RTL/core/fpu_utils.v(211)
  or \NM/u204  (\NM/n296 , \NM/n188 , \NM/n263 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u205  (\NM/n258 , M_result2[18], \NM/n182 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u21  (\NM/n349 , \NM/n18 , M_result2[17]);  // ../RTL/core/fpu_utils.v(205)
  or \NM/u214  (\NM/n312 , \NM/n209 , \NM/n227 );  // ../RTL/core/fpu_utils.v(277)
  or \NM/u219  (\NM/n142 , \NM/n146 , \NM/n143 );  // ../RTL/core/fpu_utils.v(259)
  not \NM/u22  (\NM/n22 , M_result2[14]);  // ../RTL/core/fpu_utils.v(217)
  or \NM/u223  (\NM/n253 , \NM/n258 , \NM/n180 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u224  (\NM/n209 , \NM/n214 , \NM/n211 );  // ../RTL/core/fpu_utils.v(277)
  or \NM/u225  (\NM/n143 , \NM/n273 , \NM/n189 );  // ../RTL/core/fpu_utils.v(259)
  or \NM/u226  (\NM/n211 , M_result2[6], \NM/n213 );  // ../RTL/core/fpu_utils.v(277)
  or \NM/u227  (\NM/n213 , M_result2[7], \NM/n34 );  // ../RTL/core/fpu_utils.v(277)
  or \NM/u229  (\NM/n251 , \NM/n261 , \NM/n253 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u23  (\NM/n341 , \NM/n20 , M_result2[16]);  // ../RTL/core/fpu_utils.v(211)
  not \NM/u230  (\NM/n46 , \NM/n216 );  // ../RTL/core/fpu_utils.v(283)
  or \NM/u232  (\NM/n216 , \NM/n234 , \NM/n251 );  // ../RTL/core/fpu_utils.v(283)
  or \NM/u235  (\NM/n249 , \NM/n268 , \NM/n251 );  // ../RTL/core/fpu_utils.v(289)
  not \NM/u24  (\NM/n24 , M_result2[13]);  // ../RTL/core/fpu_utils.v(223)
  or \NM/u240  (\NM/n286 , \NM/n296 , \NM/n253 );  // ../RTL/core/fpu_utils.v(295)
  not \NM/u241  (\NM/n48 , \NM/n249 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u243  (\NM/n146 , \NM/n176 , \NM/n242 );  // ../RTL/core/fpu_utils.v(259)
  or \NM/u246  (\NM/n284 , \NM/n304 , \NM/n286 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u247  (\NM/n246 , M_result2[6], M_result2[7]);  // ../RTL/core/fpu_utils.v(283)
  or \NM/u25  (\NM/n332 , \NM/n22 , M_result2[15]);  // ../RTL/core/fpu_utils.v(217)
  not \NM/u252  (\NM/n50 , \NM/n284 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u253  (\NM/n244 , M_result2[5], \NM/n246 );  // ../RTL/core/fpu_utils.v(283)
  or \NM/u254  (\NM/n234 , \NM/n243 , \NM/n236 );  // ../RTL/core/fpu_utils.v(283)
  not \NM/u255  (\NM/n39 , \NM/n177 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u256  (\NM/n236 , \NM/n276 , \NM/n271 );  // ../RTL/core/fpu_utils.v(283)
  or \NM/u258  (\NM/n281 , M_result2[5], M_result2[6]);  // ../RTL/core/fpu_utils.v(289)
  or \NM/u259  (\NM/n243 , \NM/n248 , \NM/n244 );  // ../RTL/core/fpu_utils.v(283)
  not \NM/u26  (\NM/n26 , M_result2[12]);  // ../RTL/core/fpu_utils.v(229)
  or \NM/u261  (\NM/n177 , \NM/n186 , \NM/n134 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u264  (\NM/n319 , \NM/n49 , M_result2[2]);  // ../RTL/core/fpu_utils.v(295)
  or \NM/u265  (\NM/n320 , \NM/n260 , \NM/n374 );  // ../RTL/core/fpu_utils.v(253)
  or \NM/u266  (\NM/n315 , \NM/n265 , \NM/n320 );  // ../RTL/core/fpu_utils.v(253)
  or \NM/u267  (\NM/n310 , \NM/n126 , \NM/n315 );  // ../RTL/core/fpu_utils.v(253)
  not \NM/u268  (\NM/n35 , \NM/n310 );  // ../RTL/core/fpu_utils.v(253)
  or \NM/u269  (\NM/n300 , \NM/n32 , \NM/n190 );  // ../RTL/core/fpu_utils.v(247)
  or \NM/u27  (\NM/n322 , \NM/n24 , M_result2[14]);  // ../RTL/core/fpu_utils.v(223)
  or \NM/u273  (\NM/n280 , \NM/n300 , \NM/n127 );  // ../RTL/core/fpu_utils.v(247)
  or \NM/u276  (\NM/n265 , \NM/n125 , \NM/n124 );  // ../RTL/core/fpu_utils.v(247)
  or \NM/u277  (\NM/n260 , M_result2[20], M_result2[21]);  // ../RTL/core/fpu_utils.v(247)
  not \NM/u28  (\NM/n28 , M_result2[11]);  // ../RTL/core/fpu_utils.v(235)
  or \NM/u281  (\NM/n240 , \NM/n280 , \NM/n315 );  // ../RTL/core/fpu_utils.v(247)
  not \NM/u282  (\NM/n33 , \NM/n240 );  // ../RTL/core/fpu_utils.v(247)
  or \NM/u283  (\NM/n230 , \NM/n30 , \NM/n273 );  // ../RTL/core/fpu_utils.v(241)
  or \NM/u286  (\NM/n215 , \NM/n189 , \NM/n185 );  // ../RTL/core/fpu_utils.v(241)
  or \NM/u287  (\NM/n210 , \NM/n230 , \NM/n215 );  // ../RTL/core/fpu_utils.v(241)
  or \NM/u289  (\NM/n175 , M_result2[17], \NM/n124 );  // ../RTL/core/fpu_utils.v(241)
  or \NM/u293  (\NM/n171 , \NM/n175 , \NM/n320 );  // ../RTL/core/fpu_utils.v(241)
  or \NM/u294  (\NM/n170 , \NM/n210 , \NM/n171 );  // ../RTL/core/fpu_utils.v(241)
  not \NM/u295  (\NM/n31 , \NM/n170 );  // ../RTL/core/fpu_utils.v(241)
  or \NM/u296  (\NM/n168 , \NM/n28 , \NM/n129 );  // ../RTL/core/fpu_utils.v(235)
  or \NM/u298  (\NM/n166 , M_result2[14], \NM/n185 );  // ../RTL/core/fpu_utils.v(235)
  or \NM/u299  (\NM/n165 , \NM/n168 , \NM/n166 );  // ../RTL/core/fpu_utils.v(235)
  not \NM/u30  (\NM/n30 , M_result2[10]);  // ../RTL/core/fpu_utils.v(241)
  or \NM/u306  (\NM/n158 , \NM/n165 , \NM/n171 );  // ../RTL/core/fpu_utils.v(235)
  not \NM/u307  (\NM/n29 , \NM/n158 );  // ../RTL/core/fpu_utils.v(235)
  or \NM/u308  (\NM/n156 , \NM/n26 , \NM/n189 );  // ../RTL/core/fpu_utils.v(229)
  or \NM/u311  (\NM/n153 , \NM/n156 , \NM/n263 );  // ../RTL/core/fpu_utils.v(229)
  or \NM/u317  (\NM/n321 , \NM/n153 , \NM/n253 );  // ../RTL/core/fpu_utils.v(229)
  not \NM/u318  (\NM/n27 , \NM/n321 );  // ../RTL/core/fpu_utils.v(229)
  not \NM/u32  (\NM/n32 , M_result2[9]);  // ../RTL/core/fpu_utils.v(247)
  or \NM/u321  (\NM/n325 , \NM/n322 , \NM/n263 );  // ../RTL/core/fpu_utils.v(223)
  or \NM/u327  (\NM/n331 , \NM/n325 , \NM/n253 );  // ../RTL/core/fpu_utils.v(223)
  not \NM/u328  (\NM/n25 , \NM/n331 );  // ../RTL/core/fpu_utils.v(223)
  or \NM/u331  (\NM/n335 , \NM/n332 , \NM/n207 );  // ../RTL/core/fpu_utils.v(217)
  or \NM/u336  (\NM/n340 , \NM/n335 , \NM/n179 );  // ../RTL/core/fpu_utils.v(217)
  not \NM/u337  (\NM/n23 , \NM/n340 );  // ../RTL/core/fpu_utils.v(217)
  or \NM/u339  (\NM/n343 , \NM/n341 , \NM/n184 );  // ../RTL/core/fpu_utils.v(211)
  not \NM/u34  (\NM/n34 , M_result2[8]);  // ../RTL/core/fpu_utils.v(253)
  or \NM/u344  (\NM/n348 , \NM/n343 , \NM/n179 );  // ../RTL/core/fpu_utils.v(211)
  not \NM/u345  (\NM/n21 , \NM/n348 );  // ../RTL/core/fpu_utils.v(211)
  or \NM/u347  (\NM/n351 , \NM/n349 , \NM/n124 );  // ../RTL/core/fpu_utils.v(205)
  or \NM/u351  (\NM/n355 , \NM/n351 , \NM/n320 );  // ../RTL/core/fpu_utils.v(205)
  not \NM/u352  (\NM/n19 , \NM/n355 );  // ../RTL/core/fpu_utils.v(205)
  or \NM/u353  (\NM/n357 , \NM/n16 , \NM/n124 );  // ../RTL/core/fpu_utils.v(199)
  or \NM/u357  (\NM/n361 , \NM/n357 , \NM/n320 );  // ../RTL/core/fpu_utils.v(199)
  not \NM/u358  (\NM/n17 , \NM/n361 );  // ../RTL/core/fpu_utils.v(199)
  or \NM/u359  (\NM/n363 , \NM/n14 , \NM/n182 );  // ../RTL/core/fpu_utils.v(193)
  not \NM/u36  (\NM/n36 , M_result2[7]);  // ../RTL/core/fpu_utils.v(259)
  or \NM/u362  (\NM/n366 , \NM/n363 , \NM/n180 );  // ../RTL/core/fpu_utils.v(193)
  not \NM/u363  (\NM/n15 , \NM/n366 );  // ../RTL/core/fpu_utils.v(193)
  or \NM/u366  (\NM/n370 , \NM/n367 , \NM/n180 );  // ../RTL/core/fpu_utils.v(187)
  not \NM/u367  (\NM/n13 , \NM/n370 );  // ../RTL/core/fpu_utils.v(187)
  or \NM/u369  (\NM/n373 , \NM/n371 , \NM/n374 );  // ../RTL/core/fpu_utils.v(181)
  or \NM/u37  (\NM/n132 , \NM/n34 , M_result2[9]);  // ../RTL/core/fpu_utils.v(253)
  not \NM/u370  (\NM/n11 , \NM/n373 );  // ../RTL/core/fpu_utils.v(181)
  or \NM/u371  (\NM/n375 , \NM/n8 , \NM/n374 );  // ../RTL/core/fpu_utils.v(175)
  not \NM/u372  (\NM/n9 , \NM/n375 );  // ../RTL/core/fpu_utils.v(175)
  not \NM/u373  (\NM/n7 , \NM/n376 );  // ../RTL/core/fpu_utils.v(169)
  not \NM/u38  (\NM/n38 , M_result2[6]);  // ../RTL/core/fpu_utils.v(265)
  or \NM/u39  (\NM/n176 , \NM/n36 , M_result2[8]);  // ../RTL/core/fpu_utils.v(259)
  not \NM/u40  (\NM/n40 , M_result2[5]);  // ../RTL/core/fpu_utils.v(271)
  or \NM/u41  (\NM/n193 , \NM/n38 , M_result2[7]);  // ../RTL/core/fpu_utils.v(265)
  not \NM/u42  (\NM/n42 , M_result2[4]);  // ../RTL/core/fpu_utils.v(277)
  or \NM/u44  (\NM/n257 , \NM/n40 , M_result2[6]);  // ../RTL/core/fpu_utils.v(271)
  not \NM/u45  (\NM/n45 , M_result2[3]);  // ../RTL/core/fpu_utils.v(283)
  or \NM/u46  (\NM/n214 , \NM/n42 , M_result2[5]);  // ../RTL/core/fpu_utils.v(277)
  not \NM/u47  (\NM/n47 , M_result2[2]);  // ../RTL/core/fpu_utils.v(289)
  or \NM/u48  (\NM/n248 , \NM/n45 , M_result2[4]);  // ../RTL/core/fpu_utils.v(283)
  not \NM/u49  (\NM/n49 , M_result2[1]);  // ../RTL/core/fpu_utils.v(295)
  and \NM/u5  (\NM/n2 , M_carry, \M04/M01/M01/invSL );  // ../RTL/core/fpu_utils.v(156)
  or \NM/u50  (\NM/n283 , \NM/n47 , M_result2[3]);  // ../RTL/core/fpu_utils.v(289)
  not \NM/u51  (\NM/n52 , M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/u52  (\NM/n53 , \NM/n7 , \NM/n52 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u53  (\NM/n54 , M_result2[23], \NM/n7 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u54  (\NM/n55 , \NM/n54 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u55  (\NM/n56 , \NM/n9 , \NM/n55 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u56  (\NM/n57 , \NM/n54 , \NM/n9 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u57  (\NM/n58 , \NM/n57 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u58  (\NM/n59 , \NM/n11 , \NM/n58 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u59  (\NM/n60 , \NM/n57 , \NM/n11 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u60  (\NM/n61 , \NM/n60 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u61  (\NM/n62 , \NM/n13 , \NM/n61 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u62  (\NM/n63 , \NM/n60 , \NM/n13 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u63  (\NM/n64 , \NM/n63 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u64  (\NM/n65 , \NM/n15 , \NM/n64 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u65  (\NM/n66 , \NM/n63 , \NM/n15 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u66  (\NM/n67 , \NM/n66 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u67  (\NM/n68 , \NM/n17 , \NM/n67 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u68  (\NM/n69 , \NM/n66 , \NM/n17 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u69  (\NM/n70 , \NM/n69 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u7  (\NM/n6 , M_result2[22]);  // ../RTL/core/fpu_utils.v(169)
  and \NM/u70  (\NM/n71 , \NM/n19 , \NM/n70 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u71  (\NM/n72 , \NM/n69 , \NM/n19 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u72  (\NM/n73 , \NM/n72 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u73  (\NM/n74 , \NM/n21 , \NM/n73 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u74  (\NM/n75 , \NM/n72 , \NM/n21 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u75  (\NM/n76 , \NM/n75 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u76  (\NM/n77 , \NM/n23 , \NM/n76 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u77  (\NM/n78 , \NM/n75 , \NM/n23 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u78  (\NM/n79 , \NM/n78 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u79  (\NM/n80 , \NM/n25 , \NM/n79 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u8  (\NM/n8 , M_result2[21]);  // ../RTL/core/fpu_utils.v(175)
  or \NM/u80  (\NM/n81 , \NM/n78 , \NM/n25 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u81  (\NM/n82 , \NM/n81 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u82  (\NM/n83 , \NM/n27 , \NM/n82 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u83  (\NM/n84 , \NM/n81 , \NM/n27 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u84  (\NM/n85 , \NM/n84 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u85  (\NM/n86 , \NM/n29 , \NM/n85 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u86  (\NM/n87 , \NM/n84 , \NM/n29 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u87  (\NM/n88 , \NM/n87 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u88  (\NM/n89 , \NM/n31 , \NM/n88 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u89  (\NM/n90 , \NM/n87 , \NM/n31 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u9  (\NM/n376 , \NM/n6 , M_result2[23]);  // ../RTL/core/fpu_utils.v(169)
  not \NM/u90  (\NM/n91 , \NM/n90 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u91  (\NM/n92 , \NM/n33 , \NM/n91 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u92  (\NM/n93 , \NM/n90 , \NM/n33 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u93  (\NM/n94 , \NM/n93 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u94  (\NM/n95 , \NM/n35 , \NM/n94 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u95  (\NM/n96 , \NM/n93 , \NM/n35 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u96  (\NM/n97 , \NM/n96 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u97  (\NM/n98 , \NM/n37 , \NM/n97 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u98  (\NM/n99 , \NM/n96 , \NM/n37 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u99  (\NM/n100 , \NM/n99 );  // ../RTL/core/fpu_utils.v(163)
  or \RO01/u0  (\RO01/w1 , n1[24], n1[23]);  // ../RTL/core/fpu_utils.v(14)
  or \RO01/u1  (\RO01/w2 , n1[25], \RO01/w1 );  // ../RTL/core/fpu_utils.v(15)
  or \RO01/u2  (\RO01/w3 , n1[26], \RO01/w2 );  // ../RTL/core/fpu_utils.v(16)
  or \RO01/u3  (\RO01/w4 , n1[27], \RO01/w3 );  // ../RTL/core/fpu_utils.v(17)
  or \RO01/u4  (\RO01/w5 , n1[28], \RO01/w4 );  // ../RTL/core/fpu_utils.v(18)
  or \RO01/u5  (\RO01/w6 , n1[29], \RO01/w5 );  // ../RTL/core/fpu_utils.v(19)
  or \RO01/u6  (reduced_or_E1, n1[30], \RO01/w6 );  // ../RTL/core/fpu_utils.v(20)
  not \exp_diff[4]_inv  (\exp_diff[4]_neg , exp_diff[4]);
  binary_mux_s1_w1 mux0_b0 (
    .i0(n37[0]),
    .i1(n1[0]),
    .sel(isE1GreaterThanE2),
    .o(M1[0]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b1 (
    .i0(n37[1]),
    .i1(n1[1]),
    .sel(isE1GreaterThanE2),
    .o(M1[1]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b10 (
    .i0(n37[10]),
    .i1(n1[10]),
    .sel(isE1GreaterThanE2),
    .o(M1[10]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b11 (
    .i0(n37[11]),
    .i1(n1[11]),
    .sel(isE1GreaterThanE2),
    .o(M1[11]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b12 (
    .i0(n37[12]),
    .i1(n1[12]),
    .sel(isE1GreaterThanE2),
    .o(M1[12]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b13 (
    .i0(n37[13]),
    .i1(n1[13]),
    .sel(isE1GreaterThanE2),
    .o(M1[13]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b14 (
    .i0(n37[14]),
    .i1(n1[14]),
    .sel(isE1GreaterThanE2),
    .o(M1[14]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b15 (
    .i0(n37[15]),
    .i1(n1[15]),
    .sel(isE1GreaterThanE2),
    .o(M1[15]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b16 (
    .i0(n37[16]),
    .i1(n1[16]),
    .sel(isE1GreaterThanE2),
    .o(M1[16]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b17 (
    .i0(n37[17]),
    .i1(n1[17]),
    .sel(isE1GreaterThanE2),
    .o(M1[17]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b18 (
    .i0(n37[18]),
    .i1(n1[18]),
    .sel(isE1GreaterThanE2),
    .o(M1[18]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b19 (
    .i0(n37[19]),
    .i1(n1[19]),
    .sel(isE1GreaterThanE2),
    .o(M1[19]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b2 (
    .i0(n37[2]),
    .i1(n1[2]),
    .sel(isE1GreaterThanE2),
    .o(M1[2]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b20 (
    .i0(n37[20]),
    .i1(n1[20]),
    .sel(isE1GreaterThanE2),
    .o(M1[20]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b21 (
    .i0(n37[21]),
    .i1(n1[21]),
    .sel(isE1GreaterThanE2),
    .o(M1[21]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b22 (
    .i0(n37[22]),
    .i1(n1[22]),
    .sel(isE1GreaterThanE2),
    .o(M1[22]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b23 (
    .i0(n62[23]),
    .i1(reduced_or_E1),
    .sel(isE1GreaterThanE2),
    .o(M1[23]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b3 (
    .i0(n37[3]),
    .i1(n1[3]),
    .sel(isE1GreaterThanE2),
    .o(M1[3]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b4 (
    .i0(n37[4]),
    .i1(n1[4]),
    .sel(isE1GreaterThanE2),
    .o(M1[4]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b5 (
    .i0(n37[5]),
    .i1(n1[5]),
    .sel(isE1GreaterThanE2),
    .o(M1[5]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b6 (
    .i0(n37[6]),
    .i1(n1[6]),
    .sel(isE1GreaterThanE2),
    .o(M1[6]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b7 (
    .i0(n37[7]),
    .i1(n1[7]),
    .sel(isE1GreaterThanE2),
    .o(M1[7]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b8 (
    .i0(n37[8]),
    .i1(n1[8]),
    .sel(isE1GreaterThanE2),
    .o(M1[8]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b9 (
    .i0(n37[9]),
    .i1(n1[9]),
    .sel(isE1GreaterThanE2),
    .o(M1[9]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux1_b0 (
    .i0(n2[0]),
    .i1(n62[0]),
    .sel(isE1GreaterThanE2),
    .o(M2[0]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b1 (
    .i0(n2[1]),
    .i1(n62[1]),
    .sel(isE1GreaterThanE2),
    .o(M2[1]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b10 (
    .i0(n2[10]),
    .i1(n62[10]),
    .sel(isE1GreaterThanE2),
    .o(M2[10]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b11 (
    .i0(n2[11]),
    .i1(n62[11]),
    .sel(isE1GreaterThanE2),
    .o(M2[11]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b12 (
    .i0(n2[12]),
    .i1(n62[12]),
    .sel(isE1GreaterThanE2),
    .o(M2[12]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b13 (
    .i0(n2[13]),
    .i1(n62[13]),
    .sel(isE1GreaterThanE2),
    .o(M2[13]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b14 (
    .i0(n2[14]),
    .i1(n62[14]),
    .sel(isE1GreaterThanE2),
    .o(M2[14]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b15 (
    .i0(n2[15]),
    .i1(n62[15]),
    .sel(isE1GreaterThanE2),
    .o(M2[15]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b16 (
    .i0(n2[16]),
    .i1(n62[16]),
    .sel(isE1GreaterThanE2),
    .o(M2[16]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b17 (
    .i0(n2[17]),
    .i1(n62[17]),
    .sel(isE1GreaterThanE2),
    .o(M2[17]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b18 (
    .i0(n2[18]),
    .i1(n62[18]),
    .sel(isE1GreaterThanE2),
    .o(M2[18]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b19 (
    .i0(n2[19]),
    .i1(n62[19]),
    .sel(isE1GreaterThanE2),
    .o(M2[19]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b2 (
    .i0(n2[2]),
    .i1(n62[2]),
    .sel(isE1GreaterThanE2),
    .o(M2[2]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b20 (
    .i0(n2[20]),
    .i1(n62[20]),
    .sel(isE1GreaterThanE2),
    .o(M2[20]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b21 (
    .i0(n2[21]),
    .i1(n62[21]),
    .sel(isE1GreaterThanE2),
    .o(M2[21]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b22 (
    .i0(n2[22]),
    .i1(n62[22]),
    .sel(isE1GreaterThanE2),
    .o(M2[22]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b23 (
    .i0(reduced_or_E1),
    .i1(n62[23]),
    .sel(isE1GreaterThanE2),
    .o(M2[23]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b3 (
    .i0(n2[3]),
    .i1(n62[3]),
    .sel(isE1GreaterThanE2),
    .o(M2[3]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b4 (
    .i0(n2[4]),
    .i1(n62[4]),
    .sel(isE1GreaterThanE2),
    .o(M2[4]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b5 (
    .i0(n2[5]),
    .i1(n62[5]),
    .sel(isE1GreaterThanE2),
    .o(M2[5]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b6 (
    .i0(n2[6]),
    .i1(n62[6]),
    .sel(isE1GreaterThanE2),
    .o(M2[6]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b7 (
    .i0(n2[7]),
    .i1(n62[7]),
    .sel(isE1GreaterThanE2),
    .o(M2[7]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b8 (
    .i0(n2[8]),
    .i1(n62[8]),
    .sel(isE1GreaterThanE2),
    .o(M2[8]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b9 (
    .i0(n2[9]),
    .i1(n62[9]),
    .sel(isE1GreaterThanE2),
    .o(M2[9]));  // ../RTL/core/fpu.v(128)
  not n110_inv (n110_neg, n110);
  not \new_E[5]_inv  (\new_E[5]_neg , new_E[5]);
  not \new_E[6]_inv  (\new_E[6]_neg , new_E[6]);
  not \new_E[7]_inv  (\new_E[7]_neg , new_E[7]);
  AL_MUX u100 (
    .i0(n229),
    .i1(n227),
    .sel(exp_diff[1]),
    .o(n123));  // ../RTL/core/fpu.v(128)
  AL_MUX u101 (
    .i0(n228),
    .i1(n226),
    .sel(exp_diff[1]),
    .o(n122));  // ../RTL/core/fpu.v(128)
  AL_MUX u102 (
    .i0(n227),
    .i1(n225),
    .sel(exp_diff[1]),
    .o(n121));  // ../RTL/core/fpu.v(128)
  AL_MUX u103 (
    .i0(n226),
    .i1(n224),
    .sel(exp_diff[1]),
    .o(n120));  // ../RTL/core/fpu.v(128)
  AL_MUX u104 (
    .i0(n225),
    .i1(n223),
    .sel(exp_diff[1]),
    .o(n119));  // ../RTL/core/fpu.v(128)
  AL_MUX u105 (
    .i0(n224),
    .i1(n222),
    .sel(exp_diff[1]),
    .o(n118));  // ../RTL/core/fpu.v(128)
  AL_MUX u106 (
    .i0(n223),
    .i1(n221),
    .sel(exp_diff[1]),
    .o(n117));  // ../RTL/core/fpu.v(128)
  AL_MUX u107 (
    .i0(n222),
    .i1(n165),
    .sel(exp_diff[1]),
    .o(n116));  // ../RTL/core/fpu.v(128)
  AL_MUX u108 (
    .i0(n221),
    .i1(n164),
    .sel(exp_diff[1]),
    .o(n115));  // ../RTL/core/fpu.v(128)
  AL_MUX u109 (
    .i0(n165),
    .i1(n86),
    .sel(exp_diff[1]),
    .o(n114));  // ../RTL/core/fpu.v(128)
  AL_MUX u110 (
    .i0(n164),
    .i1(1'b0),
    .sel(exp_diff[1]),
    .o(n113));  // ../RTL/core/fpu.v(128)
  AL_MUX u111 (
    .i0(n86),
    .i1(1'b0),
    .sel(exp_diff[1]),
    .o(n112));  // ../RTL/core/fpu.v(128)
  AL_MUX u112 (
    .i0(n161),
    .i1(n131),
    .sel(exp_diff[2]),
    .o(n111));  // ../RTL/core/fpu.v(128)
  AL_MUX u113 (
    .i0(n134),
    .i1(n130),
    .sel(exp_diff[2]),
    .o(n220));  // ../RTL/core/fpu.v(128)
  AL_MUX u114 (
    .i0(n133),
    .i1(n129),
    .sel(exp_diff[2]),
    .o(n219));  // ../RTL/core/fpu.v(128)
  AL_MUX u115 (
    .i0(n132),
    .i1(n128),
    .sel(exp_diff[2]),
    .o(n218));  // ../RTL/core/fpu.v(128)
  AL_MUX u116 (
    .i0(n131),
    .i1(n127),
    .sel(exp_diff[2]),
    .o(n217));  // ../RTL/core/fpu.v(128)
  AL_MUX u117 (
    .i0(n130),
    .i1(n126),
    .sel(exp_diff[2]),
    .o(n216));  // ../RTL/core/fpu.v(128)
  AL_MUX u118 (
    .i0(n129),
    .i1(n125),
    .sel(exp_diff[2]),
    .o(n215));  // ../RTL/core/fpu.v(128)
  AL_MUX u119 (
    .i0(n128),
    .i1(n124),
    .sel(exp_diff[2]),
    .o(n214));  // ../RTL/core/fpu.v(128)
  and u12 (w2, \M04/M01/M01/invSL , n1[31]);  // ../RTL/core/fpu.v(141)
  AL_MUX u120 (
    .i0(n127),
    .i1(n123),
    .sel(exp_diff[2]),
    .o(n213));  // ../RTL/core/fpu.v(128)
  AL_MUX u121 (
    .i0(n126),
    .i1(n122),
    .sel(exp_diff[2]),
    .o(n212));  // ../RTL/core/fpu.v(128)
  AL_MUX u122 (
    .i0(n125),
    .i1(n121),
    .sel(exp_diff[2]),
    .o(n211));  // ../RTL/core/fpu.v(128)
  AL_MUX u123 (
    .i0(n124),
    .i1(n120),
    .sel(exp_diff[2]),
    .o(n210));  // ../RTL/core/fpu.v(128)
  AL_MUX u124 (
    .i0(n123),
    .i1(n119),
    .sel(exp_diff[2]),
    .o(n209));  // ../RTL/core/fpu.v(128)
  AL_MUX u125 (
    .i0(n122),
    .i1(n118),
    .sel(exp_diff[2]),
    .o(n208));  // ../RTL/core/fpu.v(128)
  AL_MUX u126 (
    .i0(n121),
    .i1(n117),
    .sel(exp_diff[2]),
    .o(n207));  // ../RTL/core/fpu.v(128)
  AL_MUX u127 (
    .i0(n120),
    .i1(n116),
    .sel(exp_diff[2]),
    .o(n206));  // ../RTL/core/fpu.v(128)
  AL_MUX u128 (
    .i0(n119),
    .i1(n115),
    .sel(exp_diff[2]),
    .o(n205));  // ../RTL/core/fpu.v(128)
  AL_MUX u129 (
    .i0(n118),
    .i1(n114),
    .sel(exp_diff[2]),
    .o(n204));  // ../RTL/core/fpu.v(128)
  and u13 (w3, M_carry, n1[31]);  // ../RTL/core/fpu.v(142)
  AL_MUX u130 (
    .i0(n117),
    .i1(n113),
    .sel(exp_diff[2]),
    .o(n203));  // ../RTL/core/fpu.v(128)
  AL_MUX u131 (
    .i0(n116),
    .i1(n112),
    .sel(exp_diff[2]),
    .o(n202));  // ../RTL/core/fpu.v(128)
  AL_MUX u132 (
    .i0(n115),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n201));  // ../RTL/core/fpu.v(128)
  AL_MUX u133 (
    .i0(n114),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n200));  // ../RTL/core/fpu.v(128)
  AL_MUX u134 (
    .i0(n113),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n199));  // ../RTL/core/fpu.v(128)
  AL_MUX u135 (
    .i0(n112),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n198));  // ../RTL/core/fpu.v(128)
  AL_MUX u136 (
    .i0(n111),
    .i1(n213),
    .sel(exp_diff[3]),
    .o(n197));  // ../RTL/core/fpu.v(128)
  AL_MUX u137 (
    .i0(n220),
    .i1(n212),
    .sel(exp_diff[3]),
    .o(n158));  // ../RTL/core/fpu.v(128)
  AL_MUX u138 (
    .i0(n219),
    .i1(n211),
    .sel(exp_diff[3]),
    .o(n157));  // ../RTL/core/fpu.v(128)
  AL_MUX u139 (
    .i0(n218),
    .i1(n210),
    .sel(exp_diff[3]),
    .o(n156));  // ../RTL/core/fpu.v(128)
  and u14 (n243, real_oper, n159);  // ../RTL/core/fpu.v(140)
  AL_MUX u140 (
    .i0(n217),
    .i1(n209),
    .sel(exp_diff[3]),
    .o(n155));  // ../RTL/core/fpu.v(128)
  AL_MUX u141 (
    .i0(n216),
    .i1(n208),
    .sel(exp_diff[3]),
    .o(n154));  // ../RTL/core/fpu.v(128)
  AL_MUX u142 (
    .i0(n215),
    .i1(n207),
    .sel(exp_diff[3]),
    .o(n153));  // ../RTL/core/fpu.v(128)
  AL_MUX u143 (
    .i0(n214),
    .i1(n206),
    .sel(exp_diff[3]),
    .o(n152));  // ../RTL/core/fpu.v(128)
  AL_MUX u144 (
    .i0(n213),
    .i1(n205),
    .sel(exp_diff[3]),
    .o(n151));  // ../RTL/core/fpu.v(128)
  AL_MUX u145 (
    .i0(n212),
    .i1(n204),
    .sel(exp_diff[3]),
    .o(n150));  // ../RTL/core/fpu.v(128)
  AL_MUX u146 (
    .i0(n211),
    .i1(n203),
    .sel(exp_diff[3]),
    .o(n149));  // ../RTL/core/fpu.v(128)
  AL_MUX u147 (
    .i0(n210),
    .i1(n202),
    .sel(exp_diff[3]),
    .o(n148));  // ../RTL/core/fpu.v(128)
  AL_MUX u148 (
    .i0(n209),
    .i1(n201),
    .sel(exp_diff[3]),
    .o(n147));  // ../RTL/core/fpu.v(128)
  AL_MUX u149 (
    .i0(n208),
    .i1(n200),
    .sel(exp_diff[3]),
    .o(n146));  // ../RTL/core/fpu.v(128)
  AL_MUX u150 (
    .i0(n207),
    .i1(n199),
    .sel(exp_diff[3]),
    .o(n145));  // ../RTL/core/fpu.v(128)
  AL_MUX u151 (
    .i0(n206),
    .i1(n198),
    .sel(exp_diff[3]),
    .o(n144));  // ../RTL/core/fpu.v(128)
  AL_MUX u152 (
    .i0(n205),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n143));  // ../RTL/core/fpu.v(128)
  AL_MUX u153 (
    .i0(n204),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n142));  // ../RTL/core/fpu.v(128)
  AL_MUX u154 (
    .i0(n203),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n141));  // ../RTL/core/fpu.v(128)
  AL_MUX u155 (
    .i0(n202),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n140));  // ../RTL/core/fpu.v(128)
  AL_MUX u156 (
    .i0(n201),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n139));  // ../RTL/core/fpu.v(128)
  AL_MUX u157 (
    .i0(n200),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n138));  // ../RTL/core/fpu.v(128)
  AL_MUX u158 (
    .i0(n199),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n137));  // ../RTL/core/fpu.v(128)
  AL_MUX u159 (
    .i0(n198),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n136));  // ../RTL/core/fpu.v(128)
  AL_MUX u160 (
    .i0(n197),
    .i1(n143),
    .sel(exp_diff[4]),
    .o(n135));  // ../RTL/core/fpu.v(128)
  AL_MUX u161 (
    .i0(n158),
    .i1(n142),
    .sel(exp_diff[4]),
    .o(n194));  // ../RTL/core/fpu.v(128)
  AL_MUX u162 (
    .i0(n157),
    .i1(n141),
    .sel(exp_diff[4]),
    .o(n193));  // ../RTL/core/fpu.v(128)
  AL_MUX u163 (
    .i0(n156),
    .i1(n140),
    .sel(exp_diff[4]),
    .o(n192));  // ../RTL/core/fpu.v(128)
  AL_MUX u164 (
    .i0(n155),
    .i1(n139),
    .sel(exp_diff[4]),
    .o(n191));  // ../RTL/core/fpu.v(128)
  AL_MUX u165 (
    .i0(n154),
    .i1(n138),
    .sel(exp_diff[4]),
    .o(n190));  // ../RTL/core/fpu.v(128)
  AL_MUX u166 (
    .i0(n153),
    .i1(n137),
    .sel(exp_diff[4]),
    .o(n189));  // ../RTL/core/fpu.v(128)
  AL_MUX u167 (
    .i0(n152),
    .i1(n136),
    .sel(exp_diff[4]),
    .o(n188));  // ../RTL/core/fpu.v(128)
  and u18 (n196, real_oper, n160);  // ../RTL/core/fpu.v(151)
  or u184 (n171, exp_diff[6], exp_diff[7]);  // ../RTL/core/fpu.v(128)
  or u185 (n110, exp_diff[5], n171);  // ../RTL/core/fpu.v(128)
  AL_MUX u186 (
    .i0(n135),
    .i1(1'b0),
    .sel(n110),
    .o(n62[0]));  // ../RTL/core/fpu.v(128)
  AL_MUX u187 (
    .i0(n194),
    .i1(1'b0),
    .sel(n110),
    .o(n62[1]));  // ../RTL/core/fpu.v(128)
  AL_MUX u188 (
    .i0(n193),
    .i1(1'b0),
    .sel(n110),
    .o(n62[2]));  // ../RTL/core/fpu.v(128)
  AL_MUX u189 (
    .i0(n192),
    .i1(1'b0),
    .sel(n110),
    .o(n62[3]));  // ../RTL/core/fpu.v(128)
  or u19 (n244, w2, w1);  // ../RTL/core/fpu.v(143)
  AL_MUX u190 (
    .i0(n191),
    .i1(1'b0),
    .sel(n110),
    .o(n62[4]));  // ../RTL/core/fpu.v(128)
  AL_MUX u191 (
    .i0(n190),
    .i1(1'b0),
    .sel(n110),
    .o(n62[5]));  // ../RTL/core/fpu.v(128)
  AL_MUX u192 (
    .i0(n189),
    .i1(1'b0),
    .sel(n110),
    .o(n62[6]));  // ../RTL/core/fpu.v(128)
  AL_MUX u193 (
    .i0(n188),
    .i1(1'b0),
    .sel(n110),
    .o(n62[7]));  // ../RTL/core/fpu.v(128)
  AL_MUX u194 (
    .i0(1'b0),
    .i1(n151),
    .sel(u194_sel_is_0_o),
    .o(n62[8]));
  and u194_sel_is_0 (u194_sel_is_0_o, n110_neg, \exp_diff[4]_neg );
  AL_MUX u195 (
    .i0(1'b0),
    .i1(n150),
    .sel(u194_sel_is_0_o),
    .o(n62[9]));
  AL_MUX u196 (
    .i0(1'b0),
    .i1(n149),
    .sel(u194_sel_is_0_o),
    .o(n62[10]));
  AL_MUX u197 (
    .i0(1'b0),
    .i1(n148),
    .sel(u194_sel_is_0_o),
    .o(n62[11]));
  AL_MUX u198 (
    .i0(1'b0),
    .i1(n147),
    .sel(u194_sel_is_0_o),
    .o(n62[12]));
  AL_MUX u199 (
    .i0(1'b0),
    .i1(n146),
    .sel(u194_sel_is_0_o),
    .o(n62[13]));
  AL_MUX u200 (
    .i0(1'b0),
    .i1(n145),
    .sel(u194_sel_is_0_o),
    .o(n62[14]));
  AL_MUX u201 (
    .i0(1'b0),
    .i1(n144),
    .sel(u194_sel_is_0_o),
    .o(n62[15]));
  AL_MUX u202 (
    .i0(1'b0),
    .i1(n143),
    .sel(u194_sel_is_0_o),
    .o(n62[16]));
  AL_MUX u203 (
    .i0(1'b0),
    .i1(n142),
    .sel(u194_sel_is_0_o),
    .o(n62[17]));
  AL_MUX u204 (
    .i0(1'b0),
    .i1(n141),
    .sel(u194_sel_is_0_o),
    .o(n62[18]));
  AL_MUX u205 (
    .i0(1'b0),
    .i1(n140),
    .sel(u194_sel_is_0_o),
    .o(n62[19]));
  AL_MUX u206 (
    .i0(1'b0),
    .i1(n139),
    .sel(u194_sel_is_0_o),
    .o(n62[20]));
  AL_MUX u207 (
    .i0(1'b0),
    .i1(n138),
    .sel(u194_sel_is_0_o),
    .o(n62[21]));
  AL_MUX u208 (
    .i0(1'b0),
    .i1(n137),
    .sel(u194_sel_is_0_o),
    .o(n62[22]));
  AL_MUX u209 (
    .i0(1'b0),
    .i1(n136),
    .sel(u194_sel_is_0_o),
    .o(n62[23]));
  AL_MUX u210 (
    .i0(n1[1]),
    .i1(n1[2]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n108));  // ../RTL/core/fpu.v(127)
  AL_MUX u211 (
    .i0(n1[2]),
    .i1(n1[3]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n107));  // ../RTL/core/fpu.v(127)
  AL_MUX u212 (
    .i0(n1[3]),
    .i1(n1[4]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n106));  // ../RTL/core/fpu.v(127)
  AL_MUX u213 (
    .i0(n1[4]),
    .i1(n1[5]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n105));  // ../RTL/core/fpu.v(127)
  AL_MUX u214 (
    .i0(n1[5]),
    .i1(n1[6]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n104));  // ../RTL/core/fpu.v(127)
  AL_MUX u215 (
    .i0(n1[6]),
    .i1(n1[7]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n103));  // ../RTL/core/fpu.v(127)
  AL_MUX u216 (
    .i0(n1[7]),
    .i1(n1[8]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n102));  // ../RTL/core/fpu.v(127)
  AL_MUX u217 (
    .i0(n1[8]),
    .i1(n1[9]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n101));  // ../RTL/core/fpu.v(127)
  AL_MUX u218 (
    .i0(n1[9]),
    .i1(n1[10]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n100));  // ../RTL/core/fpu.v(127)
  AL_MUX u219 (
    .i0(n1[10]),
    .i1(n1[11]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n99));  // ../RTL/core/fpu.v(127)
  AL_MUX u220 (
    .i0(n1[11]),
    .i1(n1[12]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n98));  // ../RTL/core/fpu.v(127)
  AL_MUX u221 (
    .i0(n1[12]),
    .i1(n1[13]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n97));  // ../RTL/core/fpu.v(127)
  AL_MUX u222 (
    .i0(n1[13]),
    .i1(n1[14]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n96));  // ../RTL/core/fpu.v(127)
  AL_MUX u223 (
    .i0(n1[14]),
    .i1(n1[15]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n95));  // ../RTL/core/fpu.v(127)
  AL_MUX u224 (
    .i0(n1[15]),
    .i1(n1[16]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n94));  // ../RTL/core/fpu.v(127)
  AL_MUX u225 (
    .i0(n1[16]),
    .i1(n1[17]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n93));  // ../RTL/core/fpu.v(127)
  AL_MUX u226 (
    .i0(n1[17]),
    .i1(n1[18]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n92));  // ../RTL/core/fpu.v(127)
  AL_MUX u227 (
    .i0(n1[18]),
    .i1(n1[19]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n91));  // ../RTL/core/fpu.v(127)
  AL_MUX u228 (
    .i0(n1[19]),
    .i1(n1[20]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n90));  // ../RTL/core/fpu.v(127)
  AL_MUX u229 (
    .i0(n1[20]),
    .i1(n1[21]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n89));  // ../RTL/core/fpu.v(127)
  AL_MUX u230 (
    .i0(n1[21]),
    .i1(n1[22]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n88));  // ../RTL/core/fpu.v(127)
  AL_MUX u231 (
    .i0(n1[22]),
    .i1(reduced_or_E1),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n87));  // ../RTL/core/fpu.v(127)
  AL_MUX u232 (
    .i0(reduced_or_E1),
    .i1(1'b0),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n86));  // ../RTL/core/fpu.v(127)
  AL_MUX u233 (
    .i0(n109),
    .i1(n107),
    .sel(exp_diff[1]),
    .o(n85));  // ../RTL/core/fpu.v(127)
  AL_MUX u234 (
    .i0(n108),
    .i1(n106),
    .sel(exp_diff[1]),
    .o(n84));  // ../RTL/core/fpu.v(127)
  AL_MUX u235 (
    .i0(n107),
    .i1(n105),
    .sel(exp_diff[1]),
    .o(n83));  // ../RTL/core/fpu.v(127)
  AL_MUX u236 (
    .i0(n106),
    .i1(n104),
    .sel(exp_diff[1]),
    .o(n82));  // ../RTL/core/fpu.v(127)
  AL_MUX u237 (
    .i0(n105),
    .i1(n103),
    .sel(exp_diff[1]),
    .o(n81));  // ../RTL/core/fpu.v(127)
  AL_MUX u238 (
    .i0(n104),
    .i1(n102),
    .sel(exp_diff[1]),
    .o(n80));  // ../RTL/core/fpu.v(127)
  AL_MUX u239 (
    .i0(n103),
    .i1(n101),
    .sel(exp_diff[1]),
    .o(n79));  // ../RTL/core/fpu.v(127)
  AL_MUX u240 (
    .i0(n102),
    .i1(n100),
    .sel(exp_diff[1]),
    .o(n78));  // ../RTL/core/fpu.v(127)
  AL_MUX u241 (
    .i0(n101),
    .i1(n99),
    .sel(exp_diff[1]),
    .o(n77));  // ../RTL/core/fpu.v(127)
  AL_MUX u242 (
    .i0(n100),
    .i1(n98),
    .sel(exp_diff[1]),
    .o(n76));  // ../RTL/core/fpu.v(127)
  AL_MUX u243 (
    .i0(n99),
    .i1(n97),
    .sel(exp_diff[1]),
    .o(n75));  // ../RTL/core/fpu.v(127)
  AL_MUX u244 (
    .i0(n98),
    .i1(n96),
    .sel(exp_diff[1]),
    .o(n74));  // ../RTL/core/fpu.v(127)
  AL_MUX u245 (
    .i0(n97),
    .i1(n95),
    .sel(exp_diff[1]),
    .o(n73));  // ../RTL/core/fpu.v(127)
  AL_MUX u246 (
    .i0(n96),
    .i1(n94),
    .sel(exp_diff[1]),
    .o(n72));  // ../RTL/core/fpu.v(127)
  AL_MUX u247 (
    .i0(n95),
    .i1(n93),
    .sel(exp_diff[1]),
    .o(n71));  // ../RTL/core/fpu.v(127)
  AL_MUX u248 (
    .i0(n94),
    .i1(n92),
    .sel(exp_diff[1]),
    .o(n70));  // ../RTL/core/fpu.v(127)
  AL_MUX u249 (
    .i0(n93),
    .i1(n91),
    .sel(exp_diff[1]),
    .o(n69));  // ../RTL/core/fpu.v(127)
  AL_MUX u250 (
    .i0(n92),
    .i1(n90),
    .sel(exp_diff[1]),
    .o(n68));  // ../RTL/core/fpu.v(127)
  AL_MUX u251 (
    .i0(n91),
    .i1(n89),
    .sel(exp_diff[1]),
    .o(n67));  // ../RTL/core/fpu.v(127)
  AL_MUX u252 (
    .i0(n90),
    .i1(n88),
    .sel(exp_diff[1]),
    .o(n66));  // ../RTL/core/fpu.v(127)
  AL_MUX u253 (
    .i0(n89),
    .i1(n87),
    .sel(exp_diff[1]),
    .o(n65));  // ../RTL/core/fpu.v(127)
  AL_MUX u254 (
    .i0(n88),
    .i1(n86),
    .sel(exp_diff[1]),
    .o(n64));  // ../RTL/core/fpu.v(127)
  AL_MUX u255 (
    .i0(n87),
    .i1(1'b0),
    .sel(exp_diff[1]),
    .o(n63));  // ../RTL/core/fpu.v(127)
  AL_MUX u257 (
    .i0(n85),
    .i1(n81),
    .sel(exp_diff[2]),
    .o(n60));  // ../RTL/core/fpu.v(127)
  AL_MUX u258 (
    .i0(n84),
    .i1(n80),
    .sel(exp_diff[2]),
    .o(n59));  // ../RTL/core/fpu.v(127)
  AL_MUX u259 (
    .i0(n83),
    .i1(n79),
    .sel(exp_diff[2]),
    .o(n58));  // ../RTL/core/fpu.v(127)
  AL_MUX u260 (
    .i0(n82),
    .i1(n78),
    .sel(exp_diff[2]),
    .o(n57));  // ../RTL/core/fpu.v(127)
  AL_MUX u261 (
    .i0(n81),
    .i1(n77),
    .sel(exp_diff[2]),
    .o(n56));  // ../RTL/core/fpu.v(127)
  AL_MUX u262 (
    .i0(n80),
    .i1(n76),
    .sel(exp_diff[2]),
    .o(n55));  // ../RTL/core/fpu.v(127)
  AL_MUX u263 (
    .i0(n79),
    .i1(n75),
    .sel(exp_diff[2]),
    .o(n54));  // ../RTL/core/fpu.v(127)
  AL_MUX u264 (
    .i0(n78),
    .i1(n74),
    .sel(exp_diff[2]),
    .o(n53));  // ../RTL/core/fpu.v(127)
  AL_MUX u265 (
    .i0(n77),
    .i1(n73),
    .sel(exp_diff[2]),
    .o(n52));  // ../RTL/core/fpu.v(127)
  AL_MUX u266 (
    .i0(n76),
    .i1(n72),
    .sel(exp_diff[2]),
    .o(n51));  // ../RTL/core/fpu.v(127)
  AL_MUX u267 (
    .i0(n75),
    .i1(n71),
    .sel(exp_diff[2]),
    .o(n50));  // ../RTL/core/fpu.v(127)
  AL_MUX u268 (
    .i0(n74),
    .i1(n70),
    .sel(exp_diff[2]),
    .o(n49));  // ../RTL/core/fpu.v(127)
  AL_MUX u269 (
    .i0(n73),
    .i1(n69),
    .sel(exp_diff[2]),
    .o(n48));  // ../RTL/core/fpu.v(127)
  AL_MUX u270 (
    .i0(n72),
    .i1(n68),
    .sel(exp_diff[2]),
    .o(n47));  // ../RTL/core/fpu.v(127)
  AL_MUX u271 (
    .i0(n71),
    .i1(n67),
    .sel(exp_diff[2]),
    .o(n46));  // ../RTL/core/fpu.v(127)
  AL_MUX u272 (
    .i0(n70),
    .i1(n66),
    .sel(exp_diff[2]),
    .o(n45));  // ../RTL/core/fpu.v(127)
  AL_MUX u273 (
    .i0(n69),
    .i1(n65),
    .sel(exp_diff[2]),
    .o(n44));  // ../RTL/core/fpu.v(127)
  AL_MUX u274 (
    .i0(n68),
    .i1(n64),
    .sel(exp_diff[2]),
    .o(n43));  // ../RTL/core/fpu.v(127)
  AL_MUX u275 (
    .i0(n67),
    .i1(n63),
    .sel(exp_diff[2]),
    .o(n42));  // ../RTL/core/fpu.v(127)
  AL_MUX u276 (
    .i0(n66),
    .i1(n112),
    .sel(exp_diff[2]),
    .o(n41));  // ../RTL/core/fpu.v(127)
  AL_MUX u277 (
    .i0(n65),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n40));  // ../RTL/core/fpu.v(127)
  AL_MUX u278 (
    .i0(n64),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n39));  // ../RTL/core/fpu.v(127)
  AL_MUX u279 (
    .i0(n63),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n38));  // ../RTL/core/fpu.v(127)
  AL_MUX u281 (
    .i0(n60),
    .i1(n52),
    .sel(exp_diff[3]),
    .o(n263));  // ../RTL/core/fpu.v(127)
  AL_MUX u282 (
    .i0(n59),
    .i1(n51),
    .sel(exp_diff[3]),
    .o(n262));  // ../RTL/core/fpu.v(127)
  AL_MUX u283 (
    .i0(n58),
    .i1(n50),
    .sel(exp_diff[3]),
    .o(n261));  // ../RTL/core/fpu.v(127)
  AL_MUX u284 (
    .i0(n57),
    .i1(n49),
    .sel(exp_diff[3]),
    .o(n260));  // ../RTL/core/fpu.v(127)
  AL_MUX u285 (
    .i0(n56),
    .i1(n48),
    .sel(exp_diff[3]),
    .o(n259));  // ../RTL/core/fpu.v(127)
  AL_MUX u286 (
    .i0(n55),
    .i1(n47),
    .sel(exp_diff[3]),
    .o(n258));  // ../RTL/core/fpu.v(127)
  AL_MUX u287 (
    .i0(n54),
    .i1(n46),
    .sel(exp_diff[3]),
    .o(n257));  // ../RTL/core/fpu.v(127)
  AL_MUX u288 (
    .i0(n53),
    .i1(n45),
    .sel(exp_diff[3]),
    .o(n265));  // ../RTL/core/fpu.v(127)
  AL_MUX u289 (
    .i0(n52),
    .i1(n44),
    .sel(exp_diff[3]),
    .o(n256));  // ../RTL/core/fpu.v(127)
  AL_MUX u290 (
    .i0(n51),
    .i1(n43),
    .sel(exp_diff[3]),
    .o(n255));  // ../RTL/core/fpu.v(127)
  AL_MUX u291 (
    .i0(n50),
    .i1(n42),
    .sel(exp_diff[3]),
    .o(n254));  // ../RTL/core/fpu.v(127)
  AL_MUX u292 (
    .i0(n49),
    .i1(n41),
    .sel(exp_diff[3]),
    .o(n253));  // ../RTL/core/fpu.v(127)
  AL_MUX u293 (
    .i0(n48),
    .i1(n40),
    .sel(exp_diff[3]),
    .o(n252));  // ../RTL/core/fpu.v(127)
  AL_MUX u294 (
    .i0(n47),
    .i1(n39),
    .sel(exp_diff[3]),
    .o(n251));  // ../RTL/core/fpu.v(127)
  AL_MUX u295 (
    .i0(n46),
    .i1(n38),
    .sel(exp_diff[3]),
    .o(n250));  // ../RTL/core/fpu.v(127)
  AL_MUX u296 (
    .i0(n45),
    .i1(n198),
    .sel(exp_diff[3]),
    .o(n249));  // ../RTL/core/fpu.v(127)
  AL_MUX u297 (
    .i0(n44),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n11));  // ../RTL/core/fpu.v(127)
  AL_MUX u298 (
    .i0(n43),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n10));  // ../RTL/core/fpu.v(127)
  AL_MUX u299 (
    .i0(n42),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n9));  // ../RTL/core/fpu.v(127)
  AL_MUX u300 (
    .i0(n41),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n8));  // ../RTL/core/fpu.v(127)
  AL_MUX u301 (
    .i0(n40),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n7));  // ../RTL/core/fpu.v(127)
  AL_MUX u302 (
    .i0(n39),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n6));  // ../RTL/core/fpu.v(127)
  AL_MUX u303 (
    .i0(n38),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n5));  // ../RTL/core/fpu.v(127)
  AL_MUX u305 (
    .i0(n263),
    .i1(n11),
    .sel(exp_diff[4]),
    .o(n36));  // ../RTL/core/fpu.v(127)
  AL_MUX u306 (
    .i0(n262),
    .i1(n10),
    .sel(exp_diff[4]),
    .o(n35));  // ../RTL/core/fpu.v(127)
  AL_MUX u307 (
    .i0(n261),
    .i1(n9),
    .sel(exp_diff[4]),
    .o(n34));  // ../RTL/core/fpu.v(127)
  AL_MUX u308 (
    .i0(n260),
    .i1(n8),
    .sel(exp_diff[4]),
    .o(n33));  // ../RTL/core/fpu.v(127)
  AL_MUX u309 (
    .i0(n259),
    .i1(n7),
    .sel(exp_diff[4]),
    .o(n32));  // ../RTL/core/fpu.v(127)
  AL_MUX u310 (
    .i0(n258),
    .i1(n6),
    .sel(exp_diff[4]),
    .o(n31));  // ../RTL/core/fpu.v(127)
  AL_MUX u311 (
    .i0(n257),
    .i1(n5),
    .sel(exp_diff[4]),
    .o(n30));  // ../RTL/core/fpu.v(127)
  AL_MUX u312 (
    .i0(n265),
    .i1(n136),
    .sel(exp_diff[4]),
    .o(n29));  // ../RTL/core/fpu.v(127)
  AL_MUX u331 (
    .i0(n36),
    .i1(1'b0),
    .sel(n110),
    .o(n37[0]));  // ../RTL/core/fpu.v(127)
  AL_MUX u332 (
    .i0(n35),
    .i1(1'b0),
    .sel(n110),
    .o(n37[1]));  // ../RTL/core/fpu.v(127)
  AL_MUX u333 (
    .i0(n34),
    .i1(1'b0),
    .sel(n110),
    .o(n37[2]));  // ../RTL/core/fpu.v(127)
  AL_MUX u334 (
    .i0(n33),
    .i1(1'b0),
    .sel(n110),
    .o(n37[3]));  // ../RTL/core/fpu.v(127)
  AL_MUX u335 (
    .i0(n32),
    .i1(1'b0),
    .sel(n110),
    .o(n37[4]));  // ../RTL/core/fpu.v(127)
  AL_MUX u336 (
    .i0(n31),
    .i1(1'b0),
    .sel(n110),
    .o(n37[5]));  // ../RTL/core/fpu.v(127)
  AL_MUX u337 (
    .i0(n30),
    .i1(1'b0),
    .sel(n110),
    .o(n37[6]));  // ../RTL/core/fpu.v(127)
  AL_MUX u338 (
    .i0(n29),
    .i1(1'b0),
    .sel(n110),
    .o(n37[7]));  // ../RTL/core/fpu.v(127)
  AL_MUX u339 (
    .i0(1'b0),
    .i1(n256),
    .sel(u194_sel_is_0_o),
    .o(n37[8]));
  AL_MUX u340 (
    .i0(1'b0),
    .i1(n255),
    .sel(u194_sel_is_0_o),
    .o(n37[9]));
  AL_MUX u341 (
    .i0(1'b0),
    .i1(n254),
    .sel(u194_sel_is_0_o),
    .o(n37[10]));
  AL_MUX u342 (
    .i0(1'b0),
    .i1(n253),
    .sel(u194_sel_is_0_o),
    .o(n37[11]));
  AL_MUX u343 (
    .i0(1'b0),
    .i1(n252),
    .sel(u194_sel_is_0_o),
    .o(n37[12]));
  AL_MUX u344 (
    .i0(1'b0),
    .i1(n251),
    .sel(u194_sel_is_0_o),
    .o(n37[13]));
  AL_MUX u345 (
    .i0(1'b0),
    .i1(n250),
    .sel(u194_sel_is_0_o),
    .o(n37[14]));
  AL_MUX u346 (
    .i0(1'b0),
    .i1(n249),
    .sel(u194_sel_is_0_o),
    .o(n37[15]));
  AL_MUX u347 (
    .i0(1'b0),
    .i1(n11),
    .sel(u194_sel_is_0_o),
    .o(n37[16]));
  AL_MUX u348 (
    .i0(1'b0),
    .i1(n10),
    .sel(u194_sel_is_0_o),
    .o(n37[17]));
  AL_MUX u349 (
    .i0(1'b0),
    .i1(n9),
    .sel(u194_sel_is_0_o),
    .o(n37[18]));
  AL_MUX u350 (
    .i0(1'b0),
    .i1(n8),
    .sel(u194_sel_is_0_o),
    .o(n37[19]));
  AL_MUX u351 (
    .i0(1'b0),
    .i1(n7),
    .sel(u194_sel_is_0_o),
    .o(n37[20]));
  AL_MUX u352 (
    .i0(1'b0),
    .i1(n6),
    .sel(u194_sel_is_0_o),
    .o(n37[21]));
  AL_MUX u353 (
    .i0(1'b0),
    .i1(n5),
    .sel(u194_sel_is_0_o),
    .o(n37[22]));
  AL_MUX u5 (
    .i0(n1[0]),
    .i1(n1[1]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n109));  // ../RTL/core/fpu.v(127)
  AL_MUX u6 (
    .i0(n2[0]),
    .i1(n2[1]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n241));  // ../RTL/core/fpu.v(128)
  or u62 (result[31], w3, n244);  // ../RTL/core/fpu.v(143)
  and u63 (w1, n160, n243);  // ../RTL/core/fpu.v(140)
  xor u64 (real_oper, n2[31], n1[31]);  // ../RTL/core/fpu.v(131)
  AL_MUX u65 (
    .i0(n2[1]),
    .i1(n2[2]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n240));  // ../RTL/core/fpu.v(128)
  AL_MUX u66 (
    .i0(n2[2]),
    .i1(n2[3]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n239));  // ../RTL/core/fpu.v(128)
  AL_MUX u67 (
    .i0(n2[3]),
    .i1(n2[4]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n238));  // ../RTL/core/fpu.v(128)
  AL_MUX u68 (
    .i0(n2[4]),
    .i1(n2[5]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n237));  // ../RTL/core/fpu.v(128)
  AL_MUX u69 (
    .i0(n2[5]),
    .i1(n2[6]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n236));  // ../RTL/core/fpu.v(128)
  AL_MUX u70 (
    .i0(n2[6]),
    .i1(n2[7]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n235));  // ../RTL/core/fpu.v(128)
  AL_MUX u71 (
    .i0(n2[7]),
    .i1(n2[8]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n234));  // ../RTL/core/fpu.v(128)
  AL_MUX u72 (
    .i0(n2[8]),
    .i1(n2[9]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n233));  // ../RTL/core/fpu.v(128)
  AL_MUX u73 (
    .i0(n2[9]),
    .i1(n2[10]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n232));  // ../RTL/core/fpu.v(128)
  AL_MUX u74 (
    .i0(n2[10]),
    .i1(n2[11]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n231));  // ../RTL/core/fpu.v(128)
  AL_MUX u75 (
    .i0(n2[11]),
    .i1(n2[12]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n230));  // ../RTL/core/fpu.v(128)
  AL_MUX u76 (
    .i0(n2[12]),
    .i1(n2[13]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n229));  // ../RTL/core/fpu.v(128)
  AL_MUX u77 (
    .i0(n2[13]),
    .i1(n2[14]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n228));  // ../RTL/core/fpu.v(128)
  AL_MUX u78 (
    .i0(n2[14]),
    .i1(n2[15]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n227));  // ../RTL/core/fpu.v(128)
  AL_MUX u79 (
    .i0(n2[15]),
    .i1(n2[16]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n226));  // ../RTL/core/fpu.v(128)
  not u8 (n159, n1[31]);  // ../RTL/core/fpu.v(140)
  AL_MUX u80 (
    .i0(n2[16]),
    .i1(n2[17]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n225));  // ../RTL/core/fpu.v(128)
  AL_MUX u81 (
    .i0(n2[17]),
    .i1(n2[18]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n224));  // ../RTL/core/fpu.v(128)
  AL_MUX u82 (
    .i0(n2[18]),
    .i1(n2[19]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n223));  // ../RTL/core/fpu.v(128)
  AL_MUX u83 (
    .i0(n2[19]),
    .i1(n2[20]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n222));  // ../RTL/core/fpu.v(128)
  AL_MUX u84 (
    .i0(n2[20]),
    .i1(n2[21]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n221));  // ../RTL/core/fpu.v(128)
  AL_MUX u85 (
    .i0(n2[21]),
    .i1(n2[22]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n165));  // ../RTL/core/fpu.v(128)
  AL_MUX u86 (
    .i0(n2[22]),
    .i1(reduced_or_E1),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n164));  // ../RTL/core/fpu.v(128)
  AL_MUX u88 (
    .i0(n241),
    .i1(n239),
    .sel(exp_diff[1]),
    .o(n161));  // ../RTL/core/fpu.v(128)
  AL_MUX u89 (
    .i0(n240),
    .i1(n238),
    .sel(exp_diff[1]),
    .o(n134));  // ../RTL/core/fpu.v(128)
  not u9 (n160, M_carry);  // ../RTL/core/fpu.v(140)
  AL_MUX u90 (
    .i0(n239),
    .i1(n237),
    .sel(exp_diff[1]),
    .o(n133));  // ../RTL/core/fpu.v(128)
  AL_MUX u91 (
    .i0(n238),
    .i1(n236),
    .sel(exp_diff[1]),
    .o(n132));  // ../RTL/core/fpu.v(128)
  AL_MUX u92 (
    .i0(n237),
    .i1(n235),
    .sel(exp_diff[1]),
    .o(n131));  // ../RTL/core/fpu.v(128)
  AL_MUX u93 (
    .i0(n236),
    .i1(n234),
    .sel(exp_diff[1]),
    .o(n130));  // ../RTL/core/fpu.v(128)
  AL_MUX u94 (
    .i0(n235),
    .i1(n233),
    .sel(exp_diff[1]),
    .o(n129));  // ../RTL/core/fpu.v(128)
  AL_MUX u95 (
    .i0(n234),
    .i1(n232),
    .sel(exp_diff[1]),
    .o(n128));  // ../RTL/core/fpu.v(128)
  AL_MUX u96 (
    .i0(n233),
    .i1(n231),
    .sel(exp_diff[1]),
    .o(n127));  // ../RTL/core/fpu.v(128)
  AL_MUX u97 (
    .i0(n232),
    .i1(n230),
    .sel(exp_diff[1]),
    .o(n126));  // ../RTL/core/fpu.v(128)
  AL_MUX u98 (
    .i0(n231),
    .i1(n229),
    .sel(exp_diff[1]),
    .o(n125));  // ../RTL/core/fpu.v(128)
  AL_MUX u99 (
    .i0(n230),
    .i1(n228),
    .sel(exp_diff[1]),
    .o(n124));  // ../RTL/core/fpu.v(128)

endmodule 

module mult_u24_u24_o48
  (
  i0,
  i1,
  o
  );

  input [23:0] i0;
  input [23:0] i1;
  output [47:0] o;

  wire [23:0] and_0;
  wire [23:0] and_1;
  wire [23:0] and_10;
  wire [23:0] and_11;
  wire [23:0] and_12;
  wire [23:0] and_13;
  wire [23:0] and_14;
  wire [23:0] and_15;
  wire [23:0] and_16;
  wire [23:0] and_17;
  wire [23:0] and_18;
  wire [23:0] and_19;
  wire [23:0] and_2;
  wire [23:0] and_20;
  wire [23:0] and_21;
  wire [23:0] and_22;
  wire [23:0] and_23;
  wire [23:0] and_3;
  wire [23:0] and_4;
  wire [23:0] and_5;
  wire [23:0] and_6;
  wire [23:0] and_7;
  wire [23:0] and_8;
  wire [23:0] and_9;
  wire [23:0] nand_0;
  wire [23:0] nand_1;
  wire [23:0] nand_10;
  wire [23:0] nand_11;
  wire [23:0] nand_12;
  wire [23:0] nand_13;
  wire [23:0] nand_14;
  wire [23:0] nand_15;
  wire [23:0] nand_16;
  wire [23:0] nand_17;
  wire [23:0] nand_18;
  wire [23:0] nand_19;
  wire [23:0] nand_2;
  wire [23:0] nand_20;
  wire [23:0] nand_21;
  wire [23:0] nand_22;
  wire [23:0] nand_23;
  wire [23:0] nand_3;
  wire [23:0] nand_4;
  wire [23:0] nand_5;
  wire [23:0] nand_6;
  wire [23:0] nand_7;
  wire [23:0] nand_8;
  wire [23:0] nand_9;

  and and_a0_b0 (and_0[0], i0[0], i1[0]);
  and and_a0_b1 (and_1[0], i0[0], i1[1]);
  and and_a0_b10 (and_10[0], i0[0], i1[10]);
  and and_a0_b11 (and_11[0], i0[0], i1[11]);
  and and_a0_b12 (and_12[0], i0[0], i1[12]);
  and and_a0_b13 (and_13[0], i0[0], i1[13]);
  and and_a0_b14 (and_14[0], i0[0], i1[14]);
  and and_a0_b15 (and_15[0], i0[0], i1[15]);
  and and_a0_b16 (and_16[0], i0[0], i1[16]);
  and and_a0_b17 (and_17[0], i0[0], i1[17]);
  and and_a0_b18 (and_18[0], i0[0], i1[18]);
  and and_a0_b19 (and_19[0], i0[0], i1[19]);
  and and_a0_b2 (and_2[0], i0[0], i1[2]);
  and and_a0_b20 (and_20[0], i0[0], i1[20]);
  and and_a0_b21 (and_21[0], i0[0], i1[21]);
  and and_a0_b22 (and_22[0], i0[0], i1[22]);
  and and_a0_b23 (and_23[0], i0[0], i1[23]);
  and and_a0_b3 (and_3[0], i0[0], i1[3]);
  and and_a0_b4 (and_4[0], i0[0], i1[4]);
  and and_a0_b5 (and_5[0], i0[0], i1[5]);
  and and_a0_b6 (and_6[0], i0[0], i1[6]);
  and and_a0_b7 (and_7[0], i0[0], i1[7]);
  and and_a0_b8 (and_8[0], i0[0], i1[8]);
  and and_a0_b9 (and_9[0], i0[0], i1[9]);
  and and_a10_b0 (and_0[10], i0[10], i1[0]);
  and and_a10_b1 (and_1[10], i0[10], i1[1]);
  and and_a10_b10 (and_10[10], i0[10], i1[10]);
  and and_a10_b11 (and_11[10], i0[10], i1[11]);
  and and_a10_b12 (and_12[10], i0[10], i1[12]);
  and and_a10_b13 (and_13[10], i0[10], i1[13]);
  and and_a10_b14 (and_14[10], i0[10], i1[14]);
  and and_a10_b15 (and_15[10], i0[10], i1[15]);
  and and_a10_b16 (and_16[10], i0[10], i1[16]);
  and and_a10_b17 (and_17[10], i0[10], i1[17]);
  and and_a10_b18 (and_18[10], i0[10], i1[18]);
  and and_a10_b19 (and_19[10], i0[10], i1[19]);
  and and_a10_b2 (and_2[10], i0[10], i1[2]);
  and and_a10_b20 (and_20[10], i0[10], i1[20]);
  and and_a10_b21 (and_21[10], i0[10], i1[21]);
  and and_a10_b22 (and_22[10], i0[10], i1[22]);
  and and_a10_b23 (and_23[10], i0[10], i1[23]);
  and and_a10_b3 (and_3[10], i0[10], i1[3]);
  and and_a10_b4 (and_4[10], i0[10], i1[4]);
  and and_a10_b5 (and_5[10], i0[10], i1[5]);
  and and_a10_b6 (and_6[10], i0[10], i1[6]);
  and and_a10_b7 (and_7[10], i0[10], i1[7]);
  and and_a10_b8 (and_8[10], i0[10], i1[8]);
  and and_a10_b9 (and_9[10], i0[10], i1[9]);
  and and_a11_b0 (and_0[11], i0[11], i1[0]);
  and and_a11_b1 (and_1[11], i0[11], i1[1]);
  and and_a11_b10 (and_10[11], i0[11], i1[10]);
  and and_a11_b11 (and_11[11], i0[11], i1[11]);
  and and_a11_b12 (and_12[11], i0[11], i1[12]);
  and and_a11_b13 (and_13[11], i0[11], i1[13]);
  and and_a11_b14 (and_14[11], i0[11], i1[14]);
  and and_a11_b15 (and_15[11], i0[11], i1[15]);
  and and_a11_b16 (and_16[11], i0[11], i1[16]);
  and and_a11_b17 (and_17[11], i0[11], i1[17]);
  and and_a11_b18 (and_18[11], i0[11], i1[18]);
  and and_a11_b19 (and_19[11], i0[11], i1[19]);
  and and_a11_b2 (and_2[11], i0[11], i1[2]);
  and and_a11_b20 (and_20[11], i0[11], i1[20]);
  and and_a11_b21 (and_21[11], i0[11], i1[21]);
  and and_a11_b22 (and_22[11], i0[11], i1[22]);
  and and_a11_b23 (and_23[11], i0[11], i1[23]);
  and and_a11_b3 (and_3[11], i0[11], i1[3]);
  and and_a11_b4 (and_4[11], i0[11], i1[4]);
  and and_a11_b5 (and_5[11], i0[11], i1[5]);
  and and_a11_b6 (and_6[11], i0[11], i1[6]);
  and and_a11_b7 (and_7[11], i0[11], i1[7]);
  and and_a11_b8 (and_8[11], i0[11], i1[8]);
  and and_a11_b9 (and_9[11], i0[11], i1[9]);
  and and_a12_b0 (and_0[12], i0[12], i1[0]);
  and and_a12_b1 (and_1[12], i0[12], i1[1]);
  and and_a12_b10 (and_10[12], i0[12], i1[10]);
  and and_a12_b11 (and_11[12], i0[12], i1[11]);
  and and_a12_b12 (and_12[12], i0[12], i1[12]);
  and and_a12_b13 (and_13[12], i0[12], i1[13]);
  and and_a12_b14 (and_14[12], i0[12], i1[14]);
  and and_a12_b15 (and_15[12], i0[12], i1[15]);
  and and_a12_b16 (and_16[12], i0[12], i1[16]);
  and and_a12_b17 (and_17[12], i0[12], i1[17]);
  and and_a12_b18 (and_18[12], i0[12], i1[18]);
  and and_a12_b19 (and_19[12], i0[12], i1[19]);
  and and_a12_b2 (and_2[12], i0[12], i1[2]);
  and and_a12_b20 (and_20[12], i0[12], i1[20]);
  and and_a12_b21 (and_21[12], i0[12], i1[21]);
  and and_a12_b22 (and_22[12], i0[12], i1[22]);
  and and_a12_b23 (and_23[12], i0[12], i1[23]);
  and and_a12_b3 (and_3[12], i0[12], i1[3]);
  and and_a12_b4 (and_4[12], i0[12], i1[4]);
  and and_a12_b5 (and_5[12], i0[12], i1[5]);
  and and_a12_b6 (and_6[12], i0[12], i1[6]);
  and and_a12_b7 (and_7[12], i0[12], i1[7]);
  and and_a12_b8 (and_8[12], i0[12], i1[8]);
  and and_a12_b9 (and_9[12], i0[12], i1[9]);
  and and_a13_b0 (and_0[13], i0[13], i1[0]);
  and and_a13_b1 (and_1[13], i0[13], i1[1]);
  and and_a13_b10 (and_10[13], i0[13], i1[10]);
  and and_a13_b11 (and_11[13], i0[13], i1[11]);
  and and_a13_b12 (and_12[13], i0[13], i1[12]);
  and and_a13_b13 (and_13[13], i0[13], i1[13]);
  and and_a13_b14 (and_14[13], i0[13], i1[14]);
  and and_a13_b15 (and_15[13], i0[13], i1[15]);
  and and_a13_b16 (and_16[13], i0[13], i1[16]);
  and and_a13_b17 (and_17[13], i0[13], i1[17]);
  and and_a13_b18 (and_18[13], i0[13], i1[18]);
  and and_a13_b19 (and_19[13], i0[13], i1[19]);
  and and_a13_b2 (and_2[13], i0[13], i1[2]);
  and and_a13_b20 (and_20[13], i0[13], i1[20]);
  and and_a13_b21 (and_21[13], i0[13], i1[21]);
  and and_a13_b22 (and_22[13], i0[13], i1[22]);
  and and_a13_b23 (and_23[13], i0[13], i1[23]);
  and and_a13_b3 (and_3[13], i0[13], i1[3]);
  and and_a13_b4 (and_4[13], i0[13], i1[4]);
  and and_a13_b5 (and_5[13], i0[13], i1[5]);
  and and_a13_b6 (and_6[13], i0[13], i1[6]);
  and and_a13_b7 (and_7[13], i0[13], i1[7]);
  and and_a13_b8 (and_8[13], i0[13], i1[8]);
  and and_a13_b9 (and_9[13], i0[13], i1[9]);
  and and_a14_b0 (and_0[14], i0[14], i1[0]);
  and and_a14_b1 (and_1[14], i0[14], i1[1]);
  and and_a14_b10 (and_10[14], i0[14], i1[10]);
  and and_a14_b11 (and_11[14], i0[14], i1[11]);
  and and_a14_b12 (and_12[14], i0[14], i1[12]);
  and and_a14_b13 (and_13[14], i0[14], i1[13]);
  and and_a14_b14 (and_14[14], i0[14], i1[14]);
  and and_a14_b15 (and_15[14], i0[14], i1[15]);
  and and_a14_b16 (and_16[14], i0[14], i1[16]);
  and and_a14_b17 (and_17[14], i0[14], i1[17]);
  and and_a14_b18 (and_18[14], i0[14], i1[18]);
  and and_a14_b19 (and_19[14], i0[14], i1[19]);
  and and_a14_b2 (and_2[14], i0[14], i1[2]);
  and and_a14_b20 (and_20[14], i0[14], i1[20]);
  and and_a14_b21 (and_21[14], i0[14], i1[21]);
  and and_a14_b22 (and_22[14], i0[14], i1[22]);
  and and_a14_b23 (and_23[14], i0[14], i1[23]);
  and and_a14_b3 (and_3[14], i0[14], i1[3]);
  and and_a14_b4 (and_4[14], i0[14], i1[4]);
  and and_a14_b5 (and_5[14], i0[14], i1[5]);
  and and_a14_b6 (and_6[14], i0[14], i1[6]);
  and and_a14_b7 (and_7[14], i0[14], i1[7]);
  and and_a14_b8 (and_8[14], i0[14], i1[8]);
  and and_a14_b9 (and_9[14], i0[14], i1[9]);
  and and_a15_b0 (and_0[15], i0[15], i1[0]);
  and and_a15_b1 (and_1[15], i0[15], i1[1]);
  and and_a15_b10 (and_10[15], i0[15], i1[10]);
  and and_a15_b11 (and_11[15], i0[15], i1[11]);
  and and_a15_b12 (and_12[15], i0[15], i1[12]);
  and and_a15_b13 (and_13[15], i0[15], i1[13]);
  and and_a15_b14 (and_14[15], i0[15], i1[14]);
  and and_a15_b15 (and_15[15], i0[15], i1[15]);
  and and_a15_b16 (and_16[15], i0[15], i1[16]);
  and and_a15_b17 (and_17[15], i0[15], i1[17]);
  and and_a15_b18 (and_18[15], i0[15], i1[18]);
  and and_a15_b19 (and_19[15], i0[15], i1[19]);
  and and_a15_b2 (and_2[15], i0[15], i1[2]);
  and and_a15_b20 (and_20[15], i0[15], i1[20]);
  and and_a15_b21 (and_21[15], i0[15], i1[21]);
  and and_a15_b22 (and_22[15], i0[15], i1[22]);
  and and_a15_b23 (and_23[15], i0[15], i1[23]);
  and and_a15_b3 (and_3[15], i0[15], i1[3]);
  and and_a15_b4 (and_4[15], i0[15], i1[4]);
  and and_a15_b5 (and_5[15], i0[15], i1[5]);
  and and_a15_b6 (and_6[15], i0[15], i1[6]);
  and and_a15_b7 (and_7[15], i0[15], i1[7]);
  and and_a15_b8 (and_8[15], i0[15], i1[8]);
  and and_a15_b9 (and_9[15], i0[15], i1[9]);
  and and_a16_b0 (and_0[16], i0[16], i1[0]);
  and and_a16_b1 (and_1[16], i0[16], i1[1]);
  and and_a16_b10 (and_10[16], i0[16], i1[10]);
  and and_a16_b11 (and_11[16], i0[16], i1[11]);
  and and_a16_b12 (and_12[16], i0[16], i1[12]);
  and and_a16_b13 (and_13[16], i0[16], i1[13]);
  and and_a16_b14 (and_14[16], i0[16], i1[14]);
  and and_a16_b15 (and_15[16], i0[16], i1[15]);
  and and_a16_b16 (and_16[16], i0[16], i1[16]);
  and and_a16_b17 (and_17[16], i0[16], i1[17]);
  and and_a16_b18 (and_18[16], i0[16], i1[18]);
  and and_a16_b19 (and_19[16], i0[16], i1[19]);
  and and_a16_b2 (and_2[16], i0[16], i1[2]);
  and and_a16_b20 (and_20[16], i0[16], i1[20]);
  and and_a16_b21 (and_21[16], i0[16], i1[21]);
  and and_a16_b22 (and_22[16], i0[16], i1[22]);
  and and_a16_b23 (and_23[16], i0[16], i1[23]);
  and and_a16_b3 (and_3[16], i0[16], i1[3]);
  and and_a16_b4 (and_4[16], i0[16], i1[4]);
  and and_a16_b5 (and_5[16], i0[16], i1[5]);
  and and_a16_b6 (and_6[16], i0[16], i1[6]);
  and and_a16_b7 (and_7[16], i0[16], i1[7]);
  and and_a16_b8 (and_8[16], i0[16], i1[8]);
  and and_a16_b9 (and_9[16], i0[16], i1[9]);
  and and_a17_b0 (and_0[17], i0[17], i1[0]);
  and and_a17_b1 (and_1[17], i0[17], i1[1]);
  and and_a17_b10 (and_10[17], i0[17], i1[10]);
  and and_a17_b11 (and_11[17], i0[17], i1[11]);
  and and_a17_b12 (and_12[17], i0[17], i1[12]);
  and and_a17_b13 (and_13[17], i0[17], i1[13]);
  and and_a17_b14 (and_14[17], i0[17], i1[14]);
  and and_a17_b15 (and_15[17], i0[17], i1[15]);
  and and_a17_b16 (and_16[17], i0[17], i1[16]);
  and and_a17_b17 (and_17[17], i0[17], i1[17]);
  and and_a17_b18 (and_18[17], i0[17], i1[18]);
  and and_a17_b19 (and_19[17], i0[17], i1[19]);
  and and_a17_b2 (and_2[17], i0[17], i1[2]);
  and and_a17_b20 (and_20[17], i0[17], i1[20]);
  and and_a17_b21 (and_21[17], i0[17], i1[21]);
  and and_a17_b22 (and_22[17], i0[17], i1[22]);
  and and_a17_b23 (and_23[17], i0[17], i1[23]);
  and and_a17_b3 (and_3[17], i0[17], i1[3]);
  and and_a17_b4 (and_4[17], i0[17], i1[4]);
  and and_a17_b5 (and_5[17], i0[17], i1[5]);
  and and_a17_b6 (and_6[17], i0[17], i1[6]);
  and and_a17_b7 (and_7[17], i0[17], i1[7]);
  and and_a17_b8 (and_8[17], i0[17], i1[8]);
  and and_a17_b9 (and_9[17], i0[17], i1[9]);
  and and_a18_b0 (and_0[18], i0[18], i1[0]);
  and and_a18_b1 (and_1[18], i0[18], i1[1]);
  and and_a18_b10 (and_10[18], i0[18], i1[10]);
  and and_a18_b11 (and_11[18], i0[18], i1[11]);
  and and_a18_b12 (and_12[18], i0[18], i1[12]);
  and and_a18_b13 (and_13[18], i0[18], i1[13]);
  and and_a18_b14 (and_14[18], i0[18], i1[14]);
  and and_a18_b15 (and_15[18], i0[18], i1[15]);
  and and_a18_b16 (and_16[18], i0[18], i1[16]);
  and and_a18_b17 (and_17[18], i0[18], i1[17]);
  and and_a18_b18 (and_18[18], i0[18], i1[18]);
  and and_a18_b19 (and_19[18], i0[18], i1[19]);
  and and_a18_b2 (and_2[18], i0[18], i1[2]);
  and and_a18_b20 (and_20[18], i0[18], i1[20]);
  and and_a18_b21 (and_21[18], i0[18], i1[21]);
  and and_a18_b22 (and_22[18], i0[18], i1[22]);
  and and_a18_b23 (and_23[18], i0[18], i1[23]);
  and and_a18_b3 (and_3[18], i0[18], i1[3]);
  and and_a18_b4 (and_4[18], i0[18], i1[4]);
  and and_a18_b5 (and_5[18], i0[18], i1[5]);
  and and_a18_b6 (and_6[18], i0[18], i1[6]);
  and and_a18_b7 (and_7[18], i0[18], i1[7]);
  and and_a18_b8 (and_8[18], i0[18], i1[8]);
  and and_a18_b9 (and_9[18], i0[18], i1[9]);
  and and_a19_b0 (and_0[19], i0[19], i1[0]);
  and and_a19_b1 (and_1[19], i0[19], i1[1]);
  and and_a19_b10 (and_10[19], i0[19], i1[10]);
  and and_a19_b11 (and_11[19], i0[19], i1[11]);
  and and_a19_b12 (and_12[19], i0[19], i1[12]);
  and and_a19_b13 (and_13[19], i0[19], i1[13]);
  and and_a19_b14 (and_14[19], i0[19], i1[14]);
  and and_a19_b15 (and_15[19], i0[19], i1[15]);
  and and_a19_b16 (and_16[19], i0[19], i1[16]);
  and and_a19_b17 (and_17[19], i0[19], i1[17]);
  and and_a19_b18 (and_18[19], i0[19], i1[18]);
  and and_a19_b19 (and_19[19], i0[19], i1[19]);
  and and_a19_b2 (and_2[19], i0[19], i1[2]);
  and and_a19_b20 (and_20[19], i0[19], i1[20]);
  and and_a19_b21 (and_21[19], i0[19], i1[21]);
  and and_a19_b22 (and_22[19], i0[19], i1[22]);
  and and_a19_b23 (and_23[19], i0[19], i1[23]);
  and and_a19_b3 (and_3[19], i0[19], i1[3]);
  and and_a19_b4 (and_4[19], i0[19], i1[4]);
  and and_a19_b5 (and_5[19], i0[19], i1[5]);
  and and_a19_b6 (and_6[19], i0[19], i1[6]);
  and and_a19_b7 (and_7[19], i0[19], i1[7]);
  and and_a19_b8 (and_8[19], i0[19], i1[8]);
  and and_a19_b9 (and_9[19], i0[19], i1[9]);
  and and_a1_b0 (and_0[1], i0[1], i1[0]);
  and and_a1_b1 (and_1[1], i0[1], i1[1]);
  and and_a1_b10 (and_10[1], i0[1], i1[10]);
  and and_a1_b11 (and_11[1], i0[1], i1[11]);
  and and_a1_b12 (and_12[1], i0[1], i1[12]);
  and and_a1_b13 (and_13[1], i0[1], i1[13]);
  and and_a1_b14 (and_14[1], i0[1], i1[14]);
  and and_a1_b15 (and_15[1], i0[1], i1[15]);
  and and_a1_b16 (and_16[1], i0[1], i1[16]);
  and and_a1_b17 (and_17[1], i0[1], i1[17]);
  and and_a1_b18 (and_18[1], i0[1], i1[18]);
  and and_a1_b19 (and_19[1], i0[1], i1[19]);
  and and_a1_b2 (and_2[1], i0[1], i1[2]);
  and and_a1_b20 (and_20[1], i0[1], i1[20]);
  and and_a1_b21 (and_21[1], i0[1], i1[21]);
  and and_a1_b22 (and_22[1], i0[1], i1[22]);
  and and_a1_b23 (and_23[1], i0[1], i1[23]);
  and and_a1_b3 (and_3[1], i0[1], i1[3]);
  and and_a1_b4 (and_4[1], i0[1], i1[4]);
  and and_a1_b5 (and_5[1], i0[1], i1[5]);
  and and_a1_b6 (and_6[1], i0[1], i1[6]);
  and and_a1_b7 (and_7[1], i0[1], i1[7]);
  and and_a1_b8 (and_8[1], i0[1], i1[8]);
  and and_a1_b9 (and_9[1], i0[1], i1[9]);
  and and_a20_b0 (and_0[20], i0[20], i1[0]);
  and and_a20_b1 (and_1[20], i0[20], i1[1]);
  and and_a20_b10 (and_10[20], i0[20], i1[10]);
  and and_a20_b11 (and_11[20], i0[20], i1[11]);
  and and_a20_b12 (and_12[20], i0[20], i1[12]);
  and and_a20_b13 (and_13[20], i0[20], i1[13]);
  and and_a20_b14 (and_14[20], i0[20], i1[14]);
  and and_a20_b15 (and_15[20], i0[20], i1[15]);
  and and_a20_b16 (and_16[20], i0[20], i1[16]);
  and and_a20_b17 (and_17[20], i0[20], i1[17]);
  and and_a20_b18 (and_18[20], i0[20], i1[18]);
  and and_a20_b19 (and_19[20], i0[20], i1[19]);
  and and_a20_b2 (and_2[20], i0[20], i1[2]);
  and and_a20_b20 (and_20[20], i0[20], i1[20]);
  and and_a20_b21 (and_21[20], i0[20], i1[21]);
  and and_a20_b22 (and_22[20], i0[20], i1[22]);
  and and_a20_b23 (and_23[20], i0[20], i1[23]);
  and and_a20_b3 (and_3[20], i0[20], i1[3]);
  and and_a20_b4 (and_4[20], i0[20], i1[4]);
  and and_a20_b5 (and_5[20], i0[20], i1[5]);
  and and_a20_b6 (and_6[20], i0[20], i1[6]);
  and and_a20_b7 (and_7[20], i0[20], i1[7]);
  and and_a20_b8 (and_8[20], i0[20], i1[8]);
  and and_a20_b9 (and_9[20], i0[20], i1[9]);
  and and_a21_b0 (and_0[21], i0[21], i1[0]);
  and and_a21_b1 (and_1[21], i0[21], i1[1]);
  and and_a21_b10 (and_10[21], i0[21], i1[10]);
  and and_a21_b11 (and_11[21], i0[21], i1[11]);
  and and_a21_b12 (and_12[21], i0[21], i1[12]);
  and and_a21_b13 (and_13[21], i0[21], i1[13]);
  and and_a21_b14 (and_14[21], i0[21], i1[14]);
  and and_a21_b15 (and_15[21], i0[21], i1[15]);
  and and_a21_b16 (and_16[21], i0[21], i1[16]);
  and and_a21_b17 (and_17[21], i0[21], i1[17]);
  and and_a21_b18 (and_18[21], i0[21], i1[18]);
  and and_a21_b19 (and_19[21], i0[21], i1[19]);
  and and_a21_b2 (and_2[21], i0[21], i1[2]);
  and and_a21_b20 (and_20[21], i0[21], i1[20]);
  and and_a21_b21 (and_21[21], i0[21], i1[21]);
  and and_a21_b22 (and_22[21], i0[21], i1[22]);
  and and_a21_b23 (and_23[21], i0[21], i1[23]);
  and and_a21_b3 (and_3[21], i0[21], i1[3]);
  and and_a21_b4 (and_4[21], i0[21], i1[4]);
  and and_a21_b5 (and_5[21], i0[21], i1[5]);
  and and_a21_b6 (and_6[21], i0[21], i1[6]);
  and and_a21_b7 (and_7[21], i0[21], i1[7]);
  and and_a21_b8 (and_8[21], i0[21], i1[8]);
  and and_a21_b9 (and_9[21], i0[21], i1[9]);
  and and_a22_b0 (and_0[22], i0[22], i1[0]);
  and and_a22_b1 (and_1[22], i0[22], i1[1]);
  and and_a22_b10 (and_10[22], i0[22], i1[10]);
  and and_a22_b11 (and_11[22], i0[22], i1[11]);
  and and_a22_b12 (and_12[22], i0[22], i1[12]);
  and and_a22_b13 (and_13[22], i0[22], i1[13]);
  and and_a22_b14 (and_14[22], i0[22], i1[14]);
  and and_a22_b15 (and_15[22], i0[22], i1[15]);
  and and_a22_b16 (and_16[22], i0[22], i1[16]);
  and and_a22_b17 (and_17[22], i0[22], i1[17]);
  and and_a22_b18 (and_18[22], i0[22], i1[18]);
  and and_a22_b19 (and_19[22], i0[22], i1[19]);
  and and_a22_b2 (and_2[22], i0[22], i1[2]);
  and and_a22_b20 (and_20[22], i0[22], i1[20]);
  and and_a22_b21 (and_21[22], i0[22], i1[21]);
  and and_a22_b22 (and_22[22], i0[22], i1[22]);
  and and_a22_b23 (and_23[22], i0[22], i1[23]);
  and and_a22_b3 (and_3[22], i0[22], i1[3]);
  and and_a22_b4 (and_4[22], i0[22], i1[4]);
  and and_a22_b5 (and_5[22], i0[22], i1[5]);
  and and_a22_b6 (and_6[22], i0[22], i1[6]);
  and and_a22_b7 (and_7[22], i0[22], i1[7]);
  and and_a22_b8 (and_8[22], i0[22], i1[8]);
  and and_a22_b9 (and_9[22], i0[22], i1[9]);
  and and_a23_b0 (and_0[23], i0[23], i1[0]);
  and and_a23_b1 (and_1[23], i0[23], i1[1]);
  and and_a23_b10 (and_10[23], i0[23], i1[10]);
  and and_a23_b11 (and_11[23], i0[23], i1[11]);
  and and_a23_b12 (and_12[23], i0[23], i1[12]);
  and and_a23_b13 (and_13[23], i0[23], i1[13]);
  and and_a23_b14 (and_14[23], i0[23], i1[14]);
  and and_a23_b15 (and_15[23], i0[23], i1[15]);
  and and_a23_b16 (and_16[23], i0[23], i1[16]);
  and and_a23_b17 (and_17[23], i0[23], i1[17]);
  and and_a23_b18 (and_18[23], i0[23], i1[18]);
  and and_a23_b19 (and_19[23], i0[23], i1[19]);
  and and_a23_b2 (and_2[23], i0[23], i1[2]);
  and and_a23_b20 (and_20[23], i0[23], i1[20]);
  and and_a23_b21 (and_21[23], i0[23], i1[21]);
  and and_a23_b22 (and_22[23], i0[23], i1[22]);
  and and_a23_b23 (and_23[23], i0[23], i1[23]);
  and and_a23_b3 (and_3[23], i0[23], i1[3]);
  and and_a23_b4 (and_4[23], i0[23], i1[4]);
  and and_a23_b5 (and_5[23], i0[23], i1[5]);
  and and_a23_b6 (and_6[23], i0[23], i1[6]);
  and and_a23_b7 (and_7[23], i0[23], i1[7]);
  and and_a23_b8 (and_8[23], i0[23], i1[8]);
  and and_a23_b9 (and_9[23], i0[23], i1[9]);
  and and_a2_b0 (and_0[2], i0[2], i1[0]);
  and and_a2_b1 (and_1[2], i0[2], i1[1]);
  and and_a2_b10 (and_10[2], i0[2], i1[10]);
  and and_a2_b11 (and_11[2], i0[2], i1[11]);
  and and_a2_b12 (and_12[2], i0[2], i1[12]);
  and and_a2_b13 (and_13[2], i0[2], i1[13]);
  and and_a2_b14 (and_14[2], i0[2], i1[14]);
  and and_a2_b15 (and_15[2], i0[2], i1[15]);
  and and_a2_b16 (and_16[2], i0[2], i1[16]);
  and and_a2_b17 (and_17[2], i0[2], i1[17]);
  and and_a2_b18 (and_18[2], i0[2], i1[18]);
  and and_a2_b19 (and_19[2], i0[2], i1[19]);
  and and_a2_b2 (and_2[2], i0[2], i1[2]);
  and and_a2_b20 (and_20[2], i0[2], i1[20]);
  and and_a2_b21 (and_21[2], i0[2], i1[21]);
  and and_a2_b22 (and_22[2], i0[2], i1[22]);
  and and_a2_b23 (and_23[2], i0[2], i1[23]);
  and and_a2_b3 (and_3[2], i0[2], i1[3]);
  and and_a2_b4 (and_4[2], i0[2], i1[4]);
  and and_a2_b5 (and_5[2], i0[2], i1[5]);
  and and_a2_b6 (and_6[2], i0[2], i1[6]);
  and and_a2_b7 (and_7[2], i0[2], i1[7]);
  and and_a2_b8 (and_8[2], i0[2], i1[8]);
  and and_a2_b9 (and_9[2], i0[2], i1[9]);
  and and_a3_b0 (and_0[3], i0[3], i1[0]);
  and and_a3_b1 (and_1[3], i0[3], i1[1]);
  and and_a3_b10 (and_10[3], i0[3], i1[10]);
  and and_a3_b11 (and_11[3], i0[3], i1[11]);
  and and_a3_b12 (and_12[3], i0[3], i1[12]);
  and and_a3_b13 (and_13[3], i0[3], i1[13]);
  and and_a3_b14 (and_14[3], i0[3], i1[14]);
  and and_a3_b15 (and_15[3], i0[3], i1[15]);
  and and_a3_b16 (and_16[3], i0[3], i1[16]);
  and and_a3_b17 (and_17[3], i0[3], i1[17]);
  and and_a3_b18 (and_18[3], i0[3], i1[18]);
  and and_a3_b19 (and_19[3], i0[3], i1[19]);
  and and_a3_b2 (and_2[3], i0[3], i1[2]);
  and and_a3_b20 (and_20[3], i0[3], i1[20]);
  and and_a3_b21 (and_21[3], i0[3], i1[21]);
  and and_a3_b22 (and_22[3], i0[3], i1[22]);
  and and_a3_b23 (and_23[3], i0[3], i1[23]);
  and and_a3_b3 (and_3[3], i0[3], i1[3]);
  and and_a3_b4 (and_4[3], i0[3], i1[4]);
  and and_a3_b5 (and_5[3], i0[3], i1[5]);
  and and_a3_b6 (and_6[3], i0[3], i1[6]);
  and and_a3_b7 (and_7[3], i0[3], i1[7]);
  and and_a3_b8 (and_8[3], i0[3], i1[8]);
  and and_a3_b9 (and_9[3], i0[3], i1[9]);
  and and_a4_b0 (and_0[4], i0[4], i1[0]);
  and and_a4_b1 (and_1[4], i0[4], i1[1]);
  and and_a4_b10 (and_10[4], i0[4], i1[10]);
  and and_a4_b11 (and_11[4], i0[4], i1[11]);
  and and_a4_b12 (and_12[4], i0[4], i1[12]);
  and and_a4_b13 (and_13[4], i0[4], i1[13]);
  and and_a4_b14 (and_14[4], i0[4], i1[14]);
  and and_a4_b15 (and_15[4], i0[4], i1[15]);
  and and_a4_b16 (and_16[4], i0[4], i1[16]);
  and and_a4_b17 (and_17[4], i0[4], i1[17]);
  and and_a4_b18 (and_18[4], i0[4], i1[18]);
  and and_a4_b19 (and_19[4], i0[4], i1[19]);
  and and_a4_b2 (and_2[4], i0[4], i1[2]);
  and and_a4_b20 (and_20[4], i0[4], i1[20]);
  and and_a4_b21 (and_21[4], i0[4], i1[21]);
  and and_a4_b22 (and_22[4], i0[4], i1[22]);
  and and_a4_b23 (and_23[4], i0[4], i1[23]);
  and and_a4_b3 (and_3[4], i0[4], i1[3]);
  and and_a4_b4 (and_4[4], i0[4], i1[4]);
  and and_a4_b5 (and_5[4], i0[4], i1[5]);
  and and_a4_b6 (and_6[4], i0[4], i1[6]);
  and and_a4_b7 (and_7[4], i0[4], i1[7]);
  and and_a4_b8 (and_8[4], i0[4], i1[8]);
  and and_a4_b9 (and_9[4], i0[4], i1[9]);
  and and_a5_b0 (and_0[5], i0[5], i1[0]);
  and and_a5_b1 (and_1[5], i0[5], i1[1]);
  and and_a5_b10 (and_10[5], i0[5], i1[10]);
  and and_a5_b11 (and_11[5], i0[5], i1[11]);
  and and_a5_b12 (and_12[5], i0[5], i1[12]);
  and and_a5_b13 (and_13[5], i0[5], i1[13]);
  and and_a5_b14 (and_14[5], i0[5], i1[14]);
  and and_a5_b15 (and_15[5], i0[5], i1[15]);
  and and_a5_b16 (and_16[5], i0[5], i1[16]);
  and and_a5_b17 (and_17[5], i0[5], i1[17]);
  and and_a5_b18 (and_18[5], i0[5], i1[18]);
  and and_a5_b19 (and_19[5], i0[5], i1[19]);
  and and_a5_b2 (and_2[5], i0[5], i1[2]);
  and and_a5_b20 (and_20[5], i0[5], i1[20]);
  and and_a5_b21 (and_21[5], i0[5], i1[21]);
  and and_a5_b22 (and_22[5], i0[5], i1[22]);
  and and_a5_b23 (and_23[5], i0[5], i1[23]);
  and and_a5_b3 (and_3[5], i0[5], i1[3]);
  and and_a5_b4 (and_4[5], i0[5], i1[4]);
  and and_a5_b5 (and_5[5], i0[5], i1[5]);
  and and_a5_b6 (and_6[5], i0[5], i1[6]);
  and and_a5_b7 (and_7[5], i0[5], i1[7]);
  and and_a5_b8 (and_8[5], i0[5], i1[8]);
  and and_a5_b9 (and_9[5], i0[5], i1[9]);
  and and_a6_b0 (and_0[6], i0[6], i1[0]);
  and and_a6_b1 (and_1[6], i0[6], i1[1]);
  and and_a6_b10 (and_10[6], i0[6], i1[10]);
  and and_a6_b11 (and_11[6], i0[6], i1[11]);
  and and_a6_b12 (and_12[6], i0[6], i1[12]);
  and and_a6_b13 (and_13[6], i0[6], i1[13]);
  and and_a6_b14 (and_14[6], i0[6], i1[14]);
  and and_a6_b15 (and_15[6], i0[6], i1[15]);
  and and_a6_b16 (and_16[6], i0[6], i1[16]);
  and and_a6_b17 (and_17[6], i0[6], i1[17]);
  and and_a6_b18 (and_18[6], i0[6], i1[18]);
  and and_a6_b19 (and_19[6], i0[6], i1[19]);
  and and_a6_b2 (and_2[6], i0[6], i1[2]);
  and and_a6_b20 (and_20[6], i0[6], i1[20]);
  and and_a6_b21 (and_21[6], i0[6], i1[21]);
  and and_a6_b22 (and_22[6], i0[6], i1[22]);
  and and_a6_b23 (and_23[6], i0[6], i1[23]);
  and and_a6_b3 (and_3[6], i0[6], i1[3]);
  and and_a6_b4 (and_4[6], i0[6], i1[4]);
  and and_a6_b5 (and_5[6], i0[6], i1[5]);
  and and_a6_b6 (and_6[6], i0[6], i1[6]);
  and and_a6_b7 (and_7[6], i0[6], i1[7]);
  and and_a6_b8 (and_8[6], i0[6], i1[8]);
  and and_a6_b9 (and_9[6], i0[6], i1[9]);
  and and_a7_b0 (and_0[7], i0[7], i1[0]);
  and and_a7_b1 (and_1[7], i0[7], i1[1]);
  and and_a7_b10 (and_10[7], i0[7], i1[10]);
  and and_a7_b11 (and_11[7], i0[7], i1[11]);
  and and_a7_b12 (and_12[7], i0[7], i1[12]);
  and and_a7_b13 (and_13[7], i0[7], i1[13]);
  and and_a7_b14 (and_14[7], i0[7], i1[14]);
  and and_a7_b15 (and_15[7], i0[7], i1[15]);
  and and_a7_b16 (and_16[7], i0[7], i1[16]);
  and and_a7_b17 (and_17[7], i0[7], i1[17]);
  and and_a7_b18 (and_18[7], i0[7], i1[18]);
  and and_a7_b19 (and_19[7], i0[7], i1[19]);
  and and_a7_b2 (and_2[7], i0[7], i1[2]);
  and and_a7_b20 (and_20[7], i0[7], i1[20]);
  and and_a7_b21 (and_21[7], i0[7], i1[21]);
  and and_a7_b22 (and_22[7], i0[7], i1[22]);
  and and_a7_b23 (and_23[7], i0[7], i1[23]);
  and and_a7_b3 (and_3[7], i0[7], i1[3]);
  and and_a7_b4 (and_4[7], i0[7], i1[4]);
  and and_a7_b5 (and_5[7], i0[7], i1[5]);
  and and_a7_b6 (and_6[7], i0[7], i1[6]);
  and and_a7_b7 (and_7[7], i0[7], i1[7]);
  and and_a7_b8 (and_8[7], i0[7], i1[8]);
  and and_a7_b9 (and_9[7], i0[7], i1[9]);
  and and_a8_b0 (and_0[8], i0[8], i1[0]);
  and and_a8_b1 (and_1[8], i0[8], i1[1]);
  and and_a8_b10 (and_10[8], i0[8], i1[10]);
  and and_a8_b11 (and_11[8], i0[8], i1[11]);
  and and_a8_b12 (and_12[8], i0[8], i1[12]);
  and and_a8_b13 (and_13[8], i0[8], i1[13]);
  and and_a8_b14 (and_14[8], i0[8], i1[14]);
  and and_a8_b15 (and_15[8], i0[8], i1[15]);
  and and_a8_b16 (and_16[8], i0[8], i1[16]);
  and and_a8_b17 (and_17[8], i0[8], i1[17]);
  and and_a8_b18 (and_18[8], i0[8], i1[18]);
  and and_a8_b19 (and_19[8], i0[8], i1[19]);
  and and_a8_b2 (and_2[8], i0[8], i1[2]);
  and and_a8_b20 (and_20[8], i0[8], i1[20]);
  and and_a8_b21 (and_21[8], i0[8], i1[21]);
  and and_a8_b22 (and_22[8], i0[8], i1[22]);
  and and_a8_b23 (and_23[8], i0[8], i1[23]);
  and and_a8_b3 (and_3[8], i0[8], i1[3]);
  and and_a8_b4 (and_4[8], i0[8], i1[4]);
  and and_a8_b5 (and_5[8], i0[8], i1[5]);
  and and_a8_b6 (and_6[8], i0[8], i1[6]);
  and and_a8_b7 (and_7[8], i0[8], i1[7]);
  and and_a8_b8 (and_8[8], i0[8], i1[8]);
  and and_a8_b9 (and_9[8], i0[8], i1[9]);
  and and_a9_b0 (and_0[9], i0[9], i1[0]);
  and and_a9_b1 (and_1[9], i0[9], i1[1]);
  and and_a9_b10 (and_10[9], i0[9], i1[10]);
  and and_a9_b11 (and_11[9], i0[9], i1[11]);
  and and_a9_b12 (and_12[9], i0[9], i1[12]);
  and and_a9_b13 (and_13[9], i0[9], i1[13]);
  and and_a9_b14 (and_14[9], i0[9], i1[14]);
  and and_a9_b15 (and_15[9], i0[9], i1[15]);
  and and_a9_b16 (and_16[9], i0[9], i1[16]);
  and and_a9_b17 (and_17[9], i0[9], i1[17]);
  and and_a9_b18 (and_18[9], i0[9], i1[18]);
  and and_a9_b19 (and_19[9], i0[9], i1[19]);
  and and_a9_b2 (and_2[9], i0[9], i1[2]);
  and and_a9_b20 (and_20[9], i0[9], i1[20]);
  and and_a9_b21 (and_21[9], i0[9], i1[21]);
  and and_a9_b22 (and_22[9], i0[9], i1[22]);
  and and_a9_b23 (and_23[9], i0[9], i1[23]);
  and and_a9_b3 (and_3[9], i0[9], i1[3]);
  and and_a9_b4 (and_4[9], i0[9], i1[4]);
  and and_a9_b5 (and_5[9], i0[9], i1[5]);
  and and_a9_b6 (and_6[9], i0[9], i1[6]);
  and and_a9_b7 (and_7[9], i0[9], i1[7]);
  and and_a9_b8 (and_8[9], i0[9], i1[8]);
  and and_a9_b9 (and_9[9], i0[9], i1[9]);
  add_pu47_pu46_pu45_pu44_pu43_pu42_pu41_pu40_pu39_pu38_pu37_pu36_pu35_pu34_pu33_pu32_pu31_pu30_pu29_pu28_pu27_pu26_pu25_pu24_o48 sum (
    .i0({and_23[23],and_22[23],and_21[23],and_20[23],and_19[23],and_18[23],and_17[23],and_16[23],and_15[23],and_14[23],and_13[23],and_12[23],and_11[23],and_10[23],and_9[23],and_8[23],and_7[23],and_6[23],and_5[23],and_4[23],and_3[23],and_2[23],and_1[23],and_0}),
    .i1({and_23[22],and_22[22],and_21[22],and_20[22],and_19[22],and_18[22],and_17[22],and_16[22],and_15[22],and_14[22],and_13[22],and_12[22],and_11[22],and_10[22],and_9[22],and_8[22],and_7[22],and_6[22],and_5[22],and_4[22],and_3[22],and_2[22],and_1[22:0],1'b0}),
    .i10({and_23[13],and_22[13],and_21[13],and_20[13],and_19[13],and_18[13],and_17[13],and_16[13],and_15[13],and_14[13],and_13[13],and_12[13],and_11[13],and_10[13:0],10'b0000000000}),
    .i11({and_23[12],and_22[12],and_21[12],and_20[12],and_19[12],and_18[12],and_17[12],and_16[12],and_15[12],and_14[12],and_13[12],and_12[12],and_11[12:0],11'b00000000000}),
    .i12({and_23[11],and_22[11],and_21[11],and_20[11],and_19[11],and_18[11],and_17[11],and_16[11],and_15[11],and_14[11],and_13[11],and_12[11:0],12'b000000000000}),
    .i13({and_23[10],and_22[10],and_21[10],and_20[10],and_19[10],and_18[10],and_17[10],and_16[10],and_15[10],and_14[10],and_13[10:0],13'b0000000000000}),
    .i14({and_23[9],and_22[9],and_21[9],and_20[9],and_19[9],and_18[9],and_17[9],and_16[9],and_15[9],and_14[9:0],14'b00000000000000}),
    .i15({and_23[8],and_22[8],and_21[8],and_20[8],and_19[8],and_18[8],and_17[8],and_16[8],and_15[8:0],15'b000000000000000}),
    .i16({and_23[7],and_22[7],and_21[7],and_20[7],and_19[7],and_18[7],and_17[7],and_16[7:0],16'b0000000000000000}),
    .i17({and_23[6],and_22[6],and_21[6],and_20[6],and_19[6],and_18[6],and_17[6:0],17'b00000000000000000}),
    .i18({and_23[5],and_22[5],and_21[5],and_20[5],and_19[5],and_18[5:0],18'b000000000000000000}),
    .i19({and_23[4],and_22[4],and_21[4],and_20[4],and_19[4:0],19'b0000000000000000000}),
    .i2({and_23[21],and_22[21],and_21[21],and_20[21],and_19[21],and_18[21],and_17[21],and_16[21],and_15[21],and_14[21],and_13[21],and_12[21],and_11[21],and_10[21],and_9[21],and_8[21],and_7[21],and_6[21],and_5[21],and_4[21],and_3[21],and_2[21:0],2'b00}),
    .i20({and_23[3],and_22[3],and_21[3],and_20[3:0],20'b00000000000000000000}),
    .i21({and_23[2],and_22[2],and_21[2:0],21'b000000000000000000000}),
    .i22({and_23[1],and_22[1:0],22'b0000000000000000000000}),
    .i23({and_23[0],23'b00000000000000000000000}),
    .i3({and_23[20],and_22[20],and_21[20],and_20[20],and_19[20],and_18[20],and_17[20],and_16[20],and_15[20],and_14[20],and_13[20],and_12[20],and_11[20],and_10[20],and_9[20],and_8[20],and_7[20],and_6[20],and_5[20],and_4[20],and_3[20:0],3'b000}),
    .i4({and_23[19],and_22[19],and_21[19],and_20[19],and_19[19],and_18[19],and_17[19],and_16[19],and_15[19],and_14[19],and_13[19],and_12[19],and_11[19],and_10[19],and_9[19],and_8[19],and_7[19],and_6[19],and_5[19],and_4[19:0],4'b0000}),
    .i5({and_23[18],and_22[18],and_21[18],and_20[18],and_19[18],and_18[18],and_17[18],and_16[18],and_15[18],and_14[18],and_13[18],and_12[18],and_11[18],and_10[18],and_9[18],and_8[18],and_7[18],and_6[18],and_5[18:0],5'b00000}),
    .i6({and_23[17],and_22[17],and_21[17],and_20[17],and_19[17],and_18[17],and_17[17],and_16[17],and_15[17],and_14[17],and_13[17],and_12[17],and_11[17],and_10[17],and_9[17],and_8[17],and_7[17],and_6[17:0],6'b000000}),
    .i7({and_23[16],and_22[16],and_21[16],and_20[16],and_19[16],and_18[16],and_17[16],and_16[16],and_15[16],and_14[16],and_13[16],and_12[16],and_11[16],and_10[16],and_9[16],and_8[16],and_7[16:0],7'b0000000}),
    .i8({and_23[15],and_22[15],and_21[15],and_20[15],and_19[15],and_18[15],and_17[15],and_16[15],and_15[15],and_14[15],and_13[15],and_12[15],and_11[15],and_10[15],and_9[15],and_8[15:0],8'b00000000}),
    .i9({and_23[14],and_22[14],and_21[14],and_20[14],and_19[14],and_18[14],and_17[14],and_16[14],and_15[14],and_14[14],and_13[14],and_12[14],and_11[14],and_10[14],and_9[14:0],9'b000000000}),
    .o(o));

endmodule 

module add_sub  // ../RTL/core/fpu.v(83)
  (
  n1,
  n2,
  sub,
  Exception,
  Overflow,
  Underflow,
  result
  );

  input [31:0] n1;  // ../RTL/core/fpu.v(84)
  input [31:0] n2;  // ../RTL/core/fpu.v(85)
  input sub;  // ../RTL/core/fpu.v(87)
  output Exception;  // ../RTL/core/fpu.v(90)
  output Overflow;  // ../RTL/core/fpu.v(88)
  output Underflow;  // ../RTL/core/fpu.v(89)
  output [31:0] result;  // ../RTL/core/fpu.v(86)

  wire [7:0] \C023/outtemp ;  // ../RTL/core/fpu_utils.v(93)
  wire [23:0] \C03/outtemp ;  // ../RTL/core/fpu_utils.v(99)
  wire [7:0] E;  // ../RTL/core/fpu.v(95)
  wire [23:0] M1;  // ../RTL/core/fpu.v(97)
  wire [23:0] M2;  // ../RTL/core/fpu.v(97)
  wire [23:0] M_result;  // ../RTL/core/fpu.v(97)
  wire [23:0] M_result2;  // ../RTL/core/fpu.v(97)
  wire [22:0] \NM/n122 ;
  wire [22:0] \NM/n4 ;
  wire  \NM/sel0_b1/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b1/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b10/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B13 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b11/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B12 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B13 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b12/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B11 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B12 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B13 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b13/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B10 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B11 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B12 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B13 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b14/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B10 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B11 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B12 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B13 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b15/B9 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B10 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B11 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B12 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B13 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B8 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b16/B9 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B10 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B11 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B12 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B13 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B7 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B8 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b17/B9 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B10 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B11 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B12 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B13 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B6 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B7 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B8 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b18/B9 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B10 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B11 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B12 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B13 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B5 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B6 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B7 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B8 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b19/B9 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b2/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b2/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b2/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B10 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B11 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B12 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B13 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B4 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B5 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B6 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B7 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B8 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b20/B9 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B10 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B11 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B12 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B13 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B3 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B4 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B5 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B6 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B7 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B8 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b21/B9 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B10 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B11 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B12 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B13 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B14 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B2 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B3 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B4 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B5 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B6 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B7 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B8 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b22/B9 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b3/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b3/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b3/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b3/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b4/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b4/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b4/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b4/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b4/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b5/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b5/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b5/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b5/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b5/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b5/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b6/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b7/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b8/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B15 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B16 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B17 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B18 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B19 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B20 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B21 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B22 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B23 ;  // ../RTL/core/fpu_utils.v(163)
  wire  \NM/sel0_b9/B24 ;  // ../RTL/core/fpu_utils.v(163)
  wire [7:0] One_Added_E;  // ../RTL/core/fpu.v(95)
  wire [7:0] complemented_E2;  // ../RTL/core/fpu.v(95)
  wire [23:0] complemented_M_result;  // ../RTL/core/fpu.v(97)
  wire [7:0] complemented_shift_E;  // ../RTL/core/fpu.v(95)
  wire [7:0] complemented_temp_exp_diff;  // ../RTL/core/fpu.v(95)
  wire [7:0] exp_diff;  // ../RTL/core/fpu.v(95)
  wire [23:0] n37;
  wire [23:0] n62;
  wire [7:0] new_E;  // ../RTL/core/fpu.v(95)
  wire [23:0] new_M2;  // ../RTL/core/fpu.v(97)
  wire [4:0] shift_E;  // ../RTL/core/fpu.v(100)
  wire [7:0] temp_exp_diff;  // ../RTL/core/fpu.v(95)
  wire \ADD01/ADD01/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/n1 ;
  wire \ADD01/ADD01/n10 ;
  wire \ADD01/ADD01/n12 ;
  wire \ADD01/ADD01/n13 ;
  wire \ADD01/ADD01/n14 ;
  wire \ADD01/ADD01/n15 ;
  wire \ADD01/ADD01/n16 ;
  wire \ADD01/ADD01/n17 ;
  wire \ADD01/ADD01/n18 ;
  wire \ADD01/ADD01/n19 ;
  wire \ADD01/ADD01/n2 ;
  wire \ADD01/ADD01/n20 ;
  wire \ADD01/ADD01/n3 ;
  wire \ADD01/ADD01/n5 ;
  wire \ADD01/ADD01/n6 ;
  wire \ADD01/ADD01/n7 ;
  wire \ADD01/ADD01/n8 ;
  wire \ADD01/ADD01/n9 ;
  wire \ADD01/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/p0_neg ;
  wire \ADD01/ADD01/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/n0 ;
  wire \ADD01/ADD02/n1 ;
  wire \ADD01/ADD02/n10 ;
  wire \ADD01/ADD02/n11 ;
  wire \ADD01/ADD02/n12 ;
  wire \ADD01/ADD02/n13 ;
  wire \ADD01/ADD02/n14 ;
  wire \ADD01/ADD02/n15 ;
  wire \ADD01/ADD02/n16 ;
  wire \ADD01/ADD02/n17 ;
  wire \ADD01/ADD02/n18 ;
  wire \ADD01/ADD02/n19 ;
  wire \ADD01/ADD02/n2 ;
  wire \ADD01/ADD02/n20 ;
  wire \ADD01/ADD02/n21 ;
  wire \ADD01/ADD02/n3 ;
  wire \ADD01/ADD02/n4 ;
  wire \ADD01/ADD02/n5 ;
  wire \ADD01/ADD02/n6 ;
  wire \ADD01/ADD02/n7 ;
  wire \ADD01/ADD02/n8 ;
  wire \ADD01/ADD02/n9 ;
  wire \ADD01/ADD02/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ctemp ;  // ../RTL/core/fpu_utils.v(76)
  wire \ADD02/ADD01/ADD01/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/n0 ;
  wire \ADD02/ADD01/ADD01/n1 ;
  wire \ADD02/ADD01/ADD01/n10 ;
  wire \ADD02/ADD01/ADD01/n11 ;
  wire \ADD02/ADD01/ADD01/n12 ;
  wire \ADD02/ADD01/ADD01/n13 ;
  wire \ADD02/ADD01/ADD01/n14 ;
  wire \ADD02/ADD01/ADD01/n15 ;
  wire \ADD02/ADD01/ADD01/n16 ;
  wire \ADD02/ADD01/ADD01/n17 ;
  wire \ADD02/ADD01/ADD01/n18 ;
  wire \ADD02/ADD01/ADD01/n19 ;
  wire \ADD02/ADD01/ADD01/n2 ;
  wire \ADD02/ADD01/ADD01/n20 ;
  wire \ADD02/ADD01/ADD01/n21 ;
  wire \ADD02/ADD01/ADD01/n3 ;
  wire \ADD02/ADD01/ADD01/n4 ;
  wire \ADD02/ADD01/ADD01/n5 ;
  wire \ADD02/ADD01/ADD01/n6 ;
  wire \ADD02/ADD01/ADD01/n7 ;
  wire \ADD02/ADD01/ADD01/n8 ;
  wire \ADD02/ADD01/ADD01/n9 ;
  wire \ADD02/ADD01/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/n0 ;
  wire \ADD02/ADD01/ADD02/n1 ;
  wire \ADD02/ADD01/ADD02/n10 ;
  wire \ADD02/ADD01/ADD02/n11 ;
  wire \ADD02/ADD01/ADD02/n12 ;
  wire \ADD02/ADD01/ADD02/n13 ;
  wire \ADD02/ADD01/ADD02/n14 ;
  wire \ADD02/ADD01/ADD02/n15 ;
  wire \ADD02/ADD01/ADD02/n16 ;
  wire \ADD02/ADD01/ADD02/n17 ;
  wire \ADD02/ADD01/ADD02/n18 ;
  wire \ADD02/ADD01/ADD02/n19 ;
  wire \ADD02/ADD01/ADD02/n2 ;
  wire \ADD02/ADD01/ADD02/n20 ;
  wire \ADD02/ADD01/ADD02/n21 ;
  wire \ADD02/ADD01/ADD02/n3 ;
  wire \ADD02/ADD01/ADD02/n4 ;
  wire \ADD02/ADD01/ADD02/n5 ;
  wire \ADD02/ADD01/ADD02/n6 ;
  wire \ADD02/ADD01/ADD02/n7 ;
  wire \ADD02/ADD01/ADD02/n8 ;
  wire \ADD02/ADD01/ADD02/n9 ;
  wire \ADD02/ADD01/ADD02/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ctemp ;  // ../RTL/core/fpu_utils.v(76)
  wire \ADD02/ADD02/ADD01/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/n0 ;
  wire \ADD02/ADD02/ADD01/n1 ;
  wire \ADD02/ADD02/ADD01/n10 ;
  wire \ADD02/ADD02/ADD01/n11 ;
  wire \ADD02/ADD02/ADD01/n12 ;
  wire \ADD02/ADD02/ADD01/n13 ;
  wire \ADD02/ADD02/ADD01/n14 ;
  wire \ADD02/ADD02/ADD01/n15 ;
  wire \ADD02/ADD02/ADD01/n16 ;
  wire \ADD02/ADD02/ADD01/n17 ;
  wire \ADD02/ADD02/ADD01/n18 ;
  wire \ADD02/ADD02/ADD01/n19 ;
  wire \ADD02/ADD02/ADD01/n2 ;
  wire \ADD02/ADD02/ADD01/n20 ;
  wire \ADD02/ADD02/ADD01/n21 ;
  wire \ADD02/ADD02/ADD01/n3 ;
  wire \ADD02/ADD02/ADD01/n4 ;
  wire \ADD02/ADD02/ADD01/n5 ;
  wire \ADD02/ADD02/ADD01/n6 ;
  wire \ADD02/ADD02/ADD01/n7 ;
  wire \ADD02/ADD02/ADD01/n8 ;
  wire \ADD02/ADD02/ADD01/n9 ;
  wire \ADD02/ADD02/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/n0 ;
  wire \ADD02/ADD02/ADD02/n1 ;
  wire \ADD02/ADD02/ADD02/n10 ;
  wire \ADD02/ADD02/ADD02/n11 ;
  wire \ADD02/ADD02/ADD02/n12 ;
  wire \ADD02/ADD02/ADD02/n13 ;
  wire \ADD02/ADD02/ADD02/n14 ;
  wire \ADD02/ADD02/ADD02/n15 ;
  wire \ADD02/ADD02/ADD02/n16 ;
  wire \ADD02/ADD02/ADD02/n17 ;
  wire \ADD02/ADD02/ADD02/n18 ;
  wire \ADD02/ADD02/ADD02/n19 ;
  wire \ADD02/ADD02/ADD02/n2 ;
  wire \ADD02/ADD02/ADD02/n20 ;
  wire \ADD02/ADD02/ADD02/n21 ;
  wire \ADD02/ADD02/ADD02/n3 ;
  wire \ADD02/ADD02/ADD02/n4 ;
  wire \ADD02/ADD02/ADD02/n5 ;
  wire \ADD02/ADD02/ADD02/n6 ;
  wire \ADD02/ADD02/ADD02/n7 ;
  wire \ADD02/ADD02/ADD02/n8 ;
  wire \ADD02/ADD02/ADD02/n9 ;
  wire \ADD02/ADD02/ADD02/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ctemp ;  // ../RTL/core/fpu_utils.v(76)
  wire \ADD02/ADD03/ADD01/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/n0 ;
  wire \ADD02/ADD03/ADD01/n1 ;
  wire \ADD02/ADD03/ADD01/n10 ;
  wire \ADD02/ADD03/ADD01/n11 ;
  wire \ADD02/ADD03/ADD01/n12 ;
  wire \ADD02/ADD03/ADD01/n13 ;
  wire \ADD02/ADD03/ADD01/n14 ;
  wire \ADD02/ADD03/ADD01/n15 ;
  wire \ADD02/ADD03/ADD01/n16 ;
  wire \ADD02/ADD03/ADD01/n17 ;
  wire \ADD02/ADD03/ADD01/n18 ;
  wire \ADD02/ADD03/ADD01/n19 ;
  wire \ADD02/ADD03/ADD01/n2 ;
  wire \ADD02/ADD03/ADD01/n20 ;
  wire \ADD02/ADD03/ADD01/n21 ;
  wire \ADD02/ADD03/ADD01/n3 ;
  wire \ADD02/ADD03/ADD01/n4 ;
  wire \ADD02/ADD03/ADD01/n5 ;
  wire \ADD02/ADD03/ADD01/n6 ;
  wire \ADD02/ADD03/ADD01/n7 ;
  wire \ADD02/ADD03/ADD01/n8 ;
  wire \ADD02/ADD03/ADD01/n9 ;
  wire \ADD02/ADD03/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/n0 ;
  wire \ADD02/ADD03/ADD02/n1 ;
  wire \ADD02/ADD03/ADD02/n10 ;
  wire \ADD02/ADD03/ADD02/n11 ;
  wire \ADD02/ADD03/ADD02/n12 ;
  wire \ADD02/ADD03/ADD02/n13 ;
  wire \ADD02/ADD03/ADD02/n14 ;
  wire \ADD02/ADD03/ADD02/n15 ;
  wire \ADD02/ADD03/ADD02/n16 ;
  wire \ADD02/ADD03/ADD02/n17 ;
  wire \ADD02/ADD03/ADD02/n18 ;
  wire \ADD02/ADD03/ADD02/n19 ;
  wire \ADD02/ADD03/ADD02/n2 ;
  wire \ADD02/ADD03/ADD02/n20 ;
  wire \ADD02/ADD03/ADD02/n21 ;
  wire \ADD02/ADD03/ADD02/n3 ;
  wire \ADD02/ADD03/ADD02/n4 ;
  wire \ADD02/ADD03/ADD02/n5 ;
  wire \ADD02/ADD03/ADD02/n6 ;
  wire \ADD02/ADD03/ADD02/n7 ;
  wire \ADD02/ADD03/ADD02/n8 ;
  wire \ADD02/ADD03/ADD02/n9 ;
  wire \ADD02/ADD03/ADD02/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ctemp ;  // ../RTL/core/fpu_utils.v(76)
  wire \ADD02/ctemp1 ;  // ../RTL/core/fpu_utils.v(87)
  wire \ADD02/ctemp2 ;  // ../RTL/core/fpu_utils.v(88)
  wire \ADD0212/ADD01/n1 ;
  wire \ADD0212/ADD01/n14 ;
  wire \ADD0212/ADD01/n17 ;
  wire \ADD0212/ADD01/n18 ;
  wire \ADD0212/ADD01/n7 ;
  wire \ADD0212/ADD01/n8 ;
  wire \ADD0212/ADD02/n0 ;
  wire \ADD0212/ADD02/n10 ;
  wire \ADD0212/ADD02/n11 ;
  wire \ADD0212/ADD02/n3 ;
  wire \ADD0212/ADD02/n4 ;
  wire \ADD0212/ADD02/n7 ;
  wire \ADD03/ADD01/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/n1 ;
  wire \ADD03/ADD01/n10 ;
  wire \ADD03/ADD01/n12 ;
  wire \ADD03/ADD01/n13 ;
  wire \ADD03/ADD01/n14 ;
  wire \ADD03/ADD01/n15 ;
  wire \ADD03/ADD01/n16 ;
  wire \ADD03/ADD01/n17 ;
  wire \ADD03/ADD01/n18 ;
  wire \ADD03/ADD01/n19 ;
  wire \ADD03/ADD01/n2 ;
  wire \ADD03/ADD01/n20 ;
  wire \ADD03/ADD01/n3 ;
  wire \ADD03/ADD01/n5 ;
  wire \ADD03/ADD01/n6 ;
  wire \ADD03/ADD01/n7 ;
  wire \ADD03/ADD01/n8 ;
  wire \ADD03/ADD01/n9 ;
  wire \ADD03/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/p0_neg ;
  wire \ADD03/ADD01/p1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/p2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/p3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD02/c0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD02/c1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD02/c2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD02/n0 ;
  wire \ADD03/ADD02/n1 ;
  wire \ADD03/ADD02/n10 ;
  wire \ADD03/ADD02/n11 ;
  wire \ADD03/ADD02/n2 ;
  wire \ADD03/ADD02/n3 ;
  wire \ADD03/ADD02/n4 ;
  wire \ADD03/ADD02/n5 ;
  wire \ADD03/ADD02/n6 ;
  wire \ADD03/ADD02/n7 ;
  wire \ADD03/ADD02/n8 ;
  wire \ADD03/ADD02/n9 ;
  wire \ADD03/ADD02/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ctemp ;  // ../RTL/core/fpu_utils.v(76)
  wire \C023/ADD01/ADD01/n1 ;
  wire \C023/ADD01/ADD01/n14 ;
  wire \C023/ADD01/ADD01/n17 ;
  wire \C023/ADD01/ADD01/n18 ;
  wire \C023/ADD01/ADD01/n7 ;
  wire \C023/ADD01/ADD01/n8 ;
  wire \C023/ADD01/ADD02/n0 ;
  wire \C023/ADD01/ADD02/n10 ;
  wire \C023/ADD01/ADD02/n11 ;
  wire \C023/ADD01/ADD02/n3 ;
  wire \C023/ADD01/ADD02/n4 ;
  wire \C023/ADD01/ADD02/n7 ;
  wire \C03/ADD01/ADD01/ADD01/n1 ;
  wire \C03/ADD01/ADD01/ADD01/n14 ;
  wire \C03/ADD01/ADD01/ADD01/n17 ;
  wire \C03/ADD01/ADD01/ADD01/n18 ;
  wire \C03/ADD01/ADD01/ADD01/n7 ;
  wire \C03/ADD01/ADD01/ADD01/n8 ;
  wire \C03/ADD01/ADD01/ADD02/n0 ;
  wire \C03/ADD01/ADD01/ADD02/n10 ;
  wire \C03/ADD01/ADD01/ADD02/n11 ;
  wire \C03/ADD01/ADD01/ADD02/n14 ;
  wire \C03/ADD01/ADD01/ADD02/n17 ;
  wire \C03/ADD01/ADD01/ADD02/n20 ;
  wire \C03/ADD01/ADD01/ADD02/n21 ;
  wire \C03/ADD01/ADD01/ADD02/n3 ;
  wire \C03/ADD01/ADD01/ADD02/n4 ;
  wire \C03/ADD01/ADD01/ADD02/n7 ;
  wire \C03/ADD01/ADD02/ADD01/n0 ;
  wire \C03/ADD01/ADD02/ADD01/n10 ;
  wire \C03/ADD01/ADD02/ADD01/n11 ;
  wire \C03/ADD01/ADD02/ADD01/n14 ;
  wire \C03/ADD01/ADD02/ADD01/n17 ;
  wire \C03/ADD01/ADD02/ADD01/n20 ;
  wire \C03/ADD01/ADD02/ADD01/n21 ;
  wire \C03/ADD01/ADD02/ADD01/n3 ;
  wire \C03/ADD01/ADD02/ADD01/n4 ;
  wire \C03/ADD01/ADD02/ADD01/n7 ;
  wire \C03/ADD01/ADD02/ADD02/n0 ;
  wire \C03/ADD01/ADD02/ADD02/n10 ;
  wire \C03/ADD01/ADD02/ADD02/n11 ;
  wire \C03/ADD01/ADD02/ADD02/n14 ;
  wire \C03/ADD01/ADD02/ADD02/n17 ;
  wire \C03/ADD01/ADD02/ADD02/n20 ;
  wire \C03/ADD01/ADD02/ADD02/n21 ;
  wire \C03/ADD01/ADD02/ADD02/n3 ;
  wire \C03/ADD01/ADD02/ADD02/n4 ;
  wire \C03/ADD01/ADD02/ADD02/n7 ;
  wire \C03/ADD01/ADD03/ADD01/n0 ;
  wire \C03/ADD01/ADD03/ADD01/n10 ;
  wire \C03/ADD01/ADD03/ADD01/n11 ;
  wire \C03/ADD01/ADD03/ADD01/n14 ;
  wire \C03/ADD01/ADD03/ADD01/n17 ;
  wire \C03/ADD01/ADD03/ADD01/n20 ;
  wire \C03/ADD01/ADD03/ADD01/n21 ;
  wire \C03/ADD01/ADD03/ADD01/n3 ;
  wire \C03/ADD01/ADD03/ADD01/n4 ;
  wire \C03/ADD01/ADD03/ADD01/n7 ;
  wire \C03/ADD01/ADD03/ADD02/n0 ;
  wire \C03/ADD01/ADD03/ADD02/n10 ;
  wire \C03/ADD01/ADD03/ADD02/n11 ;
  wire \C03/ADD01/ADD03/ADD02/n3 ;
  wire \C03/ADD01/ADD03/ADD02/n4 ;
  wire \C03/ADD01/ADD03/ADD02/n7 ;
  wire \M031/M01/invSL ;  // ../RTL/core/fpu_utils.v(105)
  wire \M04/M01/M01/invSL ;  // ../RTL/core/fpu_utils.v(105)
  wire M_carry;  // ../RTL/core/fpu.v(93)
  wire \NM/mux1_b0_sel_is_2_o ;
  wire \NM/mux1_b1_sel_is_2_o ;
  wire \NM/mux1_b2_sel_is_2_o ;
  wire \NM/mux1_b3_sel_is_2_o ;
  wire \NM/mux1_b4_sel_is_2_o ;
  wire \NM/n10 ;
  wire \NM/n100 ;
  wire \NM/n101 ;
  wire \NM/n102 ;
  wire \NM/n103 ;
  wire \NM/n104 ;
  wire \NM/n105 ;
  wire \NM/n106 ;
  wire \NM/n107 ;
  wire \NM/n108 ;
  wire \NM/n109 ;
  wire \NM/n11 ;
  wire \NM/n110 ;
  wire \NM/n111 ;
  wire \NM/n112 ;
  wire \NM/n113 ;
  wire \NM/n114 ;
  wire \NM/n115 ;
  wire \NM/n116 ;
  wire \NM/n117 ;
  wire \NM/n118 ;
  wire \NM/n119 ;
  wire \NM/n12 ;
  wire \NM/n124 ;
  wire \NM/n125 ;
  wire \NM/n126 ;
  wire \NM/n127 ;
  wire \NM/n128 ;
  wire \NM/n129 ;
  wire \NM/n13 ;
  wire \NM/n130 ;
  wire \NM/n132 ;
  wire \NM/n133 ;
  wire \NM/n134 ;
  wire \NM/n14 ;
  wire \NM/n142 ;
  wire \NM/n143 ;
  wire \NM/n146 ;
  wire \NM/n15 ;
  wire \NM/n153 ;
  wire \NM/n156 ;
  wire \NM/n158 ;
  wire \NM/n16 ;
  wire \NM/n165 ;
  wire \NM/n166 ;
  wire \NM/n168 ;
  wire \NM/n17 ;
  wire \NM/n170 ;
  wire \NM/n171 ;
  wire \NM/n175 ;
  wire \NM/n176 ;
  wire \NM/n177 ;
  wire \NM/n179 ;
  wire \NM/n18 ;
  wire \NM/n180 ;
  wire \NM/n182 ;
  wire \NM/n183 ;
  wire \NM/n184 ;
  wire \NM/n185 ;
  wire \NM/n186 ;
  wire \NM/n187 ;
  wire \NM/n188 ;
  wire \NM/n189 ;
  wire \NM/n19 ;
  wire \NM/n190 ;
  wire \NM/n191 ;
  wire \NM/n193 ;
  wire \NM/n194 ;
  wire \NM/n195 ;
  wire \NM/n2 ;
  wire \NM/n20 ;
  wire \NM/n202 ;
  wire \NM/n207 ;
  wire \NM/n209 ;
  wire \NM/n21 ;
  wire \NM/n210 ;
  wire \NM/n211 ;
  wire \NM/n213 ;
  wire \NM/n214 ;
  wire \NM/n215 ;
  wire \NM/n216 ;
  wire \NM/n22 ;
  wire \NM/n222 ;
  wire \NM/n227 ;
  wire \NM/n23 ;
  wire \NM/n230 ;
  wire \NM/n232 ;
  wire \NM/n234 ;
  wire \NM/n236 ;
  wire \NM/n24 ;
  wire \NM/n240 ;
  wire \NM/n242 ;
  wire \NM/n243 ;
  wire \NM/n244 ;
  wire \NM/n246 ;
  wire \NM/n247 ;
  wire \NM/n248 ;
  wire \NM/n249 ;
  wire \NM/n25 ;
  wire \NM/n251 ;
  wire \NM/n253 ;
  wire \NM/n257 ;
  wire \NM/n258 ;
  wire \NM/n26 ;
  wire \NM/n260 ;
  wire \NM/n261 ;
  wire \NM/n262 ;
  wire \NM/n263 ;
  wire \NM/n265 ;
  wire \NM/n268 ;
  wire \NM/n269 ;
  wire \NM/n27 ;
  wire \NM/n271 ;
  wire \NM/n273 ;
  wire \NM/n274 ;
  wire \NM/n276 ;
  wire \NM/n278 ;
  wire \NM/n279 ;
  wire \NM/n28 ;
  wire \NM/n280 ;
  wire \NM/n281 ;
  wire \NM/n283 ;
  wire \NM/n284 ;
  wire \NM/n286 ;
  wire \NM/n29 ;
  wire \NM/n296 ;
  wire \NM/n30 ;
  wire \NM/n300 ;
  wire \NM/n304 ;
  wire \NM/n306 ;
  wire \NM/n308 ;
  wire \NM/n31 ;
  wire \NM/n310 ;
  wire \NM/n311 ;
  wire \NM/n312 ;
  wire \NM/n313 ;
  wire \NM/n314 ;
  wire \NM/n315 ;
  wire \NM/n316 ;
  wire \NM/n318 ;
  wire \NM/n319 ;
  wire \NM/n32 ;
  wire \NM/n320 ;
  wire \NM/n321 ;
  wire \NM/n322 ;
  wire \NM/n325 ;
  wire \NM/n33 ;
  wire \NM/n331 ;
  wire \NM/n332 ;
  wire \NM/n335 ;
  wire \NM/n34 ;
  wire \NM/n340 ;
  wire \NM/n341 ;
  wire \NM/n343 ;
  wire \NM/n348 ;
  wire \NM/n349 ;
  wire \NM/n35 ;
  wire \NM/n351 ;
  wire \NM/n355 ;
  wire \NM/n357 ;
  wire \NM/n36 ;
  wire \NM/n361 ;
  wire \NM/n363 ;
  wire \NM/n366 ;
  wire \NM/n367 ;
  wire \NM/n37 ;
  wire \NM/n370 ;
  wire \NM/n371 ;
  wire \NM/n373 ;
  wire \NM/n374 ;
  wire \NM/n375 ;
  wire \NM/n376 ;
  wire \NM/n38 ;
  wire \NM/n39 ;
  wire \NM/n40 ;
  wire \NM/n41 ;
  wire \NM/n42 ;
  wire \NM/n44 ;
  wire \NM/n45 ;
  wire \NM/n46 ;
  wire \NM/n47 ;
  wire \NM/n48 ;
  wire \NM/n49 ;
  wire \NM/n50 ;
  wire \NM/n51 ;
  wire \NM/n52 ;
  wire \NM/n53 ;
  wire \NM/n54 ;
  wire \NM/n55 ;
  wire \NM/n56 ;
  wire \NM/n57 ;
  wire \NM/n58 ;
  wire \NM/n59 ;
  wire \NM/n6 ;
  wire \NM/n60 ;
  wire \NM/n61 ;
  wire \NM/n62 ;
  wire \NM/n63 ;
  wire \NM/n64 ;
  wire \NM/n65 ;
  wire \NM/n66 ;
  wire \NM/n67 ;
  wire \NM/n68 ;
  wire \NM/n69 ;
  wire \NM/n7 ;
  wire \NM/n70 ;
  wire \NM/n71 ;
  wire \NM/n72 ;
  wire \NM/n73 ;
  wire \NM/n74 ;
  wire \NM/n75 ;
  wire \NM/n76 ;
  wire \NM/n77 ;
  wire \NM/n78 ;
  wire \NM/n79 ;
  wire \NM/n8 ;
  wire \NM/n80 ;
  wire \NM/n81 ;
  wire \NM/n82 ;
  wire \NM/n83 ;
  wire \NM/n84 ;
  wire \NM/n85 ;
  wire \NM/n86 ;
  wire \NM/n87 ;
  wire \NM/n88 ;
  wire \NM/n89 ;
  wire \NM/n9 ;
  wire \NM/n90 ;
  wire \NM/n91 ;
  wire \NM/n92 ;
  wire \NM/n93 ;
  wire \NM/n94 ;
  wire \NM/n95 ;
  wire \NM/n96 ;
  wire \NM/n97 ;
  wire \NM/n98 ;
  wire \NM/n99 ;
  wire \NM/sel0_b1/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b10/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b11/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B12_or_B13_B14_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b12/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B12_or_B13_B14_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b13/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B10_B11_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B12_or_B13_B14_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b14/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B10_B11_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B12_or_B13_B14_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_B9_or_B10_B11_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b15/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B10_B11_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B12_or_B13_B14_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_B9_or_B10_B11_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_or_B6_or_B7_B8_o__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b16/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B10_B11_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B12_or_B13_B14_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B7_B8_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_B9_or_B10_B11_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_or_B6_or_B7_B8_o__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b17/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B10_B11_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B12_or_B13_B14_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B6_or_B7_B8_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B7_B8_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_B9_or_B10_B11_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_or_B6_or_B7_B8_o__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b18/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B10_B11_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B12_or_B13_B14_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B6_or_B7_B8_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B7_B8_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_B9_or_B10_B11_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_or_B6_or_B7_B8_o__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_or_or_B0_or_B1_B2_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b19/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b2/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b2/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B10_B11_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B12_or_B13_B14_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B4_B5_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B6_or_B7_B8_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B7_B8_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_B9_or_B10_B11_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_or_B6_or_B7_B8_o__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_or_or_B0_or_B1_B2_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b20/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B10_B11_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B12_or_B13_B14_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B3_or_B4_B5_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B4_B5_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B6_or_B7_B8_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B7_B8_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_B9_or_B10_B11_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_or_B6_or_B7_B8_o__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_or_or_B0_or_B1_B2_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b21/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B10_B11_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B12_or_B13_B14_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B3_or_B4_B5_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B4_B5_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B6_or_B7_B8_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B7_B8_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_B9_or_B10_B11_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_B0_or_B1_B2_o__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_B12_or_B13_B14_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_B6_or_B7_B8_o__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_or_B0_or_B1_B2_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b22/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b3/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b3/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b3/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b4/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b4/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b4/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b4/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b5/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b5/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b5/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b5/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b5/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b6/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b6/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b6/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b6/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b6/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b6/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b7/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b8/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_B15_or_B16_B17_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_B16_B17_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_B18_or_B19_B20_o_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_B21_B22_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_B23_B24_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_or_B18_or_B19_B20_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_or_B21_B22_o_or_B_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel0_b9/or_or_or_B12_or_B13__o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel1_b0_sel_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel1_b1_sel_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel1_b2_sel_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel1_b3_sel_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \NM/sel1_b4_sel_o ;  // ../RTL/core/fpu_utils.v(163)
  wire \RO01/w1 ;  // ../RTL/core/fpu_utils.v(13)
  wire \RO01/w2 ;  // ../RTL/core/fpu_utils.v(13)
  wire \RO01/w3 ;  // ../RTL/core/fpu_utils.v(13)
  wire \RO01/w4 ;  // ../RTL/core/fpu_utils.v(13)
  wire \RO01/w5 ;  // ../RTL/core/fpu_utils.v(13)
  wire \RO01/w6 ;  // ../RTL/core/fpu_utils.v(13)
  wire \exp_diff[4]_neg ;
  wire isE1GreaterThanE2;  // ../RTL/core/fpu.v(116)
  wire n10;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n11;
  wire n110;
  wire n110_neg;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n160;
  wire n161;
  wire n164;
  wire n165;
  wire n171;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire \n1[31]_neg ;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n243;
  wire n244;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n265;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n5;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n6;
  wire n60;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n7;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n8;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n9;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire \new_E[5]_neg ;
  wire \new_E[6]_neg ;
  wire \new_E[7]_neg ;
  wire real_oper;  // ../RTL/core/fpu.v(93)
  wire reduced_or_E1;  // ../RTL/core/fpu.v(94)
  wire u194_sel_is_0_o;
  wire w1;  // ../RTL/core/fpu.v(98)
  wire w2;  // ../RTL/core/fpu.v(98)
  wire w3;  // ../RTL/core/fpu.v(98)

  assign result[23] = \ADD03/ADD01/p0_neg ;
  not \ADD01/ADD01/p0_inv  (\ADD01/ADD01/p0_neg , \ADD01/ADD01/p0 );
  and \ADD01/ADD01/u0  (\ADD01/ADD01/g0 , n1[23], complemented_E2[0]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD01/ADD01/u1  (\ADD01/ADD01/g1 , n1[24], complemented_E2[1]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD01/ADD01/u10  (\ADD01/ADD01/n1 , \ADD01/ADD01/p1 , \ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD01/ADD01/u11  (\ADD01/ADD01/n2 , \ADD01/ADD01/g1 , \ADD01/ADD01/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD01/ADD01/u12  (\ADD01/ADD01/n3 , \ADD01/ADD01/p1 , \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD01/ADD01/u14  (\ADD01/ADD01/c1 , \ADD01/ADD01/n2 , \ADD01/ADD01/n3 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD01/ADD01/u15  (\ADD01/ADD01/n5 , \ADD01/ADD01/p2 , \ADD01/ADD01/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD01/ADD01/u16  (\ADD01/ADD01/n6 , \ADD01/ADD01/g2 , \ADD01/ADD01/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD01/u17  (\ADD01/ADD01/n7 , \ADD01/ADD01/p2 , \ADD01/ADD01/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD01/u18  (\ADD01/ADD01/n8 , \ADD01/ADD01/n7 , \ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD01/ADD01/u19  (\ADD01/ADD01/n9 , \ADD01/ADD01/n6 , \ADD01/ADD01/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD01/u2  (\ADD01/ADD01/g2 , n1[25], complemented_E2[2]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD01/ADD01/u20  (temp_exp_diff[3], \ADD01/ADD01/p3 , \ADD01/ADD01/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD01/ADD01/u21  (\ADD01/ADD01/n10 , \ADD01/ADD01/n7 , \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD01/ADD01/u23  (\ADD01/ADD01/c2 , \ADD01/ADD01/n9 , \ADD01/ADD01/n10 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD01/u24  (\ADD01/ADD01/n12 , \ADD01/ADD01/p3 , \ADD01/ADD01/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD01/u25  (\ADD01/ADD01/n13 , \ADD01/ADD01/g3 , \ADD01/ADD01/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD01/u26  (\ADD01/ADD01/n14 , \ADD01/ADD01/p3 , \ADD01/ADD01/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD01/u27  (\ADD01/ADD01/n15 , \ADD01/ADD01/n14 , \ADD01/ADD01/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD01/u28  (\ADD01/ADD01/n16 , \ADD01/ADD01/n13 , \ADD01/ADD01/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD01/ADD01/u29  (temp_exp_diff[2], \ADD01/ADD01/p2 , \ADD01/ADD01/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD01/ADD01/u3  (\ADD01/ADD01/g3 , n1[26], complemented_E2[3]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD01/ADD01/u30  (\ADD01/ADD01/n17 , \ADD01/ADD01/n14 , \ADD01/ADD01/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD01/u31  (\ADD01/ADD01/n18 , \ADD01/ADD01/n17 , \ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD01/u32  (\ADD01/ADD01/n19 , \ADD01/ADD01/n16 , \ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD01/ADD01/u33  (temp_exp_diff[1], \ADD01/ADD01/p1 , \ADD01/ADD01/c0 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD01/ADD01/u35  (\ADD01/ADD01/n20 , \ADD01/ADD01/n17 , \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD01/u37  (\ADD01/ctemp , \ADD01/ADD01/n19 , \ADD01/ADD01/n20 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD01/ADD01/u4  (\ADD01/ADD01/p0 , n1[23], complemented_E2[0]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD01/ADD01/u5  (\ADD01/ADD01/p1 , n1[24], complemented_E2[1]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD01/ADD01/u6  (\ADD01/ADD01/p2 , n1[25], complemented_E2[2]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD01/ADD01/u7  (\ADD01/ADD01/p3 , n1[26], complemented_E2[3]);  // ../RTL/core/fpu_utils.v(62)
  or \ADD01/ADD01/u9  (\ADD01/ADD01/c0 , \ADD01/ADD01/g0 , \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD01/ADD02/u0  (\ADD01/ADD02/g0 , n1[27], complemented_E2[4]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD01/ADD02/u1  (\ADD01/ADD02/g1 , n1[28], complemented_E2[5]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD01/ADD02/u10  (\ADD01/ADD02/n1 , \ADD01/ADD02/p1 , \ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD01/ADD02/u11  (\ADD01/ADD02/n2 , \ADD01/ADD02/g1 , \ADD01/ADD02/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD01/ADD02/u12  (\ADD01/ADD02/n3 , \ADD01/ADD02/p1 , \ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD01/ADD02/u13  (\ADD01/ADD02/n4 , \ADD01/ADD02/n3 , \ADD01/ctemp );  // ../RTL/core/fpu_utils.v(64)
  or \ADD01/ADD02/u14  (\ADD01/ADD02/c1 , \ADD01/ADD02/n2 , \ADD01/ADD02/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD01/ADD02/u15  (\ADD01/ADD02/n5 , \ADD01/ADD02/p2 , \ADD01/ADD02/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD01/ADD02/u16  (\ADD01/ADD02/n6 , \ADD01/ADD02/g2 , \ADD01/ADD02/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD02/u17  (\ADD01/ADD02/n7 , \ADD01/ADD02/p2 , \ADD01/ADD02/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD02/u18  (\ADD01/ADD02/n8 , \ADD01/ADD02/n7 , \ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD01/ADD02/u19  (\ADD01/ADD02/n9 , \ADD01/ADD02/n6 , \ADD01/ADD02/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD02/u2  (\ADD01/ADD02/g2 , n1[29], complemented_E2[6]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD01/ADD02/u20  (temp_exp_diff[7], \ADD01/ADD02/p3 , \ADD01/ADD02/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD01/ADD02/u21  (\ADD01/ADD02/n10 , \ADD01/ADD02/n7 , \ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD02/u22  (\ADD01/ADD02/n11 , \ADD01/ADD02/n10 , \ADD01/ctemp );  // ../RTL/core/fpu_utils.v(65)
  or \ADD01/ADD02/u23  (\ADD01/ADD02/c2 , \ADD01/ADD02/n9 , \ADD01/ADD02/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD01/ADD02/u24  (\ADD01/ADD02/n12 , \ADD01/ADD02/p3 , \ADD01/ADD02/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD02/u25  (\ADD01/ADD02/n13 , \ADD01/ADD02/g3 , \ADD01/ADD02/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD02/u26  (\ADD01/ADD02/n14 , \ADD01/ADD02/p3 , \ADD01/ADD02/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD02/u27  (\ADD01/ADD02/n15 , \ADD01/ADD02/n14 , \ADD01/ADD02/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD02/u28  (\ADD01/ADD02/n16 , \ADD01/ADD02/n13 , \ADD01/ADD02/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD01/ADD02/u29  (temp_exp_diff[6], \ADD01/ADD02/p2 , \ADD01/ADD02/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD01/ADD02/u3  (\ADD01/ADD02/g3 , n1[30], complemented_E2[7]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD01/ADD02/u30  (\ADD01/ADD02/n17 , \ADD01/ADD02/n14 , \ADD01/ADD02/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD02/u31  (\ADD01/ADD02/n18 , \ADD01/ADD02/n17 , \ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD02/u32  (\ADD01/ADD02/n19 , \ADD01/ADD02/n16 , \ADD01/ADD02/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD01/ADD02/u33  (temp_exp_diff[5], \ADD01/ADD02/p1 , \ADD01/ADD02/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD01/ADD02/u34  (temp_exp_diff[4], \ADD01/ADD02/p0 , \ADD01/ctemp );  // ../RTL/core/fpu_utils.v(71)
  and \ADD01/ADD02/u35  (\ADD01/ADD02/n20 , \ADD01/ADD02/n17 , \ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD01/ADD02/u36  (\ADD01/ADD02/n21 , \ADD01/ADD02/n20 , \ADD01/ctemp );  // ../RTL/core/fpu_utils.v(66)
  or \ADD01/ADD02/u37  (isE1GreaterThanE2, \ADD01/ADD02/n19 , \ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD01/ADD02/u4  (\ADD01/ADD02/p0 , n1[27], complemented_E2[4]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD01/ADD02/u5  (\ADD01/ADD02/p1 , n1[28], complemented_E2[5]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD01/ADD02/u6  (\ADD01/ADD02/p2 , n1[29], complemented_E2[6]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD01/ADD02/u7  (\ADD01/ADD02/p3 , n1[30], complemented_E2[7]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD01/ADD02/u8  (\ADD01/ADD02/n0 , \ADD01/ADD02/p0 , \ADD01/ctemp );  // ../RTL/core/fpu_utils.v(63)
  or \ADD01/ADD02/u9  (\ADD01/ADD02/c0 , \ADD01/ADD02/g0 , \ADD01/ADD02/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD02/ADD01/ADD01/u0  (\ADD02/ADD01/ADD01/g0 , M1[0], new_M2[0]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD02/ADD01/ADD01/u1  (\ADD02/ADD01/ADD01/g1 , M1[1], new_M2[1]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD02/ADD01/ADD01/u10  (\ADD02/ADD01/ADD01/n1 , \ADD02/ADD01/ADD01/p1 , \ADD02/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD01/ADD01/u11  (\ADD02/ADD01/ADD01/n2 , \ADD02/ADD01/ADD01/g1 , \ADD02/ADD01/ADD01/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD01/ADD01/u12  (\ADD02/ADD01/ADD01/n3 , \ADD02/ADD01/ADD01/p1 , \ADD02/ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD01/ADD01/u13  (\ADD02/ADD01/ADD01/n4 , \ADD02/ADD01/ADD01/n3 , real_oper);  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD01/ADD01/u14  (\ADD02/ADD01/ADD01/c1 , \ADD02/ADD01/ADD01/n2 , \ADD02/ADD01/ADD01/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD01/ADD01/u15  (\ADD02/ADD01/ADD01/n5 , \ADD02/ADD01/ADD01/p2 , \ADD02/ADD01/ADD01/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD01/ADD01/u16  (\ADD02/ADD01/ADD01/n6 , \ADD02/ADD01/ADD01/g2 , \ADD02/ADD01/ADD01/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD01/u17  (\ADD02/ADD01/ADD01/n7 , \ADD02/ADD01/ADD01/p2 , \ADD02/ADD01/ADD01/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD01/u18  (\ADD02/ADD01/ADD01/n8 , \ADD02/ADD01/ADD01/n7 , \ADD02/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD01/ADD01/u19  (\ADD02/ADD01/ADD01/n9 , \ADD02/ADD01/ADD01/n6 , \ADD02/ADD01/ADD01/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD01/u2  (\ADD02/ADD01/ADD01/g2 , M1[2], new_M2[2]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD02/ADD01/ADD01/u20  (M_result[3], \ADD02/ADD01/ADD01/p3 , \ADD02/ADD01/ADD01/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD01/ADD01/u21  (\ADD02/ADD01/ADD01/n10 , \ADD02/ADD01/ADD01/n7 , \ADD02/ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD01/u22  (\ADD02/ADD01/ADD01/n11 , \ADD02/ADD01/ADD01/n10 , real_oper);  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD01/ADD01/u23  (\ADD02/ADD01/ADD01/c2 , \ADD02/ADD01/ADD01/n9 , \ADD02/ADD01/ADD01/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD01/u24  (\ADD02/ADD01/ADD01/n12 , \ADD02/ADD01/ADD01/p3 , \ADD02/ADD01/ADD01/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD01/u25  (\ADD02/ADD01/ADD01/n13 , \ADD02/ADD01/ADD01/g3 , \ADD02/ADD01/ADD01/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD01/u26  (\ADD02/ADD01/ADD01/n14 , \ADD02/ADD01/ADD01/p3 , \ADD02/ADD01/ADD01/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD01/u27  (\ADD02/ADD01/ADD01/n15 , \ADD02/ADD01/ADD01/n14 , \ADD02/ADD01/ADD01/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD01/u28  (\ADD02/ADD01/ADD01/n16 , \ADD02/ADD01/ADD01/n13 , \ADD02/ADD01/ADD01/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD01/ADD01/u29  (M_result[2], \ADD02/ADD01/ADD01/p2 , \ADD02/ADD01/ADD01/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD01/ADD01/u3  (\ADD02/ADD01/ADD01/g3 , M1[3], new_M2[3]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD02/ADD01/ADD01/u30  (\ADD02/ADD01/ADD01/n17 , \ADD02/ADD01/ADD01/n14 , \ADD02/ADD01/ADD01/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD01/u31  (\ADD02/ADD01/ADD01/n18 , \ADD02/ADD01/ADD01/n17 , \ADD02/ADD01/ADD01/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD01/u32  (\ADD02/ADD01/ADD01/n19 , \ADD02/ADD01/ADD01/n16 , \ADD02/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD01/ADD01/u33  (M_result[1], \ADD02/ADD01/ADD01/p1 , \ADD02/ADD01/ADD01/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD02/ADD01/ADD01/u34  (M_result[0], \ADD02/ADD01/ADD01/p0 , real_oper);  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD01/ADD01/u35  (\ADD02/ADD01/ADD01/n20 , \ADD02/ADD01/ADD01/n17 , \ADD02/ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD01/u36  (\ADD02/ADD01/ADD01/n21 , \ADD02/ADD01/ADD01/n20 , real_oper);  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD01/u37  (\ADD02/ADD01/ctemp , \ADD02/ADD01/ADD01/n19 , \ADD02/ADD01/ADD01/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD01/ADD01/u4  (\ADD02/ADD01/ADD01/p0 , M1[0], new_M2[0]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD02/ADD01/ADD01/u5  (\ADD02/ADD01/ADD01/p1 , M1[1], new_M2[1]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD02/ADD01/ADD01/u6  (\ADD02/ADD01/ADD01/p2 , M1[2], new_M2[2]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD02/ADD01/ADD01/u7  (\ADD02/ADD01/ADD01/p3 , M1[3], new_M2[3]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD02/ADD01/ADD01/u8  (\ADD02/ADD01/ADD01/n0 , \ADD02/ADD01/ADD01/p0 , real_oper);  // ../RTL/core/fpu_utils.v(63)
  or \ADD02/ADD01/ADD01/u9  (\ADD02/ADD01/ADD01/c0 , \ADD02/ADD01/ADD01/g0 , \ADD02/ADD01/ADD01/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD02/ADD01/ADD02/u0  (\ADD02/ADD01/ADD02/g0 , M1[4], new_M2[4]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD02/ADD01/ADD02/u1  (\ADD02/ADD01/ADD02/g1 , M1[5], new_M2[5]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD02/ADD01/ADD02/u10  (\ADD02/ADD01/ADD02/n1 , \ADD02/ADD01/ADD02/p1 , \ADD02/ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD01/ADD02/u11  (\ADD02/ADD01/ADD02/n2 , \ADD02/ADD01/ADD02/g1 , \ADD02/ADD01/ADD02/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD01/ADD02/u12  (\ADD02/ADD01/ADD02/n3 , \ADD02/ADD01/ADD02/p1 , \ADD02/ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD01/ADD02/u13  (\ADD02/ADD01/ADD02/n4 , \ADD02/ADD01/ADD02/n3 , \ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD01/ADD02/u14  (\ADD02/ADD01/ADD02/c1 , \ADD02/ADD01/ADD02/n2 , \ADD02/ADD01/ADD02/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD01/ADD02/u15  (\ADD02/ADD01/ADD02/n5 , \ADD02/ADD01/ADD02/p2 , \ADD02/ADD01/ADD02/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD01/ADD02/u16  (\ADD02/ADD01/ADD02/n6 , \ADD02/ADD01/ADD02/g2 , \ADD02/ADD01/ADD02/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD02/u17  (\ADD02/ADD01/ADD02/n7 , \ADD02/ADD01/ADD02/p2 , \ADD02/ADD01/ADD02/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD02/u18  (\ADD02/ADD01/ADD02/n8 , \ADD02/ADD01/ADD02/n7 , \ADD02/ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD01/ADD02/u19  (\ADD02/ADD01/ADD02/n9 , \ADD02/ADD01/ADD02/n6 , \ADD02/ADD01/ADD02/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD02/u2  (\ADD02/ADD01/ADD02/g2 , M1[6], new_M2[6]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD02/ADD01/ADD02/u20  (M_result[7], \ADD02/ADD01/ADD02/p3 , \ADD02/ADD01/ADD02/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD01/ADD02/u21  (\ADD02/ADD01/ADD02/n10 , \ADD02/ADD01/ADD02/n7 , \ADD02/ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD02/u22  (\ADD02/ADD01/ADD02/n11 , \ADD02/ADD01/ADD02/n10 , \ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD01/ADD02/u23  (\ADD02/ADD01/ADD02/c2 , \ADD02/ADD01/ADD02/n9 , \ADD02/ADD01/ADD02/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD01/ADD02/u24  (\ADD02/ADD01/ADD02/n12 , \ADD02/ADD01/ADD02/p3 , \ADD02/ADD01/ADD02/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD02/u25  (\ADD02/ADD01/ADD02/n13 , \ADD02/ADD01/ADD02/g3 , \ADD02/ADD01/ADD02/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD02/u26  (\ADD02/ADD01/ADD02/n14 , \ADD02/ADD01/ADD02/p3 , \ADD02/ADD01/ADD02/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD02/u27  (\ADD02/ADD01/ADD02/n15 , \ADD02/ADD01/ADD02/n14 , \ADD02/ADD01/ADD02/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD02/u28  (\ADD02/ADD01/ADD02/n16 , \ADD02/ADD01/ADD02/n13 , \ADD02/ADD01/ADD02/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD01/ADD02/u29  (M_result[6], \ADD02/ADD01/ADD02/p2 , \ADD02/ADD01/ADD02/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD01/ADD02/u3  (\ADD02/ADD01/ADD02/g3 , M1[7], new_M2[7]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD02/ADD01/ADD02/u30  (\ADD02/ADD01/ADD02/n17 , \ADD02/ADD01/ADD02/n14 , \ADD02/ADD01/ADD02/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD02/u31  (\ADD02/ADD01/ADD02/n18 , \ADD02/ADD01/ADD02/n17 , \ADD02/ADD01/ADD02/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD02/u32  (\ADD02/ADD01/ADD02/n19 , \ADD02/ADD01/ADD02/n16 , \ADD02/ADD01/ADD02/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD01/ADD02/u33  (M_result[5], \ADD02/ADD01/ADD02/p1 , \ADD02/ADD01/ADD02/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD02/ADD01/ADD02/u34  (M_result[4], \ADD02/ADD01/ADD02/p0 , \ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD01/ADD02/u35  (\ADD02/ADD01/ADD02/n20 , \ADD02/ADD01/ADD02/n17 , \ADD02/ADD01/ADD02/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD01/ADD02/u36  (\ADD02/ADD01/ADD02/n21 , \ADD02/ADD01/ADD02/n20 , \ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD01/ADD02/u37  (\ADD02/ctemp1 , \ADD02/ADD01/ADD02/n19 , \ADD02/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD01/ADD02/u4  (\ADD02/ADD01/ADD02/p0 , M1[4], new_M2[4]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD02/ADD01/ADD02/u5  (\ADD02/ADD01/ADD02/p1 , M1[5], new_M2[5]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD02/ADD01/ADD02/u6  (\ADD02/ADD01/ADD02/p2 , M1[6], new_M2[6]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD02/ADD01/ADD02/u7  (\ADD02/ADD01/ADD02/p3 , M1[7], new_M2[7]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD02/ADD01/ADD02/u8  (\ADD02/ADD01/ADD02/n0 , \ADD02/ADD01/ADD02/p0 , \ADD02/ADD01/ctemp );  // ../RTL/core/fpu_utils.v(63)
  or \ADD02/ADD01/ADD02/u9  (\ADD02/ADD01/ADD02/c0 , \ADD02/ADD01/ADD02/g0 , \ADD02/ADD01/ADD02/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD02/ADD02/ADD01/u0  (\ADD02/ADD02/ADD01/g0 , M1[8], new_M2[8]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD02/ADD02/ADD01/u1  (\ADD02/ADD02/ADD01/g1 , M1[9], new_M2[9]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD02/ADD02/ADD01/u10  (\ADD02/ADD02/ADD01/n1 , \ADD02/ADD02/ADD01/p1 , \ADD02/ADD02/ADD01/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD02/ADD01/u11  (\ADD02/ADD02/ADD01/n2 , \ADD02/ADD02/ADD01/g1 , \ADD02/ADD02/ADD01/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD02/ADD01/u12  (\ADD02/ADD02/ADD01/n3 , \ADD02/ADD02/ADD01/p1 , \ADD02/ADD02/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD02/ADD01/u13  (\ADD02/ADD02/ADD01/n4 , \ADD02/ADD02/ADD01/n3 , \ADD02/ctemp1 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD02/ADD01/u14  (\ADD02/ADD02/ADD01/c1 , \ADD02/ADD02/ADD01/n2 , \ADD02/ADD02/ADD01/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD02/ADD01/u15  (\ADD02/ADD02/ADD01/n5 , \ADD02/ADD02/ADD01/p2 , \ADD02/ADD02/ADD01/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD02/ADD01/u16  (\ADD02/ADD02/ADD01/n6 , \ADD02/ADD02/ADD01/g2 , \ADD02/ADD02/ADD01/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD01/u17  (\ADD02/ADD02/ADD01/n7 , \ADD02/ADD02/ADD01/p2 , \ADD02/ADD02/ADD01/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD01/u18  (\ADD02/ADD02/ADD01/n8 , \ADD02/ADD02/ADD01/n7 , \ADD02/ADD02/ADD01/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD02/ADD01/u19  (\ADD02/ADD02/ADD01/n9 , \ADD02/ADD02/ADD01/n6 , \ADD02/ADD02/ADD01/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD01/u2  (\ADD02/ADD02/ADD01/g2 , M1[10], new_M2[10]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD02/ADD02/ADD01/u20  (M_result[11], \ADD02/ADD02/ADD01/p3 , \ADD02/ADD02/ADD01/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD02/ADD01/u21  (\ADD02/ADD02/ADD01/n10 , \ADD02/ADD02/ADD01/n7 , \ADD02/ADD02/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD01/u22  (\ADD02/ADD02/ADD01/n11 , \ADD02/ADD02/ADD01/n10 , \ADD02/ctemp1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD02/ADD01/u23  (\ADD02/ADD02/ADD01/c2 , \ADD02/ADD02/ADD01/n9 , \ADD02/ADD02/ADD01/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD01/u24  (\ADD02/ADD02/ADD01/n12 , \ADD02/ADD02/ADD01/p3 , \ADD02/ADD02/ADD01/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD01/u25  (\ADD02/ADD02/ADD01/n13 , \ADD02/ADD02/ADD01/g3 , \ADD02/ADD02/ADD01/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD01/u26  (\ADD02/ADD02/ADD01/n14 , \ADD02/ADD02/ADD01/p3 , \ADD02/ADD02/ADD01/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD01/u27  (\ADD02/ADD02/ADD01/n15 , \ADD02/ADD02/ADD01/n14 , \ADD02/ADD02/ADD01/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD01/u28  (\ADD02/ADD02/ADD01/n16 , \ADD02/ADD02/ADD01/n13 , \ADD02/ADD02/ADD01/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD02/ADD01/u29  (M_result[10], \ADD02/ADD02/ADD01/p2 , \ADD02/ADD02/ADD01/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD02/ADD01/u3  (\ADD02/ADD02/ADD01/g3 , M1[11], new_M2[11]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD02/ADD02/ADD01/u30  (\ADD02/ADD02/ADD01/n17 , \ADD02/ADD02/ADD01/n14 , \ADD02/ADD02/ADD01/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD01/u31  (\ADD02/ADD02/ADD01/n18 , \ADD02/ADD02/ADD01/n17 , \ADD02/ADD02/ADD01/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD01/u32  (\ADD02/ADD02/ADD01/n19 , \ADD02/ADD02/ADD01/n16 , \ADD02/ADD02/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD02/ADD01/u33  (M_result[9], \ADD02/ADD02/ADD01/p1 , \ADD02/ADD02/ADD01/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD02/ADD02/ADD01/u34  (M_result[8], \ADD02/ADD02/ADD01/p0 , \ADD02/ctemp1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD02/ADD01/u35  (\ADD02/ADD02/ADD01/n20 , \ADD02/ADD02/ADD01/n17 , \ADD02/ADD02/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD01/u36  (\ADD02/ADD02/ADD01/n21 , \ADD02/ADD02/ADD01/n20 , \ADD02/ctemp1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD01/u37  (\ADD02/ADD02/ctemp , \ADD02/ADD02/ADD01/n19 , \ADD02/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD02/ADD01/u4  (\ADD02/ADD02/ADD01/p0 , M1[8], new_M2[8]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD02/ADD02/ADD01/u5  (\ADD02/ADD02/ADD01/p1 , M1[9], new_M2[9]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD02/ADD02/ADD01/u6  (\ADD02/ADD02/ADD01/p2 , M1[10], new_M2[10]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD02/ADD02/ADD01/u7  (\ADD02/ADD02/ADD01/p3 , M1[11], new_M2[11]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD02/ADD02/ADD01/u8  (\ADD02/ADD02/ADD01/n0 , \ADD02/ADD02/ADD01/p0 , \ADD02/ctemp1 );  // ../RTL/core/fpu_utils.v(63)
  or \ADD02/ADD02/ADD01/u9  (\ADD02/ADD02/ADD01/c0 , \ADD02/ADD02/ADD01/g0 , \ADD02/ADD02/ADD01/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD02/ADD02/ADD02/u0  (\ADD02/ADD02/ADD02/g0 , M1[12], new_M2[12]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD02/ADD02/ADD02/u1  (\ADD02/ADD02/ADD02/g1 , M1[13], new_M2[13]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD02/ADD02/ADD02/u10  (\ADD02/ADD02/ADD02/n1 , \ADD02/ADD02/ADD02/p1 , \ADD02/ADD02/ADD02/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD02/ADD02/u11  (\ADD02/ADD02/ADD02/n2 , \ADD02/ADD02/ADD02/g1 , \ADD02/ADD02/ADD02/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD02/ADD02/u12  (\ADD02/ADD02/ADD02/n3 , \ADD02/ADD02/ADD02/p1 , \ADD02/ADD02/ADD02/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD02/ADD02/u13  (\ADD02/ADD02/ADD02/n4 , \ADD02/ADD02/ADD02/n3 , \ADD02/ADD02/ctemp );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD02/ADD02/u14  (\ADD02/ADD02/ADD02/c1 , \ADD02/ADD02/ADD02/n2 , \ADD02/ADD02/ADD02/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD02/ADD02/u15  (\ADD02/ADD02/ADD02/n5 , \ADD02/ADD02/ADD02/p2 , \ADD02/ADD02/ADD02/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD02/ADD02/u16  (\ADD02/ADD02/ADD02/n6 , \ADD02/ADD02/ADD02/g2 , \ADD02/ADD02/ADD02/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD02/u17  (\ADD02/ADD02/ADD02/n7 , \ADD02/ADD02/ADD02/p2 , \ADD02/ADD02/ADD02/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD02/u18  (\ADD02/ADD02/ADD02/n8 , \ADD02/ADD02/ADD02/n7 , \ADD02/ADD02/ADD02/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD02/ADD02/u19  (\ADD02/ADD02/ADD02/n9 , \ADD02/ADD02/ADD02/n6 , \ADD02/ADD02/ADD02/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD02/u2  (\ADD02/ADD02/ADD02/g2 , M1[14], new_M2[14]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD02/ADD02/ADD02/u20  (M_result[15], \ADD02/ADD02/ADD02/p3 , \ADD02/ADD02/ADD02/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD02/ADD02/u21  (\ADD02/ADD02/ADD02/n10 , \ADD02/ADD02/ADD02/n7 , \ADD02/ADD02/ADD02/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD02/u22  (\ADD02/ADD02/ADD02/n11 , \ADD02/ADD02/ADD02/n10 , \ADD02/ADD02/ctemp );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD02/ADD02/u23  (\ADD02/ADD02/ADD02/c2 , \ADD02/ADD02/ADD02/n9 , \ADD02/ADD02/ADD02/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD02/ADD02/u24  (\ADD02/ADD02/ADD02/n12 , \ADD02/ADD02/ADD02/p3 , \ADD02/ADD02/ADD02/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD02/u25  (\ADD02/ADD02/ADD02/n13 , \ADD02/ADD02/ADD02/g3 , \ADD02/ADD02/ADD02/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD02/u26  (\ADD02/ADD02/ADD02/n14 , \ADD02/ADD02/ADD02/p3 , \ADD02/ADD02/ADD02/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD02/u27  (\ADD02/ADD02/ADD02/n15 , \ADD02/ADD02/ADD02/n14 , \ADD02/ADD02/ADD02/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD02/u28  (\ADD02/ADD02/ADD02/n16 , \ADD02/ADD02/ADD02/n13 , \ADD02/ADD02/ADD02/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD02/ADD02/u29  (M_result[14], \ADD02/ADD02/ADD02/p2 , \ADD02/ADD02/ADD02/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD02/ADD02/u3  (\ADD02/ADD02/ADD02/g3 , M1[15], new_M2[15]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD02/ADD02/ADD02/u30  (\ADD02/ADD02/ADD02/n17 , \ADD02/ADD02/ADD02/n14 , \ADD02/ADD02/ADD02/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD02/u31  (\ADD02/ADD02/ADD02/n18 , \ADD02/ADD02/ADD02/n17 , \ADD02/ADD02/ADD02/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD02/u32  (\ADD02/ADD02/ADD02/n19 , \ADD02/ADD02/ADD02/n16 , \ADD02/ADD02/ADD02/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD02/ADD02/u33  (M_result[13], \ADD02/ADD02/ADD02/p1 , \ADD02/ADD02/ADD02/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD02/ADD02/ADD02/u34  (M_result[12], \ADD02/ADD02/ADD02/p0 , \ADD02/ADD02/ctemp );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD02/ADD02/u35  (\ADD02/ADD02/ADD02/n20 , \ADD02/ADD02/ADD02/n17 , \ADD02/ADD02/ADD02/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD02/ADD02/u36  (\ADD02/ADD02/ADD02/n21 , \ADD02/ADD02/ADD02/n20 , \ADD02/ADD02/ctemp );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD02/ADD02/u37  (\ADD02/ctemp2 , \ADD02/ADD02/ADD02/n19 , \ADD02/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD02/ADD02/u4  (\ADD02/ADD02/ADD02/p0 , M1[12], new_M2[12]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD02/ADD02/ADD02/u5  (\ADD02/ADD02/ADD02/p1 , M1[13], new_M2[13]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD02/ADD02/ADD02/u6  (\ADD02/ADD02/ADD02/p2 , M1[14], new_M2[14]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD02/ADD02/ADD02/u7  (\ADD02/ADD02/ADD02/p3 , M1[15], new_M2[15]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD02/ADD02/ADD02/u8  (\ADD02/ADD02/ADD02/n0 , \ADD02/ADD02/ADD02/p0 , \ADD02/ADD02/ctemp );  // ../RTL/core/fpu_utils.v(63)
  or \ADD02/ADD02/ADD02/u9  (\ADD02/ADD02/ADD02/c0 , \ADD02/ADD02/ADD02/g0 , \ADD02/ADD02/ADD02/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD02/ADD03/ADD01/u0  (\ADD02/ADD03/ADD01/g0 , M1[16], new_M2[16]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD02/ADD03/ADD01/u1  (\ADD02/ADD03/ADD01/g1 , M1[17], new_M2[17]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD02/ADD03/ADD01/u10  (\ADD02/ADD03/ADD01/n1 , \ADD02/ADD03/ADD01/p1 , \ADD02/ADD03/ADD01/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD03/ADD01/u11  (\ADD02/ADD03/ADD01/n2 , \ADD02/ADD03/ADD01/g1 , \ADD02/ADD03/ADD01/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD03/ADD01/u12  (\ADD02/ADD03/ADD01/n3 , \ADD02/ADD03/ADD01/p1 , \ADD02/ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD03/ADD01/u13  (\ADD02/ADD03/ADD01/n4 , \ADD02/ADD03/ADD01/n3 , \ADD02/ctemp2 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD03/ADD01/u14  (\ADD02/ADD03/ADD01/c1 , \ADD02/ADD03/ADD01/n2 , \ADD02/ADD03/ADD01/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD03/ADD01/u15  (\ADD02/ADD03/ADD01/n5 , \ADD02/ADD03/ADD01/p2 , \ADD02/ADD03/ADD01/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD03/ADD01/u16  (\ADD02/ADD03/ADD01/n6 , \ADD02/ADD03/ADD01/g2 , \ADD02/ADD03/ADD01/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD01/u17  (\ADD02/ADD03/ADD01/n7 , \ADD02/ADD03/ADD01/p2 , \ADD02/ADD03/ADD01/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD01/u18  (\ADD02/ADD03/ADD01/n8 , \ADD02/ADD03/ADD01/n7 , \ADD02/ADD03/ADD01/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD03/ADD01/u19  (\ADD02/ADD03/ADD01/n9 , \ADD02/ADD03/ADD01/n6 , \ADD02/ADD03/ADD01/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD01/u2  (\ADD02/ADD03/ADD01/g2 , M1[18], new_M2[18]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD02/ADD03/ADD01/u20  (M_result[19], \ADD02/ADD03/ADD01/p3 , \ADD02/ADD03/ADD01/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD03/ADD01/u21  (\ADD02/ADD03/ADD01/n10 , \ADD02/ADD03/ADD01/n7 , \ADD02/ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD01/u22  (\ADD02/ADD03/ADD01/n11 , \ADD02/ADD03/ADD01/n10 , \ADD02/ctemp2 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD03/ADD01/u23  (\ADD02/ADD03/ADD01/c2 , \ADD02/ADD03/ADD01/n9 , \ADD02/ADD03/ADD01/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD01/u24  (\ADD02/ADD03/ADD01/n12 , \ADD02/ADD03/ADD01/p3 , \ADD02/ADD03/ADD01/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD01/u25  (\ADD02/ADD03/ADD01/n13 , \ADD02/ADD03/ADD01/g3 , \ADD02/ADD03/ADD01/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD01/u26  (\ADD02/ADD03/ADD01/n14 , \ADD02/ADD03/ADD01/p3 , \ADD02/ADD03/ADD01/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD01/u27  (\ADD02/ADD03/ADD01/n15 , \ADD02/ADD03/ADD01/n14 , \ADD02/ADD03/ADD01/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD01/u28  (\ADD02/ADD03/ADD01/n16 , \ADD02/ADD03/ADD01/n13 , \ADD02/ADD03/ADD01/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD03/ADD01/u29  (M_result[18], \ADD02/ADD03/ADD01/p2 , \ADD02/ADD03/ADD01/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD03/ADD01/u3  (\ADD02/ADD03/ADD01/g3 , M1[19], new_M2[19]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD02/ADD03/ADD01/u30  (\ADD02/ADD03/ADD01/n17 , \ADD02/ADD03/ADD01/n14 , \ADD02/ADD03/ADD01/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD01/u31  (\ADD02/ADD03/ADD01/n18 , \ADD02/ADD03/ADD01/n17 , \ADD02/ADD03/ADD01/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD01/u32  (\ADD02/ADD03/ADD01/n19 , \ADD02/ADD03/ADD01/n16 , \ADD02/ADD03/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD03/ADD01/u33  (M_result[17], \ADD02/ADD03/ADD01/p1 , \ADD02/ADD03/ADD01/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD02/ADD03/ADD01/u34  (M_result[16], \ADD02/ADD03/ADD01/p0 , \ADD02/ctemp2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD03/ADD01/u35  (\ADD02/ADD03/ADD01/n20 , \ADD02/ADD03/ADD01/n17 , \ADD02/ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD01/u36  (\ADD02/ADD03/ADD01/n21 , \ADD02/ADD03/ADD01/n20 , \ADD02/ctemp2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD01/u37  (\ADD02/ADD03/ctemp , \ADD02/ADD03/ADD01/n19 , \ADD02/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD03/ADD01/u4  (\ADD02/ADD03/ADD01/p0 , M1[16], new_M2[16]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD02/ADD03/ADD01/u5  (\ADD02/ADD03/ADD01/p1 , M1[17], new_M2[17]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD02/ADD03/ADD01/u6  (\ADD02/ADD03/ADD01/p2 , M1[18], new_M2[18]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD02/ADD03/ADD01/u7  (\ADD02/ADD03/ADD01/p3 , M1[19], new_M2[19]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD02/ADD03/ADD01/u8  (\ADD02/ADD03/ADD01/n0 , \ADD02/ADD03/ADD01/p0 , \ADD02/ctemp2 );  // ../RTL/core/fpu_utils.v(63)
  or \ADD02/ADD03/ADD01/u9  (\ADD02/ADD03/ADD01/c0 , \ADD02/ADD03/ADD01/g0 , \ADD02/ADD03/ADD01/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD02/ADD03/ADD02/u0  (\ADD02/ADD03/ADD02/g0 , M1[20], new_M2[20]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD02/ADD03/ADD02/u1  (\ADD02/ADD03/ADD02/g1 , M1[21], new_M2[21]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD02/ADD03/ADD02/u10  (\ADD02/ADD03/ADD02/n1 , \ADD02/ADD03/ADD02/p1 , \ADD02/ADD03/ADD02/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD03/ADD02/u11  (\ADD02/ADD03/ADD02/n2 , \ADD02/ADD03/ADD02/g1 , \ADD02/ADD03/ADD02/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD03/ADD02/u12  (\ADD02/ADD03/ADD02/n3 , \ADD02/ADD03/ADD02/p1 , \ADD02/ADD03/ADD02/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD03/ADD02/u13  (\ADD02/ADD03/ADD02/n4 , \ADD02/ADD03/ADD02/n3 , \ADD02/ADD03/ctemp );  // ../RTL/core/fpu_utils.v(64)
  or \ADD02/ADD03/ADD02/u14  (\ADD02/ADD03/ADD02/c1 , \ADD02/ADD03/ADD02/n2 , \ADD02/ADD03/ADD02/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD02/ADD03/ADD02/u15  (\ADD02/ADD03/ADD02/n5 , \ADD02/ADD03/ADD02/p2 , \ADD02/ADD03/ADD02/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD03/ADD02/u16  (\ADD02/ADD03/ADD02/n6 , \ADD02/ADD03/ADD02/g2 , \ADD02/ADD03/ADD02/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD02/u17  (\ADD02/ADD03/ADD02/n7 , \ADD02/ADD03/ADD02/p2 , \ADD02/ADD03/ADD02/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD02/u18  (\ADD02/ADD03/ADD02/n8 , \ADD02/ADD03/ADD02/n7 , \ADD02/ADD03/ADD02/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD03/ADD02/u19  (\ADD02/ADD03/ADD02/n9 , \ADD02/ADD03/ADD02/n6 , \ADD02/ADD03/ADD02/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD02/u2  (\ADD02/ADD03/ADD02/g2 , M1[22], new_M2[22]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD02/ADD03/ADD02/u20  (M_result[23], \ADD02/ADD03/ADD02/p3 , \ADD02/ADD03/ADD02/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD03/ADD02/u21  (\ADD02/ADD03/ADD02/n10 , \ADD02/ADD03/ADD02/n7 , \ADD02/ADD03/ADD02/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD02/u22  (\ADD02/ADD03/ADD02/n11 , \ADD02/ADD03/ADD02/n10 , \ADD02/ADD03/ctemp );  // ../RTL/core/fpu_utils.v(65)
  or \ADD02/ADD03/ADD02/u23  (\ADD02/ADD03/ADD02/c2 , \ADD02/ADD03/ADD02/n9 , \ADD02/ADD03/ADD02/n11 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD02/ADD03/ADD02/u24  (\ADD02/ADD03/ADD02/n12 , \ADD02/ADD03/ADD02/p3 , \ADD02/ADD03/ADD02/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD02/u25  (\ADD02/ADD03/ADD02/n13 , \ADD02/ADD03/ADD02/g3 , \ADD02/ADD03/ADD02/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD02/u26  (\ADD02/ADD03/ADD02/n14 , \ADD02/ADD03/ADD02/p3 , \ADD02/ADD03/ADD02/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD02/u27  (\ADD02/ADD03/ADD02/n15 , \ADD02/ADD03/ADD02/n14 , \ADD02/ADD03/ADD02/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD02/u28  (\ADD02/ADD03/ADD02/n16 , \ADD02/ADD03/ADD02/n13 , \ADD02/ADD03/ADD02/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD03/ADD02/u29  (M_result[22], \ADD02/ADD03/ADD02/p2 , \ADD02/ADD03/ADD02/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD03/ADD02/u3  (\ADD02/ADD03/ADD02/g3 , M1[23], new_M2[23]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD02/ADD03/ADD02/u30  (\ADD02/ADD03/ADD02/n17 , \ADD02/ADD03/ADD02/n14 , \ADD02/ADD03/ADD02/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD02/u31  (\ADD02/ADD03/ADD02/n18 , \ADD02/ADD03/ADD02/n17 , \ADD02/ADD03/ADD02/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD02/u32  (\ADD02/ADD03/ADD02/n19 , \ADD02/ADD03/ADD02/n16 , \ADD02/ADD03/ADD02/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD03/ADD02/u33  (M_result[21], \ADD02/ADD03/ADD02/p1 , \ADD02/ADD03/ADD02/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD02/ADD03/ADD02/u34  (M_result[20], \ADD02/ADD03/ADD02/p0 , \ADD02/ADD03/ctemp );  // ../RTL/core/fpu_utils.v(71)
  and \ADD02/ADD03/ADD02/u35  (\ADD02/ADD03/ADD02/n20 , \ADD02/ADD03/ADD02/n17 , \ADD02/ADD03/ADD02/p0 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD02/ADD03/ADD02/u36  (\ADD02/ADD03/ADD02/n21 , \ADD02/ADD03/ADD02/n20 , \ADD02/ADD03/ctemp );  // ../RTL/core/fpu_utils.v(66)
  or \ADD02/ADD03/ADD02/u37  (M_carry, \ADD02/ADD03/ADD02/n19 , \ADD02/ADD03/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD02/ADD03/ADD02/u4  (\ADD02/ADD03/ADD02/p0 , M1[20], new_M2[20]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD02/ADD03/ADD02/u5  (\ADD02/ADD03/ADD02/p1 , M1[21], new_M2[21]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD02/ADD03/ADD02/u6  (\ADD02/ADD03/ADD02/p2 , M1[22], new_M2[22]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD02/ADD03/ADD02/u7  (\ADD02/ADD03/ADD02/p3 , M1[23], new_M2[23]);  // ../RTL/core/fpu_utils.v(62)
  and \ADD02/ADD03/ADD02/u8  (\ADD02/ADD03/ADD02/n0 , \ADD02/ADD03/ADD02/p0 , \ADD02/ADD03/ctemp );  // ../RTL/core/fpu_utils.v(63)
  or \ADD02/ADD03/ADD02/u9  (\ADD02/ADD03/ADD02/c0 , \ADD02/ADD03/ADD02/g0 , \ADD02/ADD03/ADD02/n0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD0212/ADD01/u10  (\ADD0212/ADD01/n1 , E[1], E[0]);  // ../RTL/core/fpu_utils.v(64)
  and \ADD0212/ADD01/u17  (\ADD0212/ADD01/n7 , E[2], E[1]);  // ../RTL/core/fpu_utils.v(65)
  and \ADD0212/ADD01/u18  (\ADD0212/ADD01/n8 , \ADD0212/ADD01/n7 , E[0]);  // ../RTL/core/fpu_utils.v(65)
  xor \ADD0212/ADD01/u20  (One_Added_E[3], E[3], \ADD0212/ADD01/n8 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD0212/ADD01/u26  (\ADD0212/ADD01/n14 , E[3], E[2]);  // ../RTL/core/fpu_utils.v(66)
  xor \ADD0212/ADD01/u29  (One_Added_E[2], E[2], \ADD0212/ADD01/n1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD0212/ADD01/u30  (\ADD0212/ADD01/n17 , \ADD0212/ADD01/n14 , E[1]);  // ../RTL/core/fpu_utils.v(66)
  and \ADD0212/ADD01/u31  (\ADD0212/ADD01/n18 , \ADD0212/ADD01/n17 , E[0]);  // ../RTL/core/fpu_utils.v(66)
  xor \ADD0212/ADD01/u33  (One_Added_E[1], E[1], E[0]);  // ../RTL/core/fpu_utils.v(71)
  and \ADD0212/ADD02/u12  (\ADD0212/ADD02/n3 , E[5], E[4]);  // ../RTL/core/fpu_utils.v(64)
  and \ADD0212/ADD02/u13  (\ADD0212/ADD02/n4 , \ADD0212/ADD02/n3 , \ADD0212/ADD01/n18 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD0212/ADD02/u17  (\ADD0212/ADD02/n7 , E[6], E[5]);  // ../RTL/core/fpu_utils.v(65)
  xor \ADD0212/ADD02/u20  (One_Added_E[7], E[7], \ADD0212/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD0212/ADD02/u21  (\ADD0212/ADD02/n10 , \ADD0212/ADD02/n7 , E[4]);  // ../RTL/core/fpu_utils.v(65)
  and \ADD0212/ADD02/u22  (\ADD0212/ADD02/n11 , \ADD0212/ADD02/n10 , \ADD0212/ADD01/n18 );  // ../RTL/core/fpu_utils.v(65)
  xor \ADD0212/ADD02/u29  (One_Added_E[6], E[6], \ADD0212/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD0212/ADD02/u33  (One_Added_E[5], E[5], \ADD0212/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD0212/ADD02/u34  (One_Added_E[4], E[4], \ADD0212/ADD01/n18 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD0212/ADD02/u8  (\ADD0212/ADD02/n0 , E[4], \ADD0212/ADD01/n18 );  // ../RTL/core/fpu_utils.v(63)
  not \ADD03/ADD01/p0_inv  (\ADD03/ADD01/p0_neg , \ADD03/ADD01/p0 );
  and \ADD03/ADD01/u0  (\ADD03/ADD01/g0 , new_E[0], complemented_shift_E[0]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD03/ADD01/u1  (\ADD03/ADD01/g1 , new_E[1], complemented_shift_E[1]);  // ../RTL/core/fpu_utils.v(56)
  and \ADD03/ADD01/u10  (\ADD03/ADD01/n1 , \ADD03/ADD01/p1 , \ADD03/ADD01/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD03/ADD01/u11  (\ADD03/ADD01/n2 , \ADD03/ADD01/g1 , \ADD03/ADD01/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD03/ADD01/u12  (\ADD03/ADD01/n3 , \ADD03/ADD01/p1 , \ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD03/ADD01/u14  (\ADD03/ADD01/c1 , \ADD03/ADD01/n2 , \ADD03/ADD01/n3 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD03/ADD01/u15  (\ADD03/ADD01/n5 , \ADD03/ADD01/p2 , \ADD03/ADD01/g1 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD03/ADD01/u16  (\ADD03/ADD01/n6 , \ADD03/ADD01/g2 , \ADD03/ADD01/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD01/u17  (\ADD03/ADD01/n7 , \ADD03/ADD01/p2 , \ADD03/ADD01/p1 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD01/u18  (\ADD03/ADD01/n8 , \ADD03/ADD01/n7 , \ADD03/ADD01/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD03/ADD01/u19  (\ADD03/ADD01/n9 , \ADD03/ADD01/n6 , \ADD03/ADD01/n8 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD01/u2  (\ADD03/ADD01/g2 , new_E[2], complemented_shift_E[2]);  // ../RTL/core/fpu_utils.v(57)
  xor \ADD03/ADD01/u20  (result[26], \ADD03/ADD01/p3 , \ADD03/ADD01/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD03/ADD01/u21  (\ADD03/ADD01/n10 , \ADD03/ADD01/n7 , \ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD03/ADD01/u23  (\ADD03/ADD01/c2 , \ADD03/ADD01/n9 , \ADD03/ADD01/n10 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD01/u24  (\ADD03/ADD01/n12 , \ADD03/ADD01/p3 , \ADD03/ADD01/g2 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD03/ADD01/u25  (\ADD03/ADD01/n13 , \ADD03/ADD01/g3 , \ADD03/ADD01/n12 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD03/ADD01/u26  (\ADD03/ADD01/n14 , \ADD03/ADD01/p3 , \ADD03/ADD01/p2 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD03/ADD01/u27  (\ADD03/ADD01/n15 , \ADD03/ADD01/n14 , \ADD03/ADD01/g1 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD03/ADD01/u28  (\ADD03/ADD01/n16 , \ADD03/ADD01/n13 , \ADD03/ADD01/n15 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD03/ADD01/u29  (result[25], \ADD03/ADD01/p2 , \ADD03/ADD01/c1 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD03/ADD01/u3  (\ADD03/ADD01/g3 , new_E[3], complemented_shift_E[3]);  // ../RTL/core/fpu_utils.v(58)
  and \ADD03/ADD01/u30  (\ADD03/ADD01/n17 , \ADD03/ADD01/n14 , \ADD03/ADD01/p1 );  // ../RTL/core/fpu_utils.v(66)
  and \ADD03/ADD01/u31  (\ADD03/ADD01/n18 , \ADD03/ADD01/n17 , \ADD03/ADD01/g0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD03/ADD01/u32  (\ADD03/ADD01/n19 , \ADD03/ADD01/n16 , \ADD03/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD03/ADD01/u33  (result[24], \ADD03/ADD01/p1 , \ADD03/ADD01/c0 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD03/ADD01/u35  (\ADD03/ADD01/n20 , \ADD03/ADD01/n17 , \ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  or \ADD03/ADD01/u37  (\ADD03/ctemp , \ADD03/ADD01/n19 , \ADD03/ADD01/n20 );  // ../RTL/core/fpu_utils.v(66)
  xor \ADD03/ADD01/u4  (\ADD03/ADD01/p0 , new_E[0], complemented_shift_E[0]);  // ../RTL/core/fpu_utils.v(59)
  xor \ADD03/ADD01/u5  (\ADD03/ADD01/p1 , new_E[1], complemented_shift_E[1]);  // ../RTL/core/fpu_utils.v(60)
  xor \ADD03/ADD01/u6  (\ADD03/ADD01/p2 , new_E[2], complemented_shift_E[2]);  // ../RTL/core/fpu_utils.v(61)
  xor \ADD03/ADD01/u7  (\ADD03/ADD01/p3 , new_E[3], complemented_shift_E[3]);  // ../RTL/core/fpu_utils.v(62)
  or \ADD03/ADD01/u9  (\ADD03/ADD01/c0 , \ADD03/ADD01/g0 , \ADD03/ADD01/p0 );  // ../RTL/core/fpu_utils.v(63)
  and \ADD03/ADD02/u0  (\ADD03/ADD02/g0 , new_E[4], complemented_shift_E[4]);  // ../RTL/core/fpu_utils.v(55)
  and \ADD03/ADD02/u10  (\ADD03/ADD02/n1 , \new_E[5]_neg , \ADD03/ADD02/g0 );  // ../RTL/core/fpu_utils.v(64)
  or \ADD03/ADD02/u11  (\ADD03/ADD02/n2 , new_E[5], \ADD03/ADD02/n1 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD03/ADD02/u12  (\ADD03/ADD02/n3 , \new_E[5]_neg , \ADD03/ADD02/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD03/ADD02/u13  (\ADD03/ADD02/n4 , \ADD03/ADD02/n3 , \ADD03/ctemp );  // ../RTL/core/fpu_utils.v(64)
  or \ADD03/ADD02/u14  (\ADD03/ADD02/c1 , \ADD03/ADD02/n2 , \ADD03/ADD02/n4 );  // ../RTL/core/fpu_utils.v(64)
  and \ADD03/ADD02/u15  (\ADD03/ADD02/n5 , \new_E[6]_neg , new_E[5]);  // ../RTL/core/fpu_utils.v(65)
  or \ADD03/ADD02/u16  (\ADD03/ADD02/n6 , new_E[6], \ADD03/ADD02/n5 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD02/u17  (\ADD03/ADD02/n7 , \new_E[6]_neg , \new_E[5]_neg );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD02/u18  (\ADD03/ADD02/n8 , \ADD03/ADD02/n7 , \ADD03/ADD02/g0 );  // ../RTL/core/fpu_utils.v(65)
  or \ADD03/ADD02/u19  (\ADD03/ADD02/n9 , \ADD03/ADD02/n6 , \ADD03/ADD02/n8 );  // ../RTL/core/fpu_utils.v(65)
  xor \ADD03/ADD02/u20  (result[30], \new_E[7]_neg , \ADD03/ADD02/c2 );  // ../RTL/core/fpu_utils.v(71)
  and \ADD03/ADD02/u21  (\ADD03/ADD02/n10 , \ADD03/ADD02/n7 , \ADD03/ADD02/p0 );  // ../RTL/core/fpu_utils.v(65)
  and \ADD03/ADD02/u22  (\ADD03/ADD02/n11 , \ADD03/ADD02/n10 , \ADD03/ctemp );  // ../RTL/core/fpu_utils.v(65)
  or \ADD03/ADD02/u23  (\ADD03/ADD02/c2 , \ADD03/ADD02/n9 , \ADD03/ADD02/n11 );  // ../RTL/core/fpu_utils.v(65)
  xor \ADD03/ADD02/u29  (result[29], \new_E[6]_neg , \ADD03/ADD02/c1 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD03/ADD02/u33  (result[28], \new_E[5]_neg , \ADD03/ADD02/c0 );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD03/ADD02/u34  (result[27], \ADD03/ADD02/p0 , \ADD03/ctemp );  // ../RTL/core/fpu_utils.v(71)
  xor \ADD03/ADD02/u4  (\ADD03/ADD02/p0 , new_E[4], complemented_shift_E[4]);  // ../RTL/core/fpu_utils.v(59)
  and \ADD03/ADD02/u8  (\ADD03/ADD02/n0 , \ADD03/ADD02/p0 , \ADD03/ctemp );  // ../RTL/core/fpu_utils.v(63)
  or \ADD03/ADD02/u9  (\ADD03/ADD02/c0 , \ADD03/ADD02/g0 , \ADD03/ADD02/n0 );  // ../RTL/core/fpu_utils.v(63)
  not \C01/u0  (complemented_E2[3], n2[26]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u1  (complemented_E2[2], n2[25]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u2  (complemented_E2[1], n2[24]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u3  (complemented_E2[0], n2[23]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u4  (complemented_E2[7], n2[30]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u5  (complemented_E2[6], n2[29]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u6  (complemented_E2[5], n2[28]);  // ../RTL/core/fpu_utils.v(44)
  not \C01/u7  (complemented_E2[4], n2[27]);  // ../RTL/core/fpu_utils.v(44)
  and \C023/ADD01/ADD01/u10  (\C023/ADD01/ADD01/n1 , \C023/outtemp [1], \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(64)
  and \C023/ADD01/ADD01/u17  (\C023/ADD01/ADD01/n7 , \C023/outtemp [2], \C023/outtemp [1]);  // ../RTL/core/fpu_utils.v(65)
  and \C023/ADD01/ADD01/u18  (\C023/ADD01/ADD01/n8 , \C023/ADD01/ADD01/n7 , \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(65)
  xor \C023/ADD01/ADD01/u20  (complemented_temp_exp_diff[3], \C023/outtemp [3], \C023/ADD01/ADD01/n8 );  // ../RTL/core/fpu_utils.v(71)
  and \C023/ADD01/ADD01/u26  (\C023/ADD01/ADD01/n14 , \C023/outtemp [3], \C023/outtemp [2]);  // ../RTL/core/fpu_utils.v(66)
  xor \C023/ADD01/ADD01/u29  (complemented_temp_exp_diff[2], \C023/outtemp [2], \C023/ADD01/ADD01/n1 );  // ../RTL/core/fpu_utils.v(71)
  and \C023/ADD01/ADD01/u30  (\C023/ADD01/ADD01/n17 , \C023/ADD01/ADD01/n14 , \C023/outtemp [1]);  // ../RTL/core/fpu_utils.v(66)
  and \C023/ADD01/ADD01/u31  (\C023/ADD01/ADD01/n18 , \C023/ADD01/ADD01/n17 , \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(66)
  xor \C023/ADD01/ADD01/u33  (complemented_temp_exp_diff[1], \C023/outtemp [1], \ADD01/ADD01/p0 );  // ../RTL/core/fpu_utils.v(71)
  and \C023/ADD01/ADD02/u12  (\C023/ADD01/ADD02/n3 , \C023/outtemp [5], \C023/outtemp [4]);  // ../RTL/core/fpu_utils.v(64)
  and \C023/ADD01/ADD02/u13  (\C023/ADD01/ADD02/n4 , \C023/ADD01/ADD02/n3 , \C023/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(64)
  and \C023/ADD01/ADD02/u17  (\C023/ADD01/ADD02/n7 , \C023/outtemp [6], \C023/outtemp [5]);  // ../RTL/core/fpu_utils.v(65)
  xor \C023/ADD01/ADD02/u20  (complemented_temp_exp_diff[7], \C023/outtemp [7], \C023/ADD01/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \C023/ADD01/ADD02/u21  (\C023/ADD01/ADD02/n10 , \C023/ADD01/ADD02/n7 , \C023/outtemp [4]);  // ../RTL/core/fpu_utils.v(65)
  and \C023/ADD01/ADD02/u22  (\C023/ADD01/ADD02/n11 , \C023/ADD01/ADD02/n10 , \C023/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(65)
  xor \C023/ADD01/ADD02/u29  (complemented_temp_exp_diff[6], \C023/outtemp [6], \C023/ADD01/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  xor \C023/ADD01/ADD02/u33  (complemented_temp_exp_diff[5], \C023/outtemp [5], \C023/ADD01/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \C023/ADD01/ADD02/u34  (complemented_temp_exp_diff[4], \C023/outtemp [4], \C023/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(71)
  and \C023/ADD01/ADD02/u8  (\C023/ADD01/ADD02/n0 , \C023/outtemp [4], \C023/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(63)
  not \C023/C01/u0  (\C023/outtemp [3], temp_exp_diff[3]);  // ../RTL/core/fpu_utils.v(44)
  not \C023/C01/u1  (\C023/outtemp [2], temp_exp_diff[2]);  // ../RTL/core/fpu_utils.v(44)
  not \C023/C01/u2  (\C023/outtemp [1], temp_exp_diff[1]);  // ../RTL/core/fpu_utils.v(44)
  not \C023/C01/u4  (\C023/outtemp [7], temp_exp_diff[7]);  // ../RTL/core/fpu_utils.v(44)
  not \C023/C01/u5  (\C023/outtemp [6], temp_exp_diff[6]);  // ../RTL/core/fpu_utils.v(44)
  not \C023/C01/u6  (\C023/outtemp [5], temp_exp_diff[5]);  // ../RTL/core/fpu_utils.v(44)
  not \C023/C01/u7  (\C023/outtemp [4], temp_exp_diff[4]);  // ../RTL/core/fpu_utils.v(44)
  and \C03/ADD01/ADD01/ADD01/u10  (\C03/ADD01/ADD01/ADD01/n1 , \C03/outtemp [1], \C03/outtemp [0]);  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD01/ADD01/u17  (\C03/ADD01/ADD01/ADD01/n7 , \C03/outtemp [2], \C03/outtemp [1]);  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD01/ADD01/u18  (\C03/ADD01/ADD01/ADD01/n8 , \C03/ADD01/ADD01/ADD01/n7 , \C03/outtemp [0]);  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD01/ADD01/u20  (complemented_M_result[3], \C03/outtemp [3], \C03/ADD01/ADD01/ADD01/n8 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD01/ADD01/u26  (\C03/ADD01/ADD01/ADD01/n14 , \C03/outtemp [3], \C03/outtemp [2]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD01/ADD01/u29  (complemented_M_result[2], \C03/outtemp [2], \C03/ADD01/ADD01/ADD01/n1 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD01/ADD01/u30  (\C03/ADD01/ADD01/ADD01/n17 , \C03/ADD01/ADD01/ADD01/n14 , \C03/outtemp [1]);  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD01/ADD01/u31  (\C03/ADD01/ADD01/ADD01/n18 , \C03/ADD01/ADD01/ADD01/n17 , \C03/outtemp [0]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD01/ADD01/u33  (complemented_M_result[1], \C03/outtemp [1], \C03/outtemp [0]);  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD01/ADD02/u12  (\C03/ADD01/ADD01/ADD02/n3 , \C03/outtemp [5], \C03/outtemp [4]);  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD01/ADD02/u13  (\C03/ADD01/ADD01/ADD02/n4 , \C03/ADD01/ADD01/ADD02/n3 , \C03/ADD01/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD01/ADD02/u17  (\C03/ADD01/ADD01/ADD02/n7 , \C03/outtemp [6], \C03/outtemp [5]);  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD01/ADD02/u20  (complemented_M_result[7], \C03/outtemp [7], \C03/ADD01/ADD01/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD01/ADD02/u21  (\C03/ADD01/ADD01/ADD02/n10 , \C03/ADD01/ADD01/ADD02/n7 , \C03/outtemp [4]);  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD01/ADD02/u22  (\C03/ADD01/ADD01/ADD02/n11 , \C03/ADD01/ADD01/ADD02/n10 , \C03/ADD01/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD01/ADD02/u26  (\C03/ADD01/ADD01/ADD02/n14 , \C03/outtemp [7], \C03/outtemp [6]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD01/ADD02/u29  (complemented_M_result[6], \C03/outtemp [6], \C03/ADD01/ADD01/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD01/ADD02/u30  (\C03/ADD01/ADD01/ADD02/n17 , \C03/ADD01/ADD01/ADD02/n14 , \C03/outtemp [5]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD01/ADD02/u33  (complemented_M_result[5], \C03/outtemp [5], \C03/ADD01/ADD01/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \C03/ADD01/ADD01/ADD02/u34  (complemented_M_result[4], \C03/outtemp [4], \C03/ADD01/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD01/ADD02/u35  (\C03/ADD01/ADD01/ADD02/n20 , \C03/ADD01/ADD01/ADD02/n17 , \C03/outtemp [4]);  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD01/ADD02/u36  (\C03/ADD01/ADD01/ADD02/n21 , \C03/ADD01/ADD01/ADD02/n20 , \C03/ADD01/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD01/ADD02/u8  (\C03/ADD01/ADD01/ADD02/n0 , \C03/outtemp [4], \C03/ADD01/ADD01/ADD01/n18 );  // ../RTL/core/fpu_utils.v(63)
  and \C03/ADD01/ADD02/ADD01/u12  (\C03/ADD01/ADD02/ADD01/n3 , \C03/outtemp [9], \C03/outtemp [8]);  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD02/ADD01/u13  (\C03/ADD01/ADD02/ADD01/n4 , \C03/ADD01/ADD02/ADD01/n3 , \C03/ADD01/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD02/ADD01/u17  (\C03/ADD01/ADD02/ADD01/n7 , \C03/outtemp [10], \C03/outtemp [9]);  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD02/ADD01/u20  (complemented_M_result[11], \C03/outtemp [11], \C03/ADD01/ADD02/ADD01/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD02/ADD01/u21  (\C03/ADD01/ADD02/ADD01/n10 , \C03/ADD01/ADD02/ADD01/n7 , \C03/outtemp [8]);  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD02/ADD01/u22  (\C03/ADD01/ADD02/ADD01/n11 , \C03/ADD01/ADD02/ADD01/n10 , \C03/ADD01/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD02/ADD01/u26  (\C03/ADD01/ADD02/ADD01/n14 , \C03/outtemp [11], \C03/outtemp [10]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD02/ADD01/u29  (complemented_M_result[10], \C03/outtemp [10], \C03/ADD01/ADD02/ADD01/n4 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD02/ADD01/u30  (\C03/ADD01/ADD02/ADD01/n17 , \C03/ADD01/ADD02/ADD01/n14 , \C03/outtemp [9]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD02/ADD01/u33  (complemented_M_result[9], \C03/outtemp [9], \C03/ADD01/ADD02/ADD01/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \C03/ADD01/ADD02/ADD01/u34  (complemented_M_result[8], \C03/outtemp [8], \C03/ADD01/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD02/ADD01/u35  (\C03/ADD01/ADD02/ADD01/n20 , \C03/ADD01/ADD02/ADD01/n17 , \C03/outtemp [8]);  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD02/ADD01/u36  (\C03/ADD01/ADD02/ADD01/n21 , \C03/ADD01/ADD02/ADD01/n20 , \C03/ADD01/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD02/ADD01/u8  (\C03/ADD01/ADD02/ADD01/n0 , \C03/outtemp [8], \C03/ADD01/ADD01/ADD02/n21 );  // ../RTL/core/fpu_utils.v(63)
  and \C03/ADD01/ADD02/ADD02/u12  (\C03/ADD01/ADD02/ADD02/n3 , \C03/outtemp [13], \C03/outtemp [12]);  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD02/ADD02/u13  (\C03/ADD01/ADD02/ADD02/n4 , \C03/ADD01/ADD02/ADD02/n3 , \C03/ADD01/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD02/ADD02/u17  (\C03/ADD01/ADD02/ADD02/n7 , \C03/outtemp [14], \C03/outtemp [13]);  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD02/ADD02/u20  (complemented_M_result[15], \C03/outtemp [15], \C03/ADD01/ADD02/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD02/ADD02/u21  (\C03/ADD01/ADD02/ADD02/n10 , \C03/ADD01/ADD02/ADD02/n7 , \C03/outtemp [12]);  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD02/ADD02/u22  (\C03/ADD01/ADD02/ADD02/n11 , \C03/ADD01/ADD02/ADD02/n10 , \C03/ADD01/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD02/ADD02/u26  (\C03/ADD01/ADD02/ADD02/n14 , \C03/outtemp [15], \C03/outtemp [14]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD02/ADD02/u29  (complemented_M_result[14], \C03/outtemp [14], \C03/ADD01/ADD02/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD02/ADD02/u30  (\C03/ADD01/ADD02/ADD02/n17 , \C03/ADD01/ADD02/ADD02/n14 , \C03/outtemp [13]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD02/ADD02/u33  (complemented_M_result[13], \C03/outtemp [13], \C03/ADD01/ADD02/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \C03/ADD01/ADD02/ADD02/u34  (complemented_M_result[12], \C03/outtemp [12], \C03/ADD01/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD02/ADD02/u35  (\C03/ADD01/ADD02/ADD02/n20 , \C03/ADD01/ADD02/ADD02/n17 , \C03/outtemp [12]);  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD02/ADD02/u36  (\C03/ADD01/ADD02/ADD02/n21 , \C03/ADD01/ADD02/ADD02/n20 , \C03/ADD01/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD02/ADD02/u8  (\C03/ADD01/ADD02/ADD02/n0 , \C03/outtemp [12], \C03/ADD01/ADD02/ADD01/n21 );  // ../RTL/core/fpu_utils.v(63)
  and \C03/ADD01/ADD03/ADD01/u12  (\C03/ADD01/ADD03/ADD01/n3 , \C03/outtemp [17], \C03/outtemp [16]);  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD03/ADD01/u13  (\C03/ADD01/ADD03/ADD01/n4 , \C03/ADD01/ADD03/ADD01/n3 , \C03/ADD01/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD03/ADD01/u17  (\C03/ADD01/ADD03/ADD01/n7 , \C03/outtemp [18], \C03/outtemp [17]);  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD03/ADD01/u20  (complemented_M_result[19], \C03/outtemp [19], \C03/ADD01/ADD03/ADD01/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD03/ADD01/u21  (\C03/ADD01/ADD03/ADD01/n10 , \C03/ADD01/ADD03/ADD01/n7 , \C03/outtemp [16]);  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD03/ADD01/u22  (\C03/ADD01/ADD03/ADD01/n11 , \C03/ADD01/ADD03/ADD01/n10 , \C03/ADD01/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD03/ADD01/u26  (\C03/ADD01/ADD03/ADD01/n14 , \C03/outtemp [19], \C03/outtemp [18]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD03/ADD01/u29  (complemented_M_result[18], \C03/outtemp [18], \C03/ADD01/ADD03/ADD01/n4 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD03/ADD01/u30  (\C03/ADD01/ADD03/ADD01/n17 , \C03/ADD01/ADD03/ADD01/n14 , \C03/outtemp [17]);  // ../RTL/core/fpu_utils.v(66)
  xor \C03/ADD01/ADD03/ADD01/u33  (complemented_M_result[17], \C03/outtemp [17], \C03/ADD01/ADD03/ADD01/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \C03/ADD01/ADD03/ADD01/u34  (complemented_M_result[16], \C03/outtemp [16], \C03/ADD01/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD03/ADD01/u35  (\C03/ADD01/ADD03/ADD01/n20 , \C03/ADD01/ADD03/ADD01/n17 , \C03/outtemp [16]);  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD03/ADD01/u36  (\C03/ADD01/ADD03/ADD01/n21 , \C03/ADD01/ADD03/ADD01/n20 , \C03/ADD01/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(66)
  and \C03/ADD01/ADD03/ADD01/u8  (\C03/ADD01/ADD03/ADD01/n0 , \C03/outtemp [16], \C03/ADD01/ADD02/ADD02/n21 );  // ../RTL/core/fpu_utils.v(63)
  and \C03/ADD01/ADD03/ADD02/u12  (\C03/ADD01/ADD03/ADD02/n3 , \C03/outtemp [21], \C03/outtemp [20]);  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD03/ADD02/u13  (\C03/ADD01/ADD03/ADD02/n4 , \C03/ADD01/ADD03/ADD02/n3 , \C03/ADD01/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(64)
  and \C03/ADD01/ADD03/ADD02/u17  (\C03/ADD01/ADD03/ADD02/n7 , \C03/outtemp [22], \C03/outtemp [21]);  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD03/ADD02/u20  (complemented_M_result[23], \C03/outtemp [23], \C03/ADD01/ADD03/ADD02/n11 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD03/ADD02/u21  (\C03/ADD01/ADD03/ADD02/n10 , \C03/ADD01/ADD03/ADD02/n7 , \C03/outtemp [20]);  // ../RTL/core/fpu_utils.v(65)
  and \C03/ADD01/ADD03/ADD02/u22  (\C03/ADD01/ADD03/ADD02/n11 , \C03/ADD01/ADD03/ADD02/n10 , \C03/ADD01/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(65)
  xor \C03/ADD01/ADD03/ADD02/u29  (complemented_M_result[22], \C03/outtemp [22], \C03/ADD01/ADD03/ADD02/n4 );  // ../RTL/core/fpu_utils.v(71)
  xor \C03/ADD01/ADD03/ADD02/u33  (complemented_M_result[21], \C03/outtemp [21], \C03/ADD01/ADD03/ADD02/n0 );  // ../RTL/core/fpu_utils.v(71)
  xor \C03/ADD01/ADD03/ADD02/u34  (complemented_M_result[20], \C03/outtemp [20], \C03/ADD01/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(71)
  and \C03/ADD01/ADD03/ADD02/u8  (\C03/ADD01/ADD03/ADD02/n0 , \C03/outtemp [20], \C03/ADD01/ADD03/ADD01/n21 );  // ../RTL/core/fpu_utils.v(63)
  not \C03/C01/C01/u0  (\C03/outtemp [3], M_result[3]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u1  (\C03/outtemp [2], M_result[2]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u2  (\C03/outtemp [1], M_result[1]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u3  (\C03/outtemp [0], M_result[0]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u4  (\C03/outtemp [7], M_result[7]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u5  (\C03/outtemp [6], M_result[6]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u6  (\C03/outtemp [5], M_result[5]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C01/u7  (\C03/outtemp [4], M_result[4]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u0  (\C03/outtemp [11], M_result[11]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u1  (\C03/outtemp [10], M_result[10]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u2  (\C03/outtemp [9], M_result[9]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u3  (\C03/outtemp [8], M_result[8]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u4  (\C03/outtemp [15], M_result[15]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u5  (\C03/outtemp [14], M_result[14]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u6  (\C03/outtemp [13], M_result[13]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C02/u7  (\C03/outtemp [12], M_result[12]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u0  (\C03/outtemp [19], M_result[19]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u1  (\C03/outtemp [18], M_result[18]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u2  (\C03/outtemp [17], M_result[17]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u3  (\C03/outtemp [16], M_result[16]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u4  (\C03/outtemp [23], M_result[23]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u5  (\C03/outtemp [22], M_result[22]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u6  (\C03/outtemp [21], M_result[21]);  // ../RTL/core/fpu_utils.v(44)
  not \C03/C01/C03/u7  (\C03/outtemp [20], M_result[20]);  // ../RTL/core/fpu_utils.v(44)
  not \C04/u0  (complemented_shift_E[3], shift_E[3]);  // ../RTL/core/fpu_utils.v(44)
  not \C04/u1  (complemented_shift_E[2], shift_E[2]);  // ../RTL/core/fpu_utils.v(44)
  not \C04/u2  (complemented_shift_E[1], shift_E[1]);  // ../RTL/core/fpu_utils.v(44)
  not \C04/u3  (complemented_shift_E[0], shift_E[0]);  // ../RTL/core/fpu_utils.v(44)
  not \C04/u7  (complemented_shift_E[4], shift_E[4]);  // ../RTL/core/fpu_utils.v(44)
  AL_MUX \M011/M02/u3  (
    .i0(complemented_temp_exp_diff[1]),
    .i1(temp_exp_diff[1]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[1]));
  AL_MUX \M011/M03/u3  (
    .i0(complemented_temp_exp_diff[2]),
    .i1(temp_exp_diff[2]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[2]));
  AL_MUX \M011/M04/u3  (
    .i0(complemented_temp_exp_diff[3]),
    .i1(temp_exp_diff[3]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[3]));
  AL_MUX \M011/M05/u3  (
    .i0(complemented_temp_exp_diff[4]),
    .i1(temp_exp_diff[4]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[4]));
  AL_MUX \M011/M06/u3  (
    .i0(complemented_temp_exp_diff[5]),
    .i1(temp_exp_diff[5]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[5]));
  AL_MUX \M011/M07/u3  (
    .i0(complemented_temp_exp_diff[6]),
    .i1(temp_exp_diff[6]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[6]));
  AL_MUX \M011/M08/u3  (
    .i0(complemented_temp_exp_diff[7]),
    .i1(temp_exp_diff[7]),
    .sel(isE1GreaterThanE2),
    .o(exp_diff[7]));
  AL_MUX \M03/M01/u3  (
    .i0(n2[23]),
    .i1(n1[23]),
    .sel(isE1GreaterThanE2),
    .o(E[0]));
  AL_MUX \M03/M02/u3  (
    .i0(n2[24]),
    .i1(n1[24]),
    .sel(isE1GreaterThanE2),
    .o(E[1]));
  AL_MUX \M03/M03/u3  (
    .i0(n2[25]),
    .i1(n1[25]),
    .sel(isE1GreaterThanE2),
    .o(E[2]));
  AL_MUX \M03/M04/u3  (
    .i0(n2[26]),
    .i1(n1[26]),
    .sel(isE1GreaterThanE2),
    .o(E[3]));
  AL_MUX \M03/M05/u3  (
    .i0(n2[27]),
    .i1(n1[27]),
    .sel(isE1GreaterThanE2),
    .o(E[4]));
  AL_MUX \M03/M06/u3  (
    .i0(n2[28]),
    .i1(n1[28]),
    .sel(isE1GreaterThanE2),
    .o(E[5]));
  AL_MUX \M03/M07/u3  (
    .i0(n2[29]),
    .i1(n1[29]),
    .sel(isE1GreaterThanE2),
    .o(E[6]));
  AL_MUX \M03/M08/u3  (
    .i0(n2[30]),
    .i1(n1[30]),
    .sel(isE1GreaterThanE2),
    .o(E[7]));
  not \M031/M01/u0  (\M031/M01/invSL , \NM/n2 );  // ../RTL/core/fpu_utils.v(106)
  AL_MUX \M031/M01/u3  (
    .i0(\NM/n2 ),
    .i1(\M031/M01/invSL ),
    .sel(E[0]),
    .o(new_E[0]));
  AL_MUX \M031/M02/u3  (
    .i0(E[1]),
    .i1(One_Added_E[1]),
    .sel(\NM/n2 ),
    .o(new_E[1]));
  AL_MUX \M031/M03/u3  (
    .i0(E[2]),
    .i1(One_Added_E[2]),
    .sel(\NM/n2 ),
    .o(new_E[2]));
  AL_MUX \M031/M04/u3  (
    .i0(E[3]),
    .i1(One_Added_E[3]),
    .sel(\NM/n2 ),
    .o(new_E[3]));
  AL_MUX \M031/M05/u3  (
    .i0(E[4]),
    .i1(One_Added_E[4]),
    .sel(\NM/n2 ),
    .o(new_E[4]));
  AL_MUX \M031/M06/u3  (
    .i0(E[5]),
    .i1(One_Added_E[5]),
    .sel(\NM/n2 ),
    .o(new_E[5]));
  AL_MUX \M031/M07/u3  (
    .i0(E[6]),
    .i1(One_Added_E[6]),
    .sel(\NM/n2 ),
    .o(new_E[6]));
  AL_MUX \M031/M08/u3  (
    .i0(E[7]),
    .i1(One_Added_E[7]),
    .sel(\NM/n2 ),
    .o(new_E[7]));
  not \M04/M01/M01/u0  (\M04/M01/M01/invSL , real_oper);  // ../RTL/core/fpu_utils.v(106)
  AL_MUX \M04/M01/M01/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[0]),
    .o(new_M2[0]));
  AL_MUX \M04/M01/M02/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[1]),
    .o(new_M2[1]));
  AL_MUX \M04/M01/M03/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[2]),
    .o(new_M2[2]));
  AL_MUX \M04/M01/M04/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[3]),
    .o(new_M2[3]));
  AL_MUX \M04/M01/M05/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[4]),
    .o(new_M2[4]));
  AL_MUX \M04/M01/M06/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[5]),
    .o(new_M2[5]));
  AL_MUX \M04/M01/M07/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[6]),
    .o(new_M2[6]));
  AL_MUX \M04/M01/M08/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[7]),
    .o(new_M2[7]));
  AL_MUX \M04/M02/M01/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[8]),
    .o(new_M2[8]));
  AL_MUX \M04/M02/M02/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[9]),
    .o(new_M2[9]));
  AL_MUX \M04/M02/M03/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[10]),
    .o(new_M2[10]));
  AL_MUX \M04/M02/M04/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[11]),
    .o(new_M2[11]));
  AL_MUX \M04/M02/M05/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[12]),
    .o(new_M2[12]));
  AL_MUX \M04/M02/M06/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[13]),
    .o(new_M2[13]));
  AL_MUX \M04/M02/M07/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[14]),
    .o(new_M2[14]));
  AL_MUX \M04/M02/M08/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[15]),
    .o(new_M2[15]));
  AL_MUX \M04/M03/M01/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[16]),
    .o(new_M2[16]));
  AL_MUX \M04/M03/M02/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[17]),
    .o(new_M2[17]));
  AL_MUX \M04/M03/M03/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[18]),
    .o(new_M2[18]));
  AL_MUX \M04/M03/M04/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[19]),
    .o(new_M2[19]));
  AL_MUX \M04/M03/M05/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[20]),
    .o(new_M2[20]));
  AL_MUX \M04/M03/M06/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[21]),
    .o(new_M2[21]));
  AL_MUX \M04/M03/M07/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[22]),
    .o(new_M2[22]));
  AL_MUX \M04/M03/M08/u3  (
    .i0(real_oper),
    .i1(\M04/M01/M01/invSL ),
    .sel(M2[23]),
    .o(new_M2[23]));
  AL_MUX \M05/M01/M02/u3  (
    .i0(M_result[1]),
    .i1(complemented_M_result[1]),
    .sel(n196),
    .o(M_result2[1]));
  AL_MUX \M05/M01/M03/u3  (
    .i0(M_result[2]),
    .i1(complemented_M_result[2]),
    .sel(n196),
    .o(M_result2[2]));
  AL_MUX \M05/M01/M04/u3  (
    .i0(M_result[3]),
    .i1(complemented_M_result[3]),
    .sel(n196),
    .o(M_result2[3]));
  AL_MUX \M05/M01/M05/u3  (
    .i0(M_result[4]),
    .i1(complemented_M_result[4]),
    .sel(n196),
    .o(M_result2[4]));
  AL_MUX \M05/M01/M06/u3  (
    .i0(M_result[5]),
    .i1(complemented_M_result[5]),
    .sel(n196),
    .o(M_result2[5]));
  AL_MUX \M05/M01/M07/u3  (
    .i0(M_result[6]),
    .i1(complemented_M_result[6]),
    .sel(n196),
    .o(M_result2[6]));
  AL_MUX \M05/M01/M08/u3  (
    .i0(M_result[7]),
    .i1(complemented_M_result[7]),
    .sel(n196),
    .o(M_result2[7]));
  AL_MUX \M05/M02/M01/u3  (
    .i0(M_result[8]),
    .i1(complemented_M_result[8]),
    .sel(n196),
    .o(M_result2[8]));
  AL_MUX \M05/M02/M02/u3  (
    .i0(M_result[9]),
    .i1(complemented_M_result[9]),
    .sel(n196),
    .o(M_result2[9]));
  AL_MUX \M05/M02/M03/u3  (
    .i0(M_result[10]),
    .i1(complemented_M_result[10]),
    .sel(n196),
    .o(M_result2[10]));
  AL_MUX \M05/M02/M04/u3  (
    .i0(M_result[11]),
    .i1(complemented_M_result[11]),
    .sel(n196),
    .o(M_result2[11]));
  AL_MUX \M05/M02/M05/u3  (
    .i0(M_result[12]),
    .i1(complemented_M_result[12]),
    .sel(n196),
    .o(M_result2[12]));
  AL_MUX \M05/M02/M06/u3  (
    .i0(M_result[13]),
    .i1(complemented_M_result[13]),
    .sel(n196),
    .o(M_result2[13]));
  AL_MUX \M05/M02/M07/u3  (
    .i0(M_result[14]),
    .i1(complemented_M_result[14]),
    .sel(n196),
    .o(M_result2[14]));
  AL_MUX \M05/M02/M08/u3  (
    .i0(M_result[15]),
    .i1(complemented_M_result[15]),
    .sel(n196),
    .o(M_result2[15]));
  AL_MUX \M05/M03/M01/u3  (
    .i0(M_result[16]),
    .i1(complemented_M_result[16]),
    .sel(n196),
    .o(M_result2[16]));
  AL_MUX \M05/M03/M02/u3  (
    .i0(M_result[17]),
    .i1(complemented_M_result[17]),
    .sel(n196),
    .o(M_result2[17]));
  AL_MUX \M05/M03/M03/u3  (
    .i0(M_result[18]),
    .i1(complemented_M_result[18]),
    .sel(n196),
    .o(M_result2[18]));
  AL_MUX \M05/M03/M04/u3  (
    .i0(M_result[19]),
    .i1(complemented_M_result[19]),
    .sel(n196),
    .o(M_result2[19]));
  AL_MUX \M05/M03/M05/u3  (
    .i0(M_result[20]),
    .i1(complemented_M_result[20]),
    .sel(n196),
    .o(M_result2[20]));
  AL_MUX \M05/M03/M06/u3  (
    .i0(M_result[21]),
    .i1(complemented_M_result[21]),
    .sel(n196),
    .o(M_result2[21]));
  AL_MUX \M05/M03/M07/u3  (
    .i0(M_result[22]),
    .i1(complemented_M_result[22]),
    .sel(n196),
    .o(M_result2[22]));
  AL_MUX \M05/M03/M08/u3  (
    .i0(M_result[23]),
    .i1(complemented_M_result[23]),
    .sel(n196),
    .o(M_result2[23]));
  add_pu23_pu23_o23 \NM/add0  (
    .i0(M_result2[23:1]),
    .i1({22'b0000000000000000000000,M_result[0]}),
    .o(\NM/n4 ));  // ../RTL/core/fpu_utils.v(158)
  eq_w24 \NM/eq0  (
    .i0({M_result2[23:1],M_result[0]}),
    .i1(24'b000000000000000000000001),
    .o(\NM/n51 ));  // ../RTL/core/fpu_utils.v(301)
  binary_mux_s1_w1 \NM/mux0_b0  (
    .i0(\NM/n122 [0]),
    .i1(\NM/n4 [0]),
    .sel(\NM/n2 ),
    .o(result[0]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b1  (
    .i0(\NM/sel0_b1/or_B23_B24_o ),
    .i1(\NM/n4 [1]),
    .sel(\NM/n2 ),
    .o(result[1]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b10  (
    .i0(\NM/sel0_b10/or_or_or_B12_or_B13__o ),
    .i1(\NM/n4 [10]),
    .sel(\NM/n2 ),
    .o(result[10]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b11  (
    .i0(\NM/sel0_b11/or_or_or_B12_or_B13__o ),
    .i1(\NM/n4 [11]),
    .sel(\NM/n2 ),
    .o(result[11]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b12  (
    .i0(\NM/sel0_b12/or_or_or_B12_or_B13__o ),
    .i1(\NM/n4 [12]),
    .sel(\NM/n2 ),
    .o(result[12]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b13  (
    .i0(\NM/n122 [13]),
    .i1(\NM/n4 [13]),
    .sel(\NM/n2 ),
    .o(result[13]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b14  (
    .i0(\NM/n122 [14]),
    .i1(\NM/n4 [14]),
    .sel(\NM/n2 ),
    .o(result[14]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b15  (
    .i0(\NM/n122 [15]),
    .i1(\NM/n4 [15]),
    .sel(\NM/n2 ),
    .o(result[15]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b16  (
    .i0(\NM/n122 [16]),
    .i1(\NM/n4 [16]),
    .sel(\NM/n2 ),
    .o(result[16]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b17  (
    .i0(\NM/n122 [17]),
    .i1(\NM/n4 [17]),
    .sel(\NM/n2 ),
    .o(result[17]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b18  (
    .i0(\NM/n122 [18]),
    .i1(\NM/n4 [18]),
    .sel(\NM/n2 ),
    .o(result[18]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b19  (
    .i0(\NM/n122 [19]),
    .i1(\NM/n4 [19]),
    .sel(\NM/n2 ),
    .o(result[19]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b2  (
    .i0(\NM/sel0_b2/or_or_B21_B22_o_or_B_o ),
    .i1(\NM/n4 [2]),
    .sel(\NM/n2 ),
    .o(result[2]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b20  (
    .i0(\NM/n122 [20]),
    .i1(\NM/n4 [20]),
    .sel(\NM/n2 ),
    .o(result[20]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b21  (
    .i0(\NM/n122 [21]),
    .i1(\NM/n4 [21]),
    .sel(\NM/n2 ),
    .o(result[21]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b22  (
    .i0(\NM/n122 [22]),
    .i1(\NM/n4 [22]),
    .sel(\NM/n2 ),
    .o(result[22]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b3  (
    .i0(\NM/sel0_b3/or_or_B21_B22_o_or_B_o ),
    .i1(\NM/n4 [3]),
    .sel(\NM/n2 ),
    .o(result[3]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b4  (
    .i0(\NM/sel0_b4/or_or_B18_or_B19_B20_o ),
    .i1(\NM/n4 [4]),
    .sel(\NM/n2 ),
    .o(result[4]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b5  (
    .i0(\NM/sel0_b5/or_or_B18_or_B19_B20_o ),
    .i1(\NM/n4 [5]),
    .sel(\NM/n2 ),
    .o(result[5]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b6  (
    .i0(\NM/sel0_b6/or_or_B18_or_B19_B20_o ),
    .i1(\NM/n4 [6]),
    .sel(\NM/n2 ),
    .o(result[6]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b7  (
    .i0(\NM/sel0_b7/or_or_or_B12_or_B13__o ),
    .i1(\NM/n4 [7]),
    .sel(\NM/n2 ),
    .o(result[7]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b8  (
    .i0(\NM/sel0_b8/or_or_or_B12_or_B13__o ),
    .i1(\NM/n4 [8]),
    .sel(\NM/n2 ),
    .o(result[8]));  // ../RTL/core/fpu_utils.v(156)
  binary_mux_s1_w1 \NM/mux0_b9  (
    .i0(\NM/sel0_b9/or_or_or_B12_or_B13__o ),
    .i1(\NM/n4 [9]),
    .sel(\NM/n2 ),
    .o(result[9]));  // ../RTL/core/fpu_utils.v(156)
  AL_MUX \NM/mux1_b0  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\NM/mux1_b0_sel_is_2_o ),
    .o(shift_E[0]));
  and \NM/mux1_b0_sel_is_2  (\NM/mux1_b0_sel_is_2_o , \M031/M01/invSL , \NM/sel1_b0_sel_o );
  AL_MUX \NM/mux1_b1  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\NM/mux1_b1_sel_is_2_o ),
    .o(shift_E[1]));
  and \NM/mux1_b1_sel_is_2  (\NM/mux1_b1_sel_is_2_o , \M031/M01/invSL , \NM/sel1_b1_sel_o );
  AL_MUX \NM/mux1_b2  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\NM/mux1_b2_sel_is_2_o ),
    .o(shift_E[2]));
  and \NM/mux1_b2_sel_is_2  (\NM/mux1_b2_sel_is_2_o , \M031/M01/invSL , \NM/sel1_b2_sel_o );
  AL_MUX \NM/mux1_b3  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\NM/mux1_b3_sel_is_2_o ),
    .o(shift_E[3]));
  and \NM/mux1_b3_sel_is_2  (\NM/mux1_b3_sel_is_2_o , \M031/M01/invSL , \NM/sel1_b3_sel_o );
  AL_MUX \NM/mux1_b4  (
    .i0(1'b0),
    .i1(1'b1),
    .sel(\NM/mux1_b4_sel_is_2_o ),
    .o(shift_E[4]));
  and \NM/mux1_b4_sel_is_2  (\NM/mux1_b4_sel_is_2_o , \M031/M01/invSL , \NM/sel1_b4_sel_o );
  AL_MUX \NM/sel0_b0  (
    .i0(1'b0),
    .i1(M_result[0]),
    .sel(M_result2[23]),
    .o(\NM/n122 [0]));  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b1/and_b0_23  (\NM/sel0_b1/B23 , M_result[0], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b1/and_b0_24  (\NM/sel0_b1/B24 , M_result2[1], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b1/or_B23_B24  (\NM/sel0_b1/or_B23_B24_o , \NM/sel0_b1/B23 , \NM/sel0_b1/B24 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_14  (\NM/sel0_b10/B14 , M_result[0], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_15  (\NM/sel0_b10/B15 , M_result2[1], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_16  (\NM/sel0_b10/B16 , M_result2[2], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_17  (\NM/sel0_b10/B17 , M_result2[3], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_18  (\NM/sel0_b10/B18 , M_result2[4], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_19  (\NM/sel0_b10/B19 , M_result2[5], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_20  (\NM/sel0_b10/B20 , M_result2[6], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_21  (\NM/sel0_b10/B21 , M_result2[7], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_22  (\NM/sel0_b10/B22 , M_result2[8], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_23  (\NM/sel0_b10/B23 , M_result2[9], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b10/and_b0_24  (\NM/sel0_b10/B24 , M_result2[10], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_B15_or_B16_B17_o  (\NM/sel0_b10/or_B15_or_B16_B17_o_o , \NM/sel0_b10/B15 , \NM/sel0_b10/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_B16_B17  (\NM/sel0_b10/or_B16_B17_o , \NM/sel0_b10/B16 , \NM/sel0_b10/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_B18_or_B19_B20_o  (\NM/sel0_b10/or_B18_or_B19_B20_o_o , \NM/sel0_b10/B18 , \NM/sel0_b10/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_B19_B20  (\NM/sel0_b10/or_B19_B20_o , \NM/sel0_b10/B19 , \NM/sel0_b10/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_B21_B22  (\NM/sel0_b10/or_B21_B22_o , \NM/sel0_b10/B21 , \NM/sel0_b10/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_B23_B24  (\NM/sel0_b10/or_B23_B24_o , \NM/sel0_b10/B23 , \NM/sel0_b10/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_or_B12_or_B13_B14  (\NM/sel0_b10/or_or_B12_or_B13_B14_o , \NM/sel0_b10/B14 , \NM/sel0_b10/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_or_B18_or_B19_B20  (\NM/sel0_b10/or_or_B18_or_B19_B20_o , \NM/sel0_b10/or_B18_or_B19_B20_o_o , \NM/sel0_b10/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_or_B21_B22_o_or_B  (\NM/sel0_b10/or_or_B21_B22_o_or_B_o , \NM/sel0_b10/or_B21_B22_o , \NM/sel0_b10/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b10/or_or_or_B12_or_B13_  (\NM/sel0_b10/or_or_or_B12_or_B13__o , \NM/sel0_b10/or_or_B12_or_B13_B14_o , \NM/sel0_b10/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_13  (\NM/sel0_b11/B13 , M_result[0], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_14  (\NM/sel0_b11/B14 , M_result2[1], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_15  (\NM/sel0_b11/B15 , M_result2[2], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_16  (\NM/sel0_b11/B16 , M_result2[3], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_17  (\NM/sel0_b11/B17 , M_result2[4], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_18  (\NM/sel0_b11/B18 , M_result2[5], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_19  (\NM/sel0_b11/B19 , M_result2[6], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_20  (\NM/sel0_b11/B20 , M_result2[7], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_21  (\NM/sel0_b11/B21 , M_result2[8], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_22  (\NM/sel0_b11/B22 , M_result2[9], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_23  (\NM/sel0_b11/B23 , M_result2[10], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b11/and_b0_24  (\NM/sel0_b11/B24 , M_result2[11], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B13_B14  (\NM/sel0_b11/or_B13_B14_o , \NM/sel0_b11/B13 , \NM/sel0_b11/B14 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B15_or_B16_B17_o  (\NM/sel0_b11/or_B15_or_B16_B17_o_o , \NM/sel0_b11/B15 , \NM/sel0_b11/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B16_B17  (\NM/sel0_b11/or_B16_B17_o , \NM/sel0_b11/B16 , \NM/sel0_b11/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B18_or_B19_B20_o  (\NM/sel0_b11/or_B18_or_B19_B20_o_o , \NM/sel0_b11/B18 , \NM/sel0_b11/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B19_B20  (\NM/sel0_b11/or_B19_B20_o , \NM/sel0_b11/B19 , \NM/sel0_b11/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B21_B22  (\NM/sel0_b11/or_B21_B22_o , \NM/sel0_b11/B21 , \NM/sel0_b11/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_B23_B24  (\NM/sel0_b11/or_B23_B24_o , \NM/sel0_b11/B23 , \NM/sel0_b11/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_or_B12_or_B13_B14  (\NM/sel0_b11/or_or_B12_or_B13_B14_o , \NM/sel0_b11/or_B13_B14_o , \NM/sel0_b11/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_or_B18_or_B19_B20  (\NM/sel0_b11/or_or_B18_or_B19_B20_o , \NM/sel0_b11/or_B18_or_B19_B20_o_o , \NM/sel0_b11/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_or_B21_B22_o_or_B  (\NM/sel0_b11/or_or_B21_B22_o_or_B_o , \NM/sel0_b11/or_B21_B22_o , \NM/sel0_b11/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b11/or_or_or_B12_or_B13_  (\NM/sel0_b11/or_or_or_B12_or_B13__o , \NM/sel0_b11/or_or_B12_or_B13_B14_o , \NM/sel0_b11/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_12  (\NM/sel0_b12/B12 , M_result[0], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_13  (\NM/sel0_b12/B13 , M_result2[1], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_14  (\NM/sel0_b12/B14 , M_result2[2], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_15  (\NM/sel0_b12/B15 , M_result2[3], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_16  (\NM/sel0_b12/B16 , M_result2[4], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_17  (\NM/sel0_b12/B17 , M_result2[5], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_18  (\NM/sel0_b12/B18 , M_result2[6], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_19  (\NM/sel0_b12/B19 , M_result2[7], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_20  (\NM/sel0_b12/B20 , M_result2[8], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_21  (\NM/sel0_b12/B21 , M_result2[9], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_22  (\NM/sel0_b12/B22 , M_result2[10], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_23  (\NM/sel0_b12/B23 , M_result2[11], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b12/and_b0_24  (\NM/sel0_b12/B24 , M_result2[12], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B12_or_B13_B14_o  (\NM/sel0_b12/or_B12_or_B13_B14_o_o , \NM/sel0_b12/B12 , \NM/sel0_b12/or_B13_B14_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B13_B14  (\NM/sel0_b12/or_B13_B14_o , \NM/sel0_b12/B13 , \NM/sel0_b12/B14 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B15_or_B16_B17_o  (\NM/sel0_b12/or_B15_or_B16_B17_o_o , \NM/sel0_b12/B15 , \NM/sel0_b12/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B16_B17  (\NM/sel0_b12/or_B16_B17_o , \NM/sel0_b12/B16 , \NM/sel0_b12/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B18_or_B19_B20_o  (\NM/sel0_b12/or_B18_or_B19_B20_o_o , \NM/sel0_b12/B18 , \NM/sel0_b12/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B19_B20  (\NM/sel0_b12/or_B19_B20_o , \NM/sel0_b12/B19 , \NM/sel0_b12/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B21_B22  (\NM/sel0_b12/or_B21_B22_o , \NM/sel0_b12/B21 , \NM/sel0_b12/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_B23_B24  (\NM/sel0_b12/or_B23_B24_o , \NM/sel0_b12/B23 , \NM/sel0_b12/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_or_B12_or_B13_B14  (\NM/sel0_b12/or_or_B12_or_B13_B14_o , \NM/sel0_b12/or_B12_or_B13_B14_o_o , \NM/sel0_b12/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_or_B18_or_B19_B20  (\NM/sel0_b12/or_or_B18_or_B19_B20_o , \NM/sel0_b12/or_B18_or_B19_B20_o_o , \NM/sel0_b12/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_or_B21_B22_o_or_B  (\NM/sel0_b12/or_or_B21_B22_o_or_B_o , \NM/sel0_b12/or_B21_B22_o , \NM/sel0_b12/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b12/or_or_or_B12_or_B13_  (\NM/sel0_b12/or_or_or_B12_or_B13__o , \NM/sel0_b12/or_or_B12_or_B13_B14_o , \NM/sel0_b12/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_11  (\NM/sel0_b13/B11 , M_result[0], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_12  (\NM/sel0_b13/B12 , M_result2[1], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_13  (\NM/sel0_b13/B13 , M_result2[2], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_14  (\NM/sel0_b13/B14 , M_result2[3], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_15  (\NM/sel0_b13/B15 , M_result2[4], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_16  (\NM/sel0_b13/B16 , M_result2[5], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_17  (\NM/sel0_b13/B17 , M_result2[6], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_18  (\NM/sel0_b13/B18 , M_result2[7], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_19  (\NM/sel0_b13/B19 , M_result2[8], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_20  (\NM/sel0_b13/B20 , M_result2[9], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_21  (\NM/sel0_b13/B21 , M_result2[10], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_22  (\NM/sel0_b13/B22 , M_result2[11], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_23  (\NM/sel0_b13/B23 , M_result2[12], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b13/and_b0_24  (\NM/sel0_b13/B24 , M_result2[13], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B12_or_B13_B14_o  (\NM/sel0_b13/or_B12_or_B13_B14_o_o , \NM/sel0_b13/B12 , \NM/sel0_b13/or_B13_B14_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B13_B14  (\NM/sel0_b13/or_B13_B14_o , \NM/sel0_b13/B13 , \NM/sel0_b13/B14 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B15_or_B16_B17_o  (\NM/sel0_b13/or_B15_or_B16_B17_o_o , \NM/sel0_b13/B15 , \NM/sel0_b13/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B16_B17  (\NM/sel0_b13/or_B16_B17_o , \NM/sel0_b13/B16 , \NM/sel0_b13/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B18_or_B19_B20_o  (\NM/sel0_b13/or_B18_or_B19_B20_o_o , \NM/sel0_b13/B18 , \NM/sel0_b13/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B19_B20  (\NM/sel0_b13/or_B19_B20_o , \NM/sel0_b13/B19 , \NM/sel0_b13/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B21_B22  (\NM/sel0_b13/or_B21_B22_o , \NM/sel0_b13/B21 , \NM/sel0_b13/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_B23_B24  (\NM/sel0_b13/or_B23_B24_o , \NM/sel0_b13/B23 , \NM/sel0_b13/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_or_B12_or_B13_B14  (\NM/sel0_b13/or_or_B12_or_B13_B14_o , \NM/sel0_b13/or_B12_or_B13_B14_o_o , \NM/sel0_b13/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_or_B18_or_B19_B20  (\NM/sel0_b13/or_or_B18_or_B19_B20_o , \NM/sel0_b13/or_B18_or_B19_B20_o_o , \NM/sel0_b13/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_or_B21_B22_o_or_B  (\NM/sel0_b13/or_or_B21_B22_o_or_B_o , \NM/sel0_b13/or_B21_B22_o , \NM/sel0_b13/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_or_or_B12_or_B13_  (\NM/sel0_b13/or_or_or_B12_or_B13__o , \NM/sel0_b13/or_or_B12_or_B13_B14_o , \NM/sel0_b13/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b13/or_or_or_or_B0_or_B1  (\NM/n122 [13], \NM/sel0_b13/B11 , \NM/sel0_b13/or_or_or_B12_or_B13__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_10  (\NM/sel0_b14/B10 , M_result[0], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_11  (\NM/sel0_b14/B11 , M_result2[1], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_12  (\NM/sel0_b14/B12 , M_result2[2], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_13  (\NM/sel0_b14/B13 , M_result2[3], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_14  (\NM/sel0_b14/B14 , M_result2[4], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_15  (\NM/sel0_b14/B15 , M_result2[5], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_16  (\NM/sel0_b14/B16 , M_result2[6], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_17  (\NM/sel0_b14/B17 , M_result2[7], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_18  (\NM/sel0_b14/B18 , M_result2[8], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_19  (\NM/sel0_b14/B19 , M_result2[9], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_20  (\NM/sel0_b14/B20 , M_result2[10], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_21  (\NM/sel0_b14/B21 , M_result2[11], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_22  (\NM/sel0_b14/B22 , M_result2[12], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_23  (\NM/sel0_b14/B23 , M_result2[13], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b14/and_b0_24  (\NM/sel0_b14/B24 , M_result2[14], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B10_B11  (\NM/sel0_b14/or_B10_B11_o , \NM/sel0_b14/B10 , \NM/sel0_b14/B11 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B12_or_B13_B14_o  (\NM/sel0_b14/or_B12_or_B13_B14_o_o , \NM/sel0_b14/B12 , \NM/sel0_b14/or_B13_B14_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B13_B14  (\NM/sel0_b14/or_B13_B14_o , \NM/sel0_b14/B13 , \NM/sel0_b14/B14 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B15_or_B16_B17_o  (\NM/sel0_b14/or_B15_or_B16_B17_o_o , \NM/sel0_b14/B15 , \NM/sel0_b14/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B16_B17  (\NM/sel0_b14/or_B16_B17_o , \NM/sel0_b14/B16 , \NM/sel0_b14/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B18_or_B19_B20_o  (\NM/sel0_b14/or_B18_or_B19_B20_o_o , \NM/sel0_b14/B18 , \NM/sel0_b14/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B19_B20  (\NM/sel0_b14/or_B19_B20_o , \NM/sel0_b14/B19 , \NM/sel0_b14/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B21_B22  (\NM/sel0_b14/or_B21_B22_o , \NM/sel0_b14/B21 , \NM/sel0_b14/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_B23_B24  (\NM/sel0_b14/or_B23_B24_o , \NM/sel0_b14/B23 , \NM/sel0_b14/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_or_B12_or_B13_B14  (\NM/sel0_b14/or_or_B12_or_B13_B14_o , \NM/sel0_b14/or_B12_or_B13_B14_o_o , \NM/sel0_b14/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_or_B18_or_B19_B20  (\NM/sel0_b14/or_or_B18_or_B19_B20_o , \NM/sel0_b14/or_B18_or_B19_B20_o_o , \NM/sel0_b14/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_or_B21_B22_o_or_B  (\NM/sel0_b14/or_or_B21_B22_o_or_B_o , \NM/sel0_b14/or_B21_B22_o , \NM/sel0_b14/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_or_or_B12_or_B13_  (\NM/sel0_b14/or_or_or_B12_or_B13__o , \NM/sel0_b14/or_or_B12_or_B13_B14_o , \NM/sel0_b14/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b14/or_or_or_or_B0_or_B1  (\NM/n122 [14], \NM/sel0_b14/or_B10_B11_o , \NM/sel0_b14/or_or_or_B12_or_B13__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_10  (\NM/sel0_b15/B10 , M_result2[1], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_11  (\NM/sel0_b15/B11 , M_result2[2], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_12  (\NM/sel0_b15/B12 , M_result2[3], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_13  (\NM/sel0_b15/B13 , M_result2[4], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_14  (\NM/sel0_b15/B14 , M_result2[5], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_15  (\NM/sel0_b15/B15 , M_result2[6], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_16  (\NM/sel0_b15/B16 , M_result2[7], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_17  (\NM/sel0_b15/B17 , M_result2[8], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_18  (\NM/sel0_b15/B18 , M_result2[9], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_19  (\NM/sel0_b15/B19 , M_result2[10], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_20  (\NM/sel0_b15/B20 , M_result2[11], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_21  (\NM/sel0_b15/B21 , M_result2[12], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_22  (\NM/sel0_b15/B22 , M_result2[13], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_23  (\NM/sel0_b15/B23 , M_result2[14], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_24  (\NM/sel0_b15/B24 , M_result2[15], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b15/and_b0_9  (\NM/sel0_b15/B9 , M_result[0], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B10_B11  (\NM/sel0_b15/or_B10_B11_o , \NM/sel0_b15/B10 , \NM/sel0_b15/B11 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B12_or_B13_B14_o  (\NM/sel0_b15/or_B12_or_B13_B14_o_o , \NM/sel0_b15/B12 , \NM/sel0_b15/or_B13_B14_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B13_B14  (\NM/sel0_b15/or_B13_B14_o , \NM/sel0_b15/B13 , \NM/sel0_b15/B14 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B15_or_B16_B17_o  (\NM/sel0_b15/or_B15_or_B16_B17_o_o , \NM/sel0_b15/B15 , \NM/sel0_b15/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B16_B17  (\NM/sel0_b15/or_B16_B17_o , \NM/sel0_b15/B16 , \NM/sel0_b15/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B18_or_B19_B20_o  (\NM/sel0_b15/or_B18_or_B19_B20_o_o , \NM/sel0_b15/B18 , \NM/sel0_b15/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B19_B20  (\NM/sel0_b15/or_B19_B20_o , \NM/sel0_b15/B19 , \NM/sel0_b15/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B21_B22  (\NM/sel0_b15/or_B21_B22_o , \NM/sel0_b15/B21 , \NM/sel0_b15/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B23_B24  (\NM/sel0_b15/or_B23_B24_o , \NM/sel0_b15/B23 , \NM/sel0_b15/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_B9_or_B10_B11_o  (\NM/sel0_b15/or_B9_or_B10_B11_o_o , \NM/sel0_b15/B9 , \NM/sel0_b15/or_B10_B11_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_or_B12_or_B13_B14  (\NM/sel0_b15/or_or_B12_or_B13_B14_o , \NM/sel0_b15/or_B12_or_B13_B14_o_o , \NM/sel0_b15/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_or_B18_or_B19_B20  (\NM/sel0_b15/or_or_B18_or_B19_B20_o , \NM/sel0_b15/or_B18_or_B19_B20_o_o , \NM/sel0_b15/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_or_B21_B22_o_or_B  (\NM/sel0_b15/or_or_B21_B22_o_or_B_o , \NM/sel0_b15/or_B21_B22_o , \NM/sel0_b15/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_or_or_B12_or_B13_  (\NM/sel0_b15/or_or_or_B12_or_B13__o , \NM/sel0_b15/or_or_B12_or_B13_B14_o , \NM/sel0_b15/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b15/or_or_or_or_B0_or_B1  (\NM/n122 [15], \NM/sel0_b15/or_B9_or_B10_B11_o_o , \NM/sel0_b15/or_or_or_B12_or_B13__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_10  (\NM/sel0_b16/B10 , M_result2[2], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_11  (\NM/sel0_b16/B11 , M_result2[3], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_12  (\NM/sel0_b16/B12 , M_result2[4], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_13  (\NM/sel0_b16/B13 , M_result2[5], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_14  (\NM/sel0_b16/B14 , M_result2[6], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_15  (\NM/sel0_b16/B15 , M_result2[7], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_16  (\NM/sel0_b16/B16 , M_result2[8], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_17  (\NM/sel0_b16/B17 , M_result2[9], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_18  (\NM/sel0_b16/B18 , M_result2[10], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_19  (\NM/sel0_b16/B19 , M_result2[11], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_20  (\NM/sel0_b16/B20 , M_result2[12], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_21  (\NM/sel0_b16/B21 , M_result2[13], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_22  (\NM/sel0_b16/B22 , M_result2[14], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_23  (\NM/sel0_b16/B23 , M_result2[15], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_24  (\NM/sel0_b16/B24 , M_result2[16], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_8  (\NM/sel0_b16/B8 , M_result[0], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b16/and_b0_9  (\NM/sel0_b16/B9 , M_result2[1], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B10_B11  (\NM/sel0_b16/or_B10_B11_o , \NM/sel0_b16/B10 , \NM/sel0_b16/B11 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B12_or_B13_B14_o  (\NM/sel0_b16/or_B12_or_B13_B14_o_o , \NM/sel0_b16/B12 , \NM/sel0_b16/or_B13_B14_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B13_B14  (\NM/sel0_b16/or_B13_B14_o , \NM/sel0_b16/B13 , \NM/sel0_b16/B14 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B15_or_B16_B17_o  (\NM/sel0_b16/or_B15_or_B16_B17_o_o , \NM/sel0_b16/B15 , \NM/sel0_b16/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B16_B17  (\NM/sel0_b16/or_B16_B17_o , \NM/sel0_b16/B16 , \NM/sel0_b16/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B18_or_B19_B20_o  (\NM/sel0_b16/or_B18_or_B19_B20_o_o , \NM/sel0_b16/B18 , \NM/sel0_b16/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B19_B20  (\NM/sel0_b16/or_B19_B20_o , \NM/sel0_b16/B19 , \NM/sel0_b16/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B21_B22  (\NM/sel0_b16/or_B21_B22_o , \NM/sel0_b16/B21 , \NM/sel0_b16/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B23_B24  (\NM/sel0_b16/or_B23_B24_o , \NM/sel0_b16/B23 , \NM/sel0_b16/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_B9_or_B10_B11_o  (\NM/sel0_b16/or_B9_or_B10_B11_o_o , \NM/sel0_b16/B9 , \NM/sel0_b16/or_B10_B11_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_or_B12_or_B13_B14  (\NM/sel0_b16/or_or_B12_or_B13_B14_o , \NM/sel0_b16/or_B12_or_B13_B14_o_o , \NM/sel0_b16/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_or_B18_or_B19_B20  (\NM/sel0_b16/or_or_B18_or_B19_B20_o , \NM/sel0_b16/or_B18_or_B19_B20_o_o , \NM/sel0_b16/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_or_B21_B22_o_or_B  (\NM/sel0_b16/or_or_B21_B22_o_or_B_o , \NM/sel0_b16/or_B21_B22_o , \NM/sel0_b16/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_or_B6_or_B7_B8_o_  (\NM/sel0_b16/or_or_B6_or_B7_B8_o__o , \NM/sel0_b16/B8 , \NM/sel0_b16/or_B9_or_B10_B11_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_or_or_B12_or_B13_  (\NM/sel0_b16/or_or_or_B12_or_B13__o , \NM/sel0_b16/or_or_B12_or_B13_B14_o , \NM/sel0_b16/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b16/or_or_or_or_B0_or_B1  (\NM/n122 [16], \NM/sel0_b16/or_or_B6_or_B7_B8_o__o , \NM/sel0_b16/or_or_or_B12_or_B13__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_10  (\NM/sel0_b17/B10 , M_result2[3], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_11  (\NM/sel0_b17/B11 , M_result2[4], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_12  (\NM/sel0_b17/B12 , M_result2[5], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_13  (\NM/sel0_b17/B13 , M_result2[6], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_14  (\NM/sel0_b17/B14 , M_result2[7], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_15  (\NM/sel0_b17/B15 , M_result2[8], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_16  (\NM/sel0_b17/B16 , M_result2[9], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_17  (\NM/sel0_b17/B17 , M_result2[10], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_18  (\NM/sel0_b17/B18 , M_result2[11], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_19  (\NM/sel0_b17/B19 , M_result2[12], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_20  (\NM/sel0_b17/B20 , M_result2[13], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_21  (\NM/sel0_b17/B21 , M_result2[14], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_22  (\NM/sel0_b17/B22 , M_result2[15], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_23  (\NM/sel0_b17/B23 , M_result2[16], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_24  (\NM/sel0_b17/B24 , M_result2[17], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_7  (\NM/sel0_b17/B7 , M_result[0], \NM/n101 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_8  (\NM/sel0_b17/B8 , M_result2[1], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b17/and_b0_9  (\NM/sel0_b17/B9 , M_result2[2], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B10_B11  (\NM/sel0_b17/or_B10_B11_o , \NM/sel0_b17/B10 , \NM/sel0_b17/B11 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B12_or_B13_B14_o  (\NM/sel0_b17/or_B12_or_B13_B14_o_o , \NM/sel0_b17/B12 , \NM/sel0_b17/or_B13_B14_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B13_B14  (\NM/sel0_b17/or_B13_B14_o , \NM/sel0_b17/B13 , \NM/sel0_b17/B14 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B15_or_B16_B17_o  (\NM/sel0_b17/or_B15_or_B16_B17_o_o , \NM/sel0_b17/B15 , \NM/sel0_b17/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B16_B17  (\NM/sel0_b17/or_B16_B17_o , \NM/sel0_b17/B16 , \NM/sel0_b17/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B18_or_B19_B20_o  (\NM/sel0_b17/or_B18_or_B19_B20_o_o , \NM/sel0_b17/B18 , \NM/sel0_b17/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B19_B20  (\NM/sel0_b17/or_B19_B20_o , \NM/sel0_b17/B19 , \NM/sel0_b17/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B21_B22  (\NM/sel0_b17/or_B21_B22_o , \NM/sel0_b17/B21 , \NM/sel0_b17/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B23_B24  (\NM/sel0_b17/or_B23_B24_o , \NM/sel0_b17/B23 , \NM/sel0_b17/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B7_B8  (\NM/sel0_b17/or_B7_B8_o , \NM/sel0_b17/B7 , \NM/sel0_b17/B8 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_B9_or_B10_B11_o  (\NM/sel0_b17/or_B9_or_B10_B11_o_o , \NM/sel0_b17/B9 , \NM/sel0_b17/or_B10_B11_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_or_B12_or_B13_B14  (\NM/sel0_b17/or_or_B12_or_B13_B14_o , \NM/sel0_b17/or_B12_or_B13_B14_o_o , \NM/sel0_b17/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_or_B18_or_B19_B20  (\NM/sel0_b17/or_or_B18_or_B19_B20_o , \NM/sel0_b17/or_B18_or_B19_B20_o_o , \NM/sel0_b17/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_or_B21_B22_o_or_B  (\NM/sel0_b17/or_or_B21_B22_o_or_B_o , \NM/sel0_b17/or_B21_B22_o , \NM/sel0_b17/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_or_B6_or_B7_B8_o_  (\NM/sel0_b17/or_or_B6_or_B7_B8_o__o , \NM/sel0_b17/or_B7_B8_o , \NM/sel0_b17/or_B9_or_B10_B11_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_or_or_B12_or_B13_  (\NM/sel0_b17/or_or_or_B12_or_B13__o , \NM/sel0_b17/or_or_B12_or_B13_B14_o , \NM/sel0_b17/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b17/or_or_or_or_B0_or_B1  (\NM/n122 [17], \NM/sel0_b17/or_or_B6_or_B7_B8_o__o , \NM/sel0_b17/or_or_or_B12_or_B13__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_10  (\NM/sel0_b18/B10 , M_result2[4], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_11  (\NM/sel0_b18/B11 , M_result2[5], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_12  (\NM/sel0_b18/B12 , M_result2[6], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_13  (\NM/sel0_b18/B13 , M_result2[7], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_14  (\NM/sel0_b18/B14 , M_result2[8], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_15  (\NM/sel0_b18/B15 , M_result2[9], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_16  (\NM/sel0_b18/B16 , M_result2[10], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_17  (\NM/sel0_b18/B17 , M_result2[11], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_18  (\NM/sel0_b18/B18 , M_result2[12], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_19  (\NM/sel0_b18/B19 , M_result2[13], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_20  (\NM/sel0_b18/B20 , M_result2[14], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_21  (\NM/sel0_b18/B21 , M_result2[15], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_22  (\NM/sel0_b18/B22 , M_result2[16], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_23  (\NM/sel0_b18/B23 , M_result2[17], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_24  (\NM/sel0_b18/B24 , M_result2[18], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_6  (\NM/sel0_b18/B6 , M_result[0], \NM/n104 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_7  (\NM/sel0_b18/B7 , M_result2[1], \NM/n101 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_8  (\NM/sel0_b18/B8 , M_result2[2], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b18/and_b0_9  (\NM/sel0_b18/B9 , M_result2[3], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B10_B11  (\NM/sel0_b18/or_B10_B11_o , \NM/sel0_b18/B10 , \NM/sel0_b18/B11 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B12_or_B13_B14_o  (\NM/sel0_b18/or_B12_or_B13_B14_o_o , \NM/sel0_b18/B12 , \NM/sel0_b18/or_B13_B14_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B13_B14  (\NM/sel0_b18/or_B13_B14_o , \NM/sel0_b18/B13 , \NM/sel0_b18/B14 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B15_or_B16_B17_o  (\NM/sel0_b18/or_B15_or_B16_B17_o_o , \NM/sel0_b18/B15 , \NM/sel0_b18/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B16_B17  (\NM/sel0_b18/or_B16_B17_o , \NM/sel0_b18/B16 , \NM/sel0_b18/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B18_or_B19_B20_o  (\NM/sel0_b18/or_B18_or_B19_B20_o_o , \NM/sel0_b18/B18 , \NM/sel0_b18/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B19_B20  (\NM/sel0_b18/or_B19_B20_o , \NM/sel0_b18/B19 , \NM/sel0_b18/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B21_B22  (\NM/sel0_b18/or_B21_B22_o , \NM/sel0_b18/B21 , \NM/sel0_b18/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B23_B24  (\NM/sel0_b18/or_B23_B24_o , \NM/sel0_b18/B23 , \NM/sel0_b18/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B6_or_B7_B8_o  (\NM/sel0_b18/or_B6_or_B7_B8_o_o , \NM/sel0_b18/B6 , \NM/sel0_b18/or_B7_B8_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B7_B8  (\NM/sel0_b18/or_B7_B8_o , \NM/sel0_b18/B7 , \NM/sel0_b18/B8 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_B9_or_B10_B11_o  (\NM/sel0_b18/or_B9_or_B10_B11_o_o , \NM/sel0_b18/B9 , \NM/sel0_b18/or_B10_B11_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_or_B12_or_B13_B14  (\NM/sel0_b18/or_or_B12_or_B13_B14_o , \NM/sel0_b18/or_B12_or_B13_B14_o_o , \NM/sel0_b18/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_or_B18_or_B19_B20  (\NM/sel0_b18/or_or_B18_or_B19_B20_o , \NM/sel0_b18/or_B18_or_B19_B20_o_o , \NM/sel0_b18/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_or_B21_B22_o_or_B  (\NM/sel0_b18/or_or_B21_B22_o_or_B_o , \NM/sel0_b18/or_B21_B22_o , \NM/sel0_b18/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_or_B6_or_B7_B8_o_  (\NM/sel0_b18/or_or_B6_or_B7_B8_o__o , \NM/sel0_b18/or_B6_or_B7_B8_o_o , \NM/sel0_b18/or_B9_or_B10_B11_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_or_or_B12_or_B13_  (\NM/sel0_b18/or_or_or_B12_or_B13__o , \NM/sel0_b18/or_or_B12_or_B13_B14_o , \NM/sel0_b18/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b18/or_or_or_or_B0_or_B1  (\NM/n122 [18], \NM/sel0_b18/or_or_B6_or_B7_B8_o__o , \NM/sel0_b18/or_or_or_B12_or_B13__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_10  (\NM/sel0_b19/B10 , M_result2[5], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_11  (\NM/sel0_b19/B11 , M_result2[6], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_12  (\NM/sel0_b19/B12 , M_result2[7], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_13  (\NM/sel0_b19/B13 , M_result2[8], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_14  (\NM/sel0_b19/B14 , M_result2[9], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_15  (\NM/sel0_b19/B15 , M_result2[10], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_16  (\NM/sel0_b19/B16 , M_result2[11], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_17  (\NM/sel0_b19/B17 , M_result2[12], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_18  (\NM/sel0_b19/B18 , M_result2[13], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_19  (\NM/sel0_b19/B19 , M_result2[14], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_20  (\NM/sel0_b19/B20 , M_result2[15], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_21  (\NM/sel0_b19/B21 , M_result2[16], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_22  (\NM/sel0_b19/B22 , M_result2[17], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_23  (\NM/sel0_b19/B23 , M_result2[18], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_24  (\NM/sel0_b19/B24 , M_result2[19], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_5  (\NM/sel0_b19/B5 , M_result[0], \NM/n107 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_6  (\NM/sel0_b19/B6 , M_result2[1], \NM/n104 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_7  (\NM/sel0_b19/B7 , M_result2[2], \NM/n101 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_8  (\NM/sel0_b19/B8 , M_result2[3], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b19/and_b0_9  (\NM/sel0_b19/B9 , M_result2[4], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B10_B11  (\NM/sel0_b19/or_B10_B11_o , \NM/sel0_b19/B10 , \NM/sel0_b19/B11 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B12_or_B13_B14_o  (\NM/sel0_b19/or_B12_or_B13_B14_o_o , \NM/sel0_b19/B12 , \NM/sel0_b19/or_B13_B14_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B13_B14  (\NM/sel0_b19/or_B13_B14_o , \NM/sel0_b19/B13 , \NM/sel0_b19/B14 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B15_or_B16_B17_o  (\NM/sel0_b19/or_B15_or_B16_B17_o_o , \NM/sel0_b19/B15 , \NM/sel0_b19/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B16_B17  (\NM/sel0_b19/or_B16_B17_o , \NM/sel0_b19/B16 , \NM/sel0_b19/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B18_or_B19_B20_o  (\NM/sel0_b19/or_B18_or_B19_B20_o_o , \NM/sel0_b19/B18 , \NM/sel0_b19/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B19_B20  (\NM/sel0_b19/or_B19_B20_o , \NM/sel0_b19/B19 , \NM/sel0_b19/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B21_B22  (\NM/sel0_b19/or_B21_B22_o , \NM/sel0_b19/B21 , \NM/sel0_b19/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B23_B24  (\NM/sel0_b19/or_B23_B24_o , \NM/sel0_b19/B23 , \NM/sel0_b19/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B6_or_B7_B8_o  (\NM/sel0_b19/or_B6_or_B7_B8_o_o , \NM/sel0_b19/B6 , \NM/sel0_b19/or_B7_B8_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B7_B8  (\NM/sel0_b19/or_B7_B8_o , \NM/sel0_b19/B7 , \NM/sel0_b19/B8 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_B9_or_B10_B11_o  (\NM/sel0_b19/or_B9_or_B10_B11_o_o , \NM/sel0_b19/B9 , \NM/sel0_b19/or_B10_B11_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_B12_or_B13_B14  (\NM/sel0_b19/or_or_B12_or_B13_B14_o , \NM/sel0_b19/or_B12_or_B13_B14_o_o , \NM/sel0_b19/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_B18_or_B19_B20  (\NM/sel0_b19/or_or_B18_or_B19_B20_o , \NM/sel0_b19/or_B18_or_B19_B20_o_o , \NM/sel0_b19/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_B21_B22_o_or_B  (\NM/sel0_b19/or_or_B21_B22_o_or_B_o , \NM/sel0_b19/or_B21_B22_o , \NM/sel0_b19/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_B6_or_B7_B8_o_  (\NM/sel0_b19/or_or_B6_or_B7_B8_o__o , \NM/sel0_b19/or_B6_or_B7_B8_o_o , \NM/sel0_b19/or_B9_or_B10_B11_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_or_B0_or_B1_B2  (\NM/sel0_b19/or_or_or_B0_or_B1_B2_o , \NM/sel0_b19/B5 , \NM/sel0_b19/or_or_B6_or_B7_B8_o__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_or_B12_or_B13_  (\NM/sel0_b19/or_or_or_B12_or_B13__o , \NM/sel0_b19/or_or_B12_or_B13_B14_o , \NM/sel0_b19/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b19/or_or_or_or_B0_or_B1  (\NM/n122 [19], \NM/sel0_b19/or_or_or_B0_or_B1_B2_o , \NM/sel0_b19/or_or_or_B12_or_B13__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b2/and_b0_22  (\NM/sel0_b2/B22 , M_result[0], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b2/and_b0_23  (\NM/sel0_b2/B23 , M_result2[1], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b2/and_b0_24  (\NM/sel0_b2/B24 , M_result2[2], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b2/or_B23_B24  (\NM/sel0_b2/or_B23_B24_o , \NM/sel0_b2/B23 , \NM/sel0_b2/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b2/or_or_B21_B22_o_or_B  (\NM/sel0_b2/or_or_B21_B22_o_or_B_o , \NM/sel0_b2/B22 , \NM/sel0_b2/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_10  (\NM/sel0_b20/B10 , M_result2[6], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_11  (\NM/sel0_b20/B11 , M_result2[7], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_12  (\NM/sel0_b20/B12 , M_result2[8], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_13  (\NM/sel0_b20/B13 , M_result2[9], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_14  (\NM/sel0_b20/B14 , M_result2[10], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_15  (\NM/sel0_b20/B15 , M_result2[11], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_16  (\NM/sel0_b20/B16 , M_result2[12], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_17  (\NM/sel0_b20/B17 , M_result2[13], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_18  (\NM/sel0_b20/B18 , M_result2[14], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_19  (\NM/sel0_b20/B19 , M_result2[15], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_20  (\NM/sel0_b20/B20 , M_result2[16], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_21  (\NM/sel0_b20/B21 , M_result2[17], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_22  (\NM/sel0_b20/B22 , M_result2[18], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_23  (\NM/sel0_b20/B23 , M_result2[19], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_24  (\NM/sel0_b20/B24 , M_result2[20], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_4  (\NM/sel0_b20/B4 , M_result[0], \NM/n110 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_5  (\NM/sel0_b20/B5 , M_result2[1], \NM/n107 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_6  (\NM/sel0_b20/B6 , M_result2[2], \NM/n104 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_7  (\NM/sel0_b20/B7 , M_result2[3], \NM/n101 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_8  (\NM/sel0_b20/B8 , M_result2[4], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b20/and_b0_9  (\NM/sel0_b20/B9 , M_result2[5], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B10_B11  (\NM/sel0_b20/or_B10_B11_o , \NM/sel0_b20/B10 , \NM/sel0_b20/B11 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B12_or_B13_B14_o  (\NM/sel0_b20/or_B12_or_B13_B14_o_o , \NM/sel0_b20/B12 , \NM/sel0_b20/or_B13_B14_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B13_B14  (\NM/sel0_b20/or_B13_B14_o , \NM/sel0_b20/B13 , \NM/sel0_b20/B14 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B15_or_B16_B17_o  (\NM/sel0_b20/or_B15_or_B16_B17_o_o , \NM/sel0_b20/B15 , \NM/sel0_b20/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B16_B17  (\NM/sel0_b20/or_B16_B17_o , \NM/sel0_b20/B16 , \NM/sel0_b20/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B18_or_B19_B20_o  (\NM/sel0_b20/or_B18_or_B19_B20_o_o , \NM/sel0_b20/B18 , \NM/sel0_b20/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B19_B20  (\NM/sel0_b20/or_B19_B20_o , \NM/sel0_b20/B19 , \NM/sel0_b20/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B21_B22  (\NM/sel0_b20/or_B21_B22_o , \NM/sel0_b20/B21 , \NM/sel0_b20/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B23_B24  (\NM/sel0_b20/or_B23_B24_o , \NM/sel0_b20/B23 , \NM/sel0_b20/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B4_B5  (\NM/sel0_b20/or_B4_B5_o , \NM/sel0_b20/B4 , \NM/sel0_b20/B5 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B6_or_B7_B8_o  (\NM/sel0_b20/or_B6_or_B7_B8_o_o , \NM/sel0_b20/B6 , \NM/sel0_b20/or_B7_B8_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B7_B8  (\NM/sel0_b20/or_B7_B8_o , \NM/sel0_b20/B7 , \NM/sel0_b20/B8 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_B9_or_B10_B11_o  (\NM/sel0_b20/or_B9_or_B10_B11_o_o , \NM/sel0_b20/B9 , \NM/sel0_b20/or_B10_B11_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_B12_or_B13_B14  (\NM/sel0_b20/or_or_B12_or_B13_B14_o , \NM/sel0_b20/or_B12_or_B13_B14_o_o , \NM/sel0_b20/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_B18_or_B19_B20  (\NM/sel0_b20/or_or_B18_or_B19_B20_o , \NM/sel0_b20/or_B18_or_B19_B20_o_o , \NM/sel0_b20/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_B21_B22_o_or_B  (\NM/sel0_b20/or_or_B21_B22_o_or_B_o , \NM/sel0_b20/or_B21_B22_o , \NM/sel0_b20/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_B6_or_B7_B8_o_  (\NM/sel0_b20/or_or_B6_or_B7_B8_o__o , \NM/sel0_b20/or_B6_or_B7_B8_o_o , \NM/sel0_b20/or_B9_or_B10_B11_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_or_B0_or_B1_B2  (\NM/sel0_b20/or_or_or_B0_or_B1_B2_o , \NM/sel0_b20/or_B4_B5_o , \NM/sel0_b20/or_or_B6_or_B7_B8_o__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_or_B12_or_B13_  (\NM/sel0_b20/or_or_or_B12_or_B13__o , \NM/sel0_b20/or_or_B12_or_B13_B14_o , \NM/sel0_b20/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b20/or_or_or_or_B0_or_B1  (\NM/n122 [20], \NM/sel0_b20/or_or_or_B0_or_B1_B2_o , \NM/sel0_b20/or_or_or_B12_or_B13__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_10  (\NM/sel0_b21/B10 , M_result2[7], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_11  (\NM/sel0_b21/B11 , M_result2[8], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_12  (\NM/sel0_b21/B12 , M_result2[9], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_13  (\NM/sel0_b21/B13 , M_result2[10], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_14  (\NM/sel0_b21/B14 , M_result2[11], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_15  (\NM/sel0_b21/B15 , M_result2[12], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_16  (\NM/sel0_b21/B16 , M_result2[13], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_17  (\NM/sel0_b21/B17 , M_result2[14], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_18  (\NM/sel0_b21/B18 , M_result2[15], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_19  (\NM/sel0_b21/B19 , M_result2[16], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_20  (\NM/sel0_b21/B20 , M_result2[17], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_21  (\NM/sel0_b21/B21 , M_result2[18], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_22  (\NM/sel0_b21/B22 , M_result2[19], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_23  (\NM/sel0_b21/B23 , M_result2[20], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_24  (\NM/sel0_b21/B24 , M_result2[21], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_3  (\NM/sel0_b21/B3 , M_result[0], \NM/n113 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_4  (\NM/sel0_b21/B4 , M_result2[1], \NM/n110 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_5  (\NM/sel0_b21/B5 , M_result2[2], \NM/n107 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_6  (\NM/sel0_b21/B6 , M_result2[3], \NM/n104 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_7  (\NM/sel0_b21/B7 , M_result2[4], \NM/n101 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_8  (\NM/sel0_b21/B8 , M_result2[5], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b21/and_b0_9  (\NM/sel0_b21/B9 , M_result2[6], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B10_B11  (\NM/sel0_b21/or_B10_B11_o , \NM/sel0_b21/B10 , \NM/sel0_b21/B11 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B12_or_B13_B14_o  (\NM/sel0_b21/or_B12_or_B13_B14_o_o , \NM/sel0_b21/B12 , \NM/sel0_b21/or_B13_B14_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B13_B14  (\NM/sel0_b21/or_B13_B14_o , \NM/sel0_b21/B13 , \NM/sel0_b21/B14 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B15_or_B16_B17_o  (\NM/sel0_b21/or_B15_or_B16_B17_o_o , \NM/sel0_b21/B15 , \NM/sel0_b21/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B16_B17  (\NM/sel0_b21/or_B16_B17_o , \NM/sel0_b21/B16 , \NM/sel0_b21/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B18_or_B19_B20_o  (\NM/sel0_b21/or_B18_or_B19_B20_o_o , \NM/sel0_b21/B18 , \NM/sel0_b21/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B19_B20  (\NM/sel0_b21/or_B19_B20_o , \NM/sel0_b21/B19 , \NM/sel0_b21/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B21_B22  (\NM/sel0_b21/or_B21_B22_o , \NM/sel0_b21/B21 , \NM/sel0_b21/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B23_B24  (\NM/sel0_b21/or_B23_B24_o , \NM/sel0_b21/B23 , \NM/sel0_b21/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B3_or_B4_B5_o  (\NM/sel0_b21/or_B3_or_B4_B5_o_o , \NM/sel0_b21/B3 , \NM/sel0_b21/or_B4_B5_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B4_B5  (\NM/sel0_b21/or_B4_B5_o , \NM/sel0_b21/B4 , \NM/sel0_b21/B5 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B6_or_B7_B8_o  (\NM/sel0_b21/or_B6_or_B7_B8_o_o , \NM/sel0_b21/B6 , \NM/sel0_b21/or_B7_B8_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B7_B8  (\NM/sel0_b21/or_B7_B8_o , \NM/sel0_b21/B7 , \NM/sel0_b21/B8 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_B9_or_B10_B11_o  (\NM/sel0_b21/or_B9_or_B10_B11_o_o , \NM/sel0_b21/B9 , \NM/sel0_b21/or_B10_B11_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_B12_or_B13_B14  (\NM/sel0_b21/or_or_B12_or_B13_B14_o , \NM/sel0_b21/or_B12_or_B13_B14_o_o , \NM/sel0_b21/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_B18_or_B19_B20  (\NM/sel0_b21/or_or_B18_or_B19_B20_o , \NM/sel0_b21/or_B18_or_B19_B20_o_o , \NM/sel0_b21/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_B21_B22_o_or_B  (\NM/sel0_b21/or_or_B21_B22_o_or_B_o , \NM/sel0_b21/or_B21_B22_o , \NM/sel0_b21/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_B6_or_B7_B8_o_  (\NM/sel0_b21/or_or_B6_or_B7_B8_o__o , \NM/sel0_b21/or_B6_or_B7_B8_o_o , \NM/sel0_b21/or_B9_or_B10_B11_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_or_B0_or_B1_B2  (\NM/sel0_b21/or_or_or_B0_or_B1_B2_o , \NM/sel0_b21/or_B3_or_B4_B5_o_o , \NM/sel0_b21/or_or_B6_or_B7_B8_o__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_or_B12_or_B13_  (\NM/sel0_b21/or_or_or_B12_or_B13__o , \NM/sel0_b21/or_or_B12_or_B13_B14_o , \NM/sel0_b21/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b21/or_or_or_or_B0_or_B1  (\NM/n122 [21], \NM/sel0_b21/or_or_or_B0_or_B1_B2_o , \NM/sel0_b21/or_or_or_B12_or_B13__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_10  (\NM/sel0_b22/B10 , M_result2[8], \NM/n92 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_11  (\NM/sel0_b22/B11 , M_result2[9], \NM/n89 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_12  (\NM/sel0_b22/B12 , M_result2[10], \NM/n86 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_13  (\NM/sel0_b22/B13 , M_result2[11], \NM/n83 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_14  (\NM/sel0_b22/B14 , M_result2[12], \NM/n80 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_15  (\NM/sel0_b22/B15 , M_result2[13], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_16  (\NM/sel0_b22/B16 , M_result2[14], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_17  (\NM/sel0_b22/B17 , M_result2[15], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_18  (\NM/sel0_b22/B18 , M_result2[16], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_19  (\NM/sel0_b22/B19 , M_result2[17], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_2  (\NM/sel0_b22/B2 , M_result[0], \NM/n116 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_20  (\NM/sel0_b22/B20 , M_result2[18], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_21  (\NM/sel0_b22/B21 , M_result2[19], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_22  (\NM/sel0_b22/B22 , M_result2[20], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_23  (\NM/sel0_b22/B23 , M_result2[21], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_24  (\NM/sel0_b22/B24 , M_result2[22], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_3  (\NM/sel0_b22/B3 , M_result2[1], \NM/n113 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_4  (\NM/sel0_b22/B4 , M_result2[2], \NM/n110 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_5  (\NM/sel0_b22/B5 , M_result2[3], \NM/n107 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_6  (\NM/sel0_b22/B6 , M_result2[4], \NM/n104 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_7  (\NM/sel0_b22/B7 , M_result2[5], \NM/n101 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_8  (\NM/sel0_b22/B8 , M_result2[6], \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b22/and_b0_9  (\NM/sel0_b22/B9 , M_result2[7], \NM/n95 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B10_B11  (\NM/sel0_b22/or_B10_B11_o , \NM/sel0_b22/B10 , \NM/sel0_b22/B11 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B12_or_B13_B14_o  (\NM/sel0_b22/or_B12_or_B13_B14_o_o , \NM/sel0_b22/B12 , \NM/sel0_b22/or_B13_B14_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B13_B14  (\NM/sel0_b22/or_B13_B14_o , \NM/sel0_b22/B13 , \NM/sel0_b22/B14 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B15_or_B16_B17_o  (\NM/sel0_b22/or_B15_or_B16_B17_o_o , \NM/sel0_b22/B15 , \NM/sel0_b22/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B16_B17  (\NM/sel0_b22/or_B16_B17_o , \NM/sel0_b22/B16 , \NM/sel0_b22/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B18_or_B19_B20_o  (\NM/sel0_b22/or_B18_or_B19_B20_o_o , \NM/sel0_b22/B18 , \NM/sel0_b22/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B19_B20  (\NM/sel0_b22/or_B19_B20_o , \NM/sel0_b22/B19 , \NM/sel0_b22/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B21_B22  (\NM/sel0_b22/or_B21_B22_o , \NM/sel0_b22/B21 , \NM/sel0_b22/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B23_B24  (\NM/sel0_b22/or_B23_B24_o , \NM/sel0_b22/B23 , \NM/sel0_b22/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B3_or_B4_B5_o  (\NM/sel0_b22/or_B3_or_B4_B5_o_o , \NM/sel0_b22/B3 , \NM/sel0_b22/or_B4_B5_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B4_B5  (\NM/sel0_b22/or_B4_B5_o , \NM/sel0_b22/B4 , \NM/sel0_b22/B5 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B6_or_B7_B8_o  (\NM/sel0_b22/or_B6_or_B7_B8_o_o , \NM/sel0_b22/B6 , \NM/sel0_b22/or_B7_B8_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B7_B8  (\NM/sel0_b22/or_B7_B8_o , \NM/sel0_b22/B7 , \NM/sel0_b22/B8 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_B9_or_B10_B11_o  (\NM/sel0_b22/or_B9_or_B10_B11_o_o , \NM/sel0_b22/B9 , \NM/sel0_b22/or_B10_B11_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_B0_or_B1_B2_o_  (\NM/sel0_b22/or_or_B0_or_B1_B2_o__o , \NM/sel0_b22/B2 , \NM/sel0_b22/or_B3_or_B4_B5_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_B12_or_B13_B14  (\NM/sel0_b22/or_or_B12_or_B13_B14_o , \NM/sel0_b22/or_B12_or_B13_B14_o_o , \NM/sel0_b22/or_B15_or_B16_B17_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_B18_or_B19_B20  (\NM/sel0_b22/or_or_B18_or_B19_B20_o , \NM/sel0_b22/or_B18_or_B19_B20_o_o , \NM/sel0_b22/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_B21_B22_o_or_B  (\NM/sel0_b22/or_or_B21_B22_o_or_B_o , \NM/sel0_b22/or_B21_B22_o , \NM/sel0_b22/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_B6_or_B7_B8_o_  (\NM/sel0_b22/or_or_B6_or_B7_B8_o__o , \NM/sel0_b22/or_B6_or_B7_B8_o_o , \NM/sel0_b22/or_B9_or_B10_B11_o_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_or_B0_or_B1_B2  (\NM/sel0_b22/or_or_or_B0_or_B1_B2_o , \NM/sel0_b22/or_or_B0_or_B1_B2_o__o , \NM/sel0_b22/or_or_B6_or_B7_B8_o__o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_or_B12_or_B13_  (\NM/sel0_b22/or_or_or_B12_or_B13__o , \NM/sel0_b22/or_or_B12_or_B13_B14_o , \NM/sel0_b22/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b22/or_or_or_or_B0_or_B1  (\NM/n122 [22], \NM/sel0_b22/or_or_or_B0_or_B1_B2_o , \NM/sel0_b22/or_or_or_B12_or_B13__o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b3/and_b0_21  (\NM/sel0_b3/B21 , M_result[0], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b3/and_b0_22  (\NM/sel0_b3/B22 , M_result2[1], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b3/and_b0_23  (\NM/sel0_b3/B23 , M_result2[2], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b3/and_b0_24  (\NM/sel0_b3/B24 , M_result2[3], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b3/or_B21_B22  (\NM/sel0_b3/or_B21_B22_o , \NM/sel0_b3/B21 , \NM/sel0_b3/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b3/or_B23_B24  (\NM/sel0_b3/or_B23_B24_o , \NM/sel0_b3/B23 , \NM/sel0_b3/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b3/or_or_B21_B22_o_or_B  (\NM/sel0_b3/or_or_B21_B22_o_or_B_o , \NM/sel0_b3/or_B21_B22_o , \NM/sel0_b3/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b4/and_b0_20  (\NM/sel0_b4/B20 , M_result[0], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b4/and_b0_21  (\NM/sel0_b4/B21 , M_result2[1], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b4/and_b0_22  (\NM/sel0_b4/B22 , M_result2[2], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b4/and_b0_23  (\NM/sel0_b4/B23 , M_result2[3], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b4/and_b0_24  (\NM/sel0_b4/B24 , M_result2[4], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b4/or_B21_B22  (\NM/sel0_b4/or_B21_B22_o , \NM/sel0_b4/B21 , \NM/sel0_b4/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b4/or_B23_B24  (\NM/sel0_b4/or_B23_B24_o , \NM/sel0_b4/B23 , \NM/sel0_b4/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b4/or_or_B18_or_B19_B20  (\NM/sel0_b4/or_or_B18_or_B19_B20_o , \NM/sel0_b4/B20 , \NM/sel0_b4/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b4/or_or_B21_B22_o_or_B  (\NM/sel0_b4/or_or_B21_B22_o_or_B_o , \NM/sel0_b4/or_B21_B22_o , \NM/sel0_b4/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b5/and_b0_19  (\NM/sel0_b5/B19 , M_result[0], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b5/and_b0_20  (\NM/sel0_b5/B20 , M_result2[1], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b5/and_b0_21  (\NM/sel0_b5/B21 , M_result2[2], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b5/and_b0_22  (\NM/sel0_b5/B22 , M_result2[3], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b5/and_b0_23  (\NM/sel0_b5/B23 , M_result2[4], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b5/and_b0_24  (\NM/sel0_b5/B24 , M_result2[5], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b5/or_B19_B20  (\NM/sel0_b5/or_B19_B20_o , \NM/sel0_b5/B19 , \NM/sel0_b5/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b5/or_B21_B22  (\NM/sel0_b5/or_B21_B22_o , \NM/sel0_b5/B21 , \NM/sel0_b5/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b5/or_B23_B24  (\NM/sel0_b5/or_B23_B24_o , \NM/sel0_b5/B23 , \NM/sel0_b5/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b5/or_or_B18_or_B19_B20  (\NM/sel0_b5/or_or_B18_or_B19_B20_o , \NM/sel0_b5/or_B19_B20_o , \NM/sel0_b5/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b5/or_or_B21_B22_o_or_B  (\NM/sel0_b5/or_or_B21_B22_o_or_B_o , \NM/sel0_b5/or_B21_B22_o , \NM/sel0_b5/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_18  (\NM/sel0_b6/B18 , M_result[0], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_19  (\NM/sel0_b6/B19 , M_result2[1], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_20  (\NM/sel0_b6/B20 , M_result2[2], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_21  (\NM/sel0_b6/B21 , M_result2[3], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_22  (\NM/sel0_b6/B22 , M_result2[4], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_23  (\NM/sel0_b6/B23 , M_result2[5], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b6/and_b0_24  (\NM/sel0_b6/B24 , M_result2[6], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b6/or_B18_or_B19_B20_o  (\NM/sel0_b6/or_B18_or_B19_B20_o_o , \NM/sel0_b6/B18 , \NM/sel0_b6/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b6/or_B19_B20  (\NM/sel0_b6/or_B19_B20_o , \NM/sel0_b6/B19 , \NM/sel0_b6/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b6/or_B21_B22  (\NM/sel0_b6/or_B21_B22_o , \NM/sel0_b6/B21 , \NM/sel0_b6/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b6/or_B23_B24  (\NM/sel0_b6/or_B23_B24_o , \NM/sel0_b6/B23 , \NM/sel0_b6/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b6/or_or_B18_or_B19_B20  (\NM/sel0_b6/or_or_B18_or_B19_B20_o , \NM/sel0_b6/or_B18_or_B19_B20_o_o , \NM/sel0_b6/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b6/or_or_B21_B22_o_or_B  (\NM/sel0_b6/or_or_B21_B22_o_or_B_o , \NM/sel0_b6/or_B21_B22_o , \NM/sel0_b6/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_17  (\NM/sel0_b7/B17 , M_result[0], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_18  (\NM/sel0_b7/B18 , M_result2[1], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_19  (\NM/sel0_b7/B19 , M_result2[2], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_20  (\NM/sel0_b7/B20 , M_result2[3], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_21  (\NM/sel0_b7/B21 , M_result2[4], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_22  (\NM/sel0_b7/B22 , M_result2[5], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_23  (\NM/sel0_b7/B23 , M_result2[6], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b7/and_b0_24  (\NM/sel0_b7/B24 , M_result2[7], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_B18_or_B19_B20_o  (\NM/sel0_b7/or_B18_or_B19_B20_o_o , \NM/sel0_b7/B18 , \NM/sel0_b7/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_B19_B20  (\NM/sel0_b7/or_B19_B20_o , \NM/sel0_b7/B19 , \NM/sel0_b7/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_B21_B22  (\NM/sel0_b7/or_B21_B22_o , \NM/sel0_b7/B21 , \NM/sel0_b7/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_B23_B24  (\NM/sel0_b7/or_B23_B24_o , \NM/sel0_b7/B23 , \NM/sel0_b7/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_or_B18_or_B19_B20  (\NM/sel0_b7/or_or_B18_or_B19_B20_o , \NM/sel0_b7/or_B18_or_B19_B20_o_o , \NM/sel0_b7/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_or_B21_B22_o_or_B  (\NM/sel0_b7/or_or_B21_B22_o_or_B_o , \NM/sel0_b7/or_B21_B22_o , \NM/sel0_b7/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b7/or_or_or_B12_or_B13_  (\NM/sel0_b7/or_or_or_B12_or_B13__o , \NM/sel0_b7/B17 , \NM/sel0_b7/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_16  (\NM/sel0_b8/B16 , M_result[0], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_17  (\NM/sel0_b8/B17 , M_result2[1], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_18  (\NM/sel0_b8/B18 , M_result2[2], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_19  (\NM/sel0_b8/B19 , M_result2[3], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_20  (\NM/sel0_b8/B20 , M_result2[4], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_21  (\NM/sel0_b8/B21 , M_result2[5], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_22  (\NM/sel0_b8/B22 , M_result2[6], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_23  (\NM/sel0_b8/B23 , M_result2[7], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b8/and_b0_24  (\NM/sel0_b8/B24 , M_result2[8], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_B16_B17  (\NM/sel0_b8/or_B16_B17_o , \NM/sel0_b8/B16 , \NM/sel0_b8/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_B18_or_B19_B20_o  (\NM/sel0_b8/or_B18_or_B19_B20_o_o , \NM/sel0_b8/B18 , \NM/sel0_b8/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_B19_B20  (\NM/sel0_b8/or_B19_B20_o , \NM/sel0_b8/B19 , \NM/sel0_b8/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_B21_B22  (\NM/sel0_b8/or_B21_B22_o , \NM/sel0_b8/B21 , \NM/sel0_b8/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_B23_B24  (\NM/sel0_b8/or_B23_B24_o , \NM/sel0_b8/B23 , \NM/sel0_b8/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_or_B18_or_B19_B20  (\NM/sel0_b8/or_or_B18_or_B19_B20_o , \NM/sel0_b8/or_B18_or_B19_B20_o_o , \NM/sel0_b8/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_or_B21_B22_o_or_B  (\NM/sel0_b8/or_or_B21_B22_o_or_B_o , \NM/sel0_b8/or_B21_B22_o , \NM/sel0_b8/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b8/or_or_or_B12_or_B13_  (\NM/sel0_b8/or_or_or_B12_or_B13__o , \NM/sel0_b8/or_B16_B17_o , \NM/sel0_b8/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_15  (\NM/sel0_b9/B15 , M_result[0], \NM/n77 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_16  (\NM/sel0_b9/B16 , M_result2[1], \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_17  (\NM/sel0_b9/B17 , M_result2[2], \NM/n71 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_18  (\NM/sel0_b9/B18 , M_result2[3], \NM/n68 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_19  (\NM/sel0_b9/B19 , M_result2[4], \NM/n65 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_20  (\NM/sel0_b9/B20 , M_result2[5], \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_21  (\NM/sel0_b9/B21 , M_result2[6], \NM/n59 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_22  (\NM/sel0_b9/B22 , M_result2[7], \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_23  (\NM/sel0_b9/B23 , M_result2[8], \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/sel0_b9/and_b0_24  (\NM/sel0_b9/B24 , M_result2[9], M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_B15_or_B16_B17_o  (\NM/sel0_b9/or_B15_or_B16_B17_o_o , \NM/sel0_b9/B15 , \NM/sel0_b9/or_B16_B17_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_B16_B17  (\NM/sel0_b9/or_B16_B17_o , \NM/sel0_b9/B16 , \NM/sel0_b9/B17 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_B18_or_B19_B20_o  (\NM/sel0_b9/or_B18_or_B19_B20_o_o , \NM/sel0_b9/B18 , \NM/sel0_b9/or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_B19_B20  (\NM/sel0_b9/or_B19_B20_o , \NM/sel0_b9/B19 , \NM/sel0_b9/B20 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_B21_B22  (\NM/sel0_b9/or_B21_B22_o , \NM/sel0_b9/B21 , \NM/sel0_b9/B22 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_B23_B24  (\NM/sel0_b9/or_B23_B24_o , \NM/sel0_b9/B23 , \NM/sel0_b9/B24 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_or_B18_or_B19_B20  (\NM/sel0_b9/or_or_B18_or_B19_B20_o , \NM/sel0_b9/or_B18_or_B19_B20_o_o , \NM/sel0_b9/or_or_B21_B22_o_or_B_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_or_B21_B22_o_or_B  (\NM/sel0_b9/or_or_B21_B22_o_or_B_o , \NM/sel0_b9/or_B21_B22_o , \NM/sel0_b9/or_B23_B24_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel0_b9/or_or_or_B12_or_B13_  (\NM/sel0_b9/or_or_or_B12_or_B13__o , \NM/sel0_b9/or_B15_or_B16_B17_o_o , \NM/sel0_b9/or_or_B18_or_B19_B20_o );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel1_b0_sel  (\NM/sel1_b0_sel_o , \NM/n119 , \NM/n113 , \NM/n107 , \NM/n101 , \NM/n95 , \NM/n89 , \NM/n83 , \NM/n77 , \NM/n71 , \NM/n65 , \NM/n59 , \NM/n53 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel1_b1_sel  (\NM/sel1_b1_sel_o , \NM/n119 , \NM/n116 , \NM/n107 , \NM/n104 , \NM/n95 , \NM/n92 , \NM/n83 , \NM/n80 , \NM/n71 , \NM/n68 , \NM/n59 , \NM/n56 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel1_b2_sel  (\NM/sel1_b2_sel_o , \NM/n119 , \NM/n116 , \NM/n113 , \NM/n110 , \NM/n95 , \NM/n92 , \NM/n89 , \NM/n86 , \NM/n71 , \NM/n68 , \NM/n65 , \NM/n62 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel1_b3_sel  (\NM/sel1_b3_sel_o , \NM/n95 , \NM/n92 , \NM/n89 , \NM/n86 , \NM/n83 , \NM/n80 , \NM/n77 , \NM/n74 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/sel1_b4_sel  (\NM/sel1_b4_sel_o , \NM/n119 , \NM/n116 , \NM/n113 , \NM/n110 , \NM/n107 , \NM/n104 , \NM/n101 , \NM/n98 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u10  (\NM/n10 , M_result2[20]);  // ../RTL/core/fpu_utils.v(181)
  and \NM/u100  (\NM/n101 , \NM/n39 , \NM/n100 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u101  (\NM/n102 , \NM/n99 , \NM/n39 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u102  (\NM/n103 , \NM/n102 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u103  (\NM/n104 , \NM/n41 , \NM/n103 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u104  (\NM/n105 , \NM/n102 , \NM/n41 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u105  (\NM/n106 , \NM/n105 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u106  (\NM/n107 , \NM/n44 , \NM/n106 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u107  (\NM/n108 , \NM/n105 , \NM/n44 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u108  (\NM/n109 , \NM/n108 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u109  (\NM/n110 , \NM/n46 , \NM/n109 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u11  (\NM/n374 , M_result2[22], M_result2[23]);  // ../RTL/core/fpu_utils.v(175)
  or \NM/u110  (\NM/n111 , \NM/n108 , \NM/n46 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u111  (\NM/n112 , \NM/n111 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u112  (\NM/n113 , \NM/n48 , \NM/n112 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u113  (\NM/n114 , \NM/n111 , \NM/n48 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u114  (\NM/n115 , \NM/n114 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u115  (\NM/n116 , \NM/n50 , \NM/n115 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u116  (\NM/n117 , \NM/n114 , \NM/n50 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u117  (\NM/n118 , \NM/n117 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u118  (\NM/n119 , \NM/n51 , \NM/n118 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u12  (\NM/n12 , M_result2[19]);  // ../RTL/core/fpu_utils.v(187)
  or \NM/u121  (\NM/n124 , M_result2[18], M_result2[19]);  // ../RTL/core/fpu_utils.v(253)
  or \NM/u122  (\NM/n125 , M_result2[16], M_result2[17]);  // ../RTL/core/fpu_utils.v(253)
  or \NM/u123  (\NM/n126 , \NM/n130 , \NM/n127 );  // ../RTL/core/fpu_utils.v(253)
  or \NM/u126  (\NM/n318 , M_result2[4], M_result2[5]);  // ../RTL/core/fpu_utils.v(295)
  or \NM/u127  (\NM/n279 , M_result2[4], \NM/n281 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u128  (\NM/n179 , \NM/n182 , \NM/n180 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u129  (\NM/n127 , \NM/n129 , \NM/n128 );  // ../RTL/core/fpu_utils.v(253)
  or \NM/u13  (\NM/n371 , \NM/n10 , M_result2[21]);  // ../RTL/core/fpu_utils.v(181)
  or \NM/u130  (\NM/n180 , M_result2[21], \NM/n374 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u132  (\NM/n316 , M_result2[3], \NM/n318 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u133  (\NM/n278 , \NM/n283 , \NM/n279 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u134  (\NM/n182 , M_result2[19], M_result2[20]);  // ../RTL/core/fpu_utils.v(265)
  or \NM/u135  (\NM/n128 , M_result2[14], M_result2[15]);  // ../RTL/core/fpu_utils.v(253)
  or \NM/u136  (\NM/n183 , \NM/n185 , \NM/n184 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u137  (\NM/n184 , M_result2[17], M_result2[18]);  // ../RTL/core/fpu_utils.v(265)
  or \NM/u138  (\NM/n314 , \NM/n319 , \NM/n316 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u139  (\NM/n276 , M_result2[8], M_result2[9]);  // ../RTL/core/fpu_utils.v(289)
  not \NM/u14  (\NM/n14 , M_result2[18]);  // ../RTL/core/fpu_utils.v(193)
  or \NM/u140  (\NM/n185 , M_result2[15], M_result2[16]);  // ../RTL/core/fpu_utils.v(265)
  or \NM/u141  (\NM/n129 , M_result2[12], M_result2[13]);  // ../RTL/core/fpu_utils.v(253)
  or \NM/u142  (\NM/n186 , \NM/n191 , \NM/n187 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u143  (\NM/n187 , \NM/n190 , \NM/n188 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u144  (\NM/n313 , M_result2[7], M_result2[8]);  // ../RTL/core/fpu_utils.v(295)
  or \NM/u145  (\NM/n274 , M_result2[7], \NM/n276 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u146  (\NM/n188 , M_result2[12], \NM/n189 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u147  (\NM/n130 , \NM/n132 , \NM/n190 );  // ../RTL/core/fpu_utils.v(253)
  or \NM/u148  (\NM/n189 , M_result2[13], M_result2[14]);  // ../RTL/core/fpu_utils.v(265)
  or \NM/u149  (\NM/n190 , M_result2[10], M_result2[11]);  // ../RTL/core/fpu_utils.v(265)
  or \NM/u15  (\NM/n367 , \NM/n12 , M_result2[20]);  // ../RTL/core/fpu_utils.v(187)
  or \NM/u150  (\NM/n311 , M_result2[6], \NM/n313 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u151  (\NM/n273 , M_result2[11], M_result2[12]);  // ../RTL/core/fpu_utils.v(289)
  or \NM/u152  (\NM/n191 , \NM/n193 , \NM/n276 );  // ../RTL/core/fpu_utils.v(265)
  not \NM/u155  (\NM/n41 , \NM/n194 );  // ../RTL/core/fpu_utils.v(271)
  or \NM/u157  (\NM/n271 , M_result2[10], \NM/n273 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u158  (\NM/n194 , \NM/n222 , \NM/n195 );  // ../RTL/core/fpu_utils.v(271)
  not \NM/u159  (\NM/n37 , \NM/n133 );  // ../RTL/core/fpu_utils.v(259)
  not \NM/u16  (\NM/n16 , M_result2[17]);  // ../RTL/core/fpu_utils.v(199)
  or \NM/u160  (\NM/n195 , \NM/n202 , \NM/n179 );  // ../RTL/core/fpu_utils.v(271)
  or \NM/u162  (\NM/n308 , M_result2[9], \NM/n190 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u163  (\NM/n269 , \NM/n274 , \NM/n271 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u165  (\NM/n133 , \NM/n142 , \NM/n134 );  // ../RTL/core/fpu_utils.v(259)
  or \NM/u168  (\NM/n306 , \NM/n311 , \NM/n308 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u169  (\NM/n268 , \NM/n278 , \NM/n269 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u170  (\NM/n202 , \NM/n128 , \NM/n207 );  // ../RTL/core/fpu_utils.v(271)
  or \NM/u171  (\NM/n134 , \NM/n183 , \NM/n179 );  // ../RTL/core/fpu_utils.v(259)
  or \NM/u172  (\NM/n207 , M_result2[16], \NM/n184 );  // ../RTL/core/fpu_utils.v(271)
  or \NM/u174  (\NM/n304 , \NM/n314 , \NM/n306 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u178  (\NM/n222 , \NM/n247 , \NM/n227 );  // ../RTL/core/fpu_utils.v(271)
  or \NM/u179  (\NM/n227 , \NM/n242 , \NM/n232 );  // ../RTL/core/fpu_utils.v(271)
  not \NM/u18  (\NM/n18 , M_result2[16]);  // ../RTL/core/fpu_utils.v(205)
  or \NM/u182  (\NM/n232 , M_result2[11], \NM/n129 );  // ../RTL/core/fpu_utils.v(271)
  or \NM/u185  (\NM/n242 , M_result2[9], M_result2[10]);  // ../RTL/core/fpu_utils.v(271)
  or \NM/u187  (\NM/n263 , M_result2[15], \NM/n125 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u188  (\NM/n247 , \NM/n257 , \NM/n313 );  // ../RTL/core/fpu_utils.v(271)
  not \NM/u191  (\NM/n44 , \NM/n262 );  // ../RTL/core/fpu_utils.v(277)
  or \NM/u193  (\NM/n261 , \NM/n189 , \NM/n263 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u194  (\NM/n262 , \NM/n312 , \NM/n195 );  // ../RTL/core/fpu_utils.v(277)
  not \NM/u20  (\NM/n20 , M_result2[15]);  // ../RTL/core/fpu_utils.v(211)
  or \NM/u204  (\NM/n296 , \NM/n188 , \NM/n263 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u205  (\NM/n258 , M_result2[18], \NM/n182 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u21  (\NM/n349 , \NM/n18 , M_result2[17]);  // ../RTL/core/fpu_utils.v(205)
  or \NM/u214  (\NM/n312 , \NM/n209 , \NM/n227 );  // ../RTL/core/fpu_utils.v(277)
  or \NM/u219  (\NM/n142 , \NM/n146 , \NM/n143 );  // ../RTL/core/fpu_utils.v(259)
  not \NM/u22  (\NM/n22 , M_result2[14]);  // ../RTL/core/fpu_utils.v(217)
  or \NM/u223  (\NM/n253 , \NM/n258 , \NM/n180 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u224  (\NM/n209 , \NM/n214 , \NM/n211 );  // ../RTL/core/fpu_utils.v(277)
  or \NM/u225  (\NM/n143 , \NM/n273 , \NM/n189 );  // ../RTL/core/fpu_utils.v(259)
  or \NM/u226  (\NM/n211 , M_result2[6], \NM/n213 );  // ../RTL/core/fpu_utils.v(277)
  or \NM/u227  (\NM/n213 , M_result2[7], \NM/n34 );  // ../RTL/core/fpu_utils.v(277)
  or \NM/u229  (\NM/n251 , \NM/n261 , \NM/n253 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u23  (\NM/n341 , \NM/n20 , M_result2[16]);  // ../RTL/core/fpu_utils.v(211)
  not \NM/u230  (\NM/n46 , \NM/n216 );  // ../RTL/core/fpu_utils.v(283)
  or \NM/u232  (\NM/n216 , \NM/n234 , \NM/n251 );  // ../RTL/core/fpu_utils.v(283)
  or \NM/u235  (\NM/n249 , \NM/n268 , \NM/n251 );  // ../RTL/core/fpu_utils.v(289)
  not \NM/u24  (\NM/n24 , M_result2[13]);  // ../RTL/core/fpu_utils.v(223)
  or \NM/u240  (\NM/n286 , \NM/n296 , \NM/n253 );  // ../RTL/core/fpu_utils.v(295)
  not \NM/u241  (\NM/n48 , \NM/n249 );  // ../RTL/core/fpu_utils.v(289)
  or \NM/u243  (\NM/n146 , \NM/n176 , \NM/n242 );  // ../RTL/core/fpu_utils.v(259)
  or \NM/u246  (\NM/n284 , \NM/n304 , \NM/n286 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u247  (\NM/n246 , M_result2[6], M_result2[7]);  // ../RTL/core/fpu_utils.v(283)
  or \NM/u25  (\NM/n332 , \NM/n22 , M_result2[15]);  // ../RTL/core/fpu_utils.v(217)
  not \NM/u252  (\NM/n50 , \NM/n284 );  // ../RTL/core/fpu_utils.v(295)
  or \NM/u253  (\NM/n244 , M_result2[5], \NM/n246 );  // ../RTL/core/fpu_utils.v(283)
  or \NM/u254  (\NM/n234 , \NM/n243 , \NM/n236 );  // ../RTL/core/fpu_utils.v(283)
  not \NM/u255  (\NM/n39 , \NM/n177 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u256  (\NM/n236 , \NM/n276 , \NM/n271 );  // ../RTL/core/fpu_utils.v(283)
  or \NM/u258  (\NM/n281 , M_result2[5], M_result2[6]);  // ../RTL/core/fpu_utils.v(289)
  or \NM/u259  (\NM/n243 , \NM/n248 , \NM/n244 );  // ../RTL/core/fpu_utils.v(283)
  not \NM/u26  (\NM/n26 , M_result2[12]);  // ../RTL/core/fpu_utils.v(229)
  or \NM/u261  (\NM/n177 , \NM/n186 , \NM/n134 );  // ../RTL/core/fpu_utils.v(265)
  or \NM/u264  (\NM/n319 , \NM/n49 , M_result2[2]);  // ../RTL/core/fpu_utils.v(295)
  or \NM/u265  (\NM/n320 , \NM/n260 , \NM/n374 );  // ../RTL/core/fpu_utils.v(253)
  or \NM/u266  (\NM/n315 , \NM/n265 , \NM/n320 );  // ../RTL/core/fpu_utils.v(253)
  or \NM/u267  (\NM/n310 , \NM/n126 , \NM/n315 );  // ../RTL/core/fpu_utils.v(253)
  not \NM/u268  (\NM/n35 , \NM/n310 );  // ../RTL/core/fpu_utils.v(253)
  or \NM/u269  (\NM/n300 , \NM/n32 , \NM/n190 );  // ../RTL/core/fpu_utils.v(247)
  or \NM/u27  (\NM/n322 , \NM/n24 , M_result2[14]);  // ../RTL/core/fpu_utils.v(223)
  or \NM/u273  (\NM/n280 , \NM/n300 , \NM/n127 );  // ../RTL/core/fpu_utils.v(247)
  or \NM/u276  (\NM/n265 , \NM/n125 , \NM/n124 );  // ../RTL/core/fpu_utils.v(247)
  or \NM/u277  (\NM/n260 , M_result2[20], M_result2[21]);  // ../RTL/core/fpu_utils.v(247)
  not \NM/u28  (\NM/n28 , M_result2[11]);  // ../RTL/core/fpu_utils.v(235)
  or \NM/u281  (\NM/n240 , \NM/n280 , \NM/n315 );  // ../RTL/core/fpu_utils.v(247)
  not \NM/u282  (\NM/n33 , \NM/n240 );  // ../RTL/core/fpu_utils.v(247)
  or \NM/u283  (\NM/n230 , \NM/n30 , \NM/n273 );  // ../RTL/core/fpu_utils.v(241)
  or \NM/u286  (\NM/n215 , \NM/n189 , \NM/n185 );  // ../RTL/core/fpu_utils.v(241)
  or \NM/u287  (\NM/n210 , \NM/n230 , \NM/n215 );  // ../RTL/core/fpu_utils.v(241)
  or \NM/u289  (\NM/n175 , M_result2[17], \NM/n124 );  // ../RTL/core/fpu_utils.v(241)
  or \NM/u293  (\NM/n171 , \NM/n175 , \NM/n320 );  // ../RTL/core/fpu_utils.v(241)
  or \NM/u294  (\NM/n170 , \NM/n210 , \NM/n171 );  // ../RTL/core/fpu_utils.v(241)
  not \NM/u295  (\NM/n31 , \NM/n170 );  // ../RTL/core/fpu_utils.v(241)
  or \NM/u296  (\NM/n168 , \NM/n28 , \NM/n129 );  // ../RTL/core/fpu_utils.v(235)
  or \NM/u298  (\NM/n166 , M_result2[14], \NM/n185 );  // ../RTL/core/fpu_utils.v(235)
  or \NM/u299  (\NM/n165 , \NM/n168 , \NM/n166 );  // ../RTL/core/fpu_utils.v(235)
  not \NM/u30  (\NM/n30 , M_result2[10]);  // ../RTL/core/fpu_utils.v(241)
  or \NM/u306  (\NM/n158 , \NM/n165 , \NM/n171 );  // ../RTL/core/fpu_utils.v(235)
  not \NM/u307  (\NM/n29 , \NM/n158 );  // ../RTL/core/fpu_utils.v(235)
  or \NM/u308  (\NM/n156 , \NM/n26 , \NM/n189 );  // ../RTL/core/fpu_utils.v(229)
  or \NM/u311  (\NM/n153 , \NM/n156 , \NM/n263 );  // ../RTL/core/fpu_utils.v(229)
  or \NM/u317  (\NM/n321 , \NM/n153 , \NM/n253 );  // ../RTL/core/fpu_utils.v(229)
  not \NM/u318  (\NM/n27 , \NM/n321 );  // ../RTL/core/fpu_utils.v(229)
  not \NM/u32  (\NM/n32 , M_result2[9]);  // ../RTL/core/fpu_utils.v(247)
  or \NM/u321  (\NM/n325 , \NM/n322 , \NM/n263 );  // ../RTL/core/fpu_utils.v(223)
  or \NM/u327  (\NM/n331 , \NM/n325 , \NM/n253 );  // ../RTL/core/fpu_utils.v(223)
  not \NM/u328  (\NM/n25 , \NM/n331 );  // ../RTL/core/fpu_utils.v(223)
  or \NM/u331  (\NM/n335 , \NM/n332 , \NM/n207 );  // ../RTL/core/fpu_utils.v(217)
  or \NM/u336  (\NM/n340 , \NM/n335 , \NM/n179 );  // ../RTL/core/fpu_utils.v(217)
  not \NM/u337  (\NM/n23 , \NM/n340 );  // ../RTL/core/fpu_utils.v(217)
  or \NM/u339  (\NM/n343 , \NM/n341 , \NM/n184 );  // ../RTL/core/fpu_utils.v(211)
  not \NM/u34  (\NM/n34 , M_result2[8]);  // ../RTL/core/fpu_utils.v(253)
  or \NM/u344  (\NM/n348 , \NM/n343 , \NM/n179 );  // ../RTL/core/fpu_utils.v(211)
  not \NM/u345  (\NM/n21 , \NM/n348 );  // ../RTL/core/fpu_utils.v(211)
  or \NM/u347  (\NM/n351 , \NM/n349 , \NM/n124 );  // ../RTL/core/fpu_utils.v(205)
  or \NM/u351  (\NM/n355 , \NM/n351 , \NM/n320 );  // ../RTL/core/fpu_utils.v(205)
  not \NM/u352  (\NM/n19 , \NM/n355 );  // ../RTL/core/fpu_utils.v(205)
  or \NM/u353  (\NM/n357 , \NM/n16 , \NM/n124 );  // ../RTL/core/fpu_utils.v(199)
  or \NM/u357  (\NM/n361 , \NM/n357 , \NM/n320 );  // ../RTL/core/fpu_utils.v(199)
  not \NM/u358  (\NM/n17 , \NM/n361 );  // ../RTL/core/fpu_utils.v(199)
  or \NM/u359  (\NM/n363 , \NM/n14 , \NM/n182 );  // ../RTL/core/fpu_utils.v(193)
  not \NM/u36  (\NM/n36 , M_result2[7]);  // ../RTL/core/fpu_utils.v(259)
  or \NM/u362  (\NM/n366 , \NM/n363 , \NM/n180 );  // ../RTL/core/fpu_utils.v(193)
  not \NM/u363  (\NM/n15 , \NM/n366 );  // ../RTL/core/fpu_utils.v(193)
  or \NM/u366  (\NM/n370 , \NM/n367 , \NM/n180 );  // ../RTL/core/fpu_utils.v(187)
  not \NM/u367  (\NM/n13 , \NM/n370 );  // ../RTL/core/fpu_utils.v(187)
  or \NM/u369  (\NM/n373 , \NM/n371 , \NM/n374 );  // ../RTL/core/fpu_utils.v(181)
  or \NM/u37  (\NM/n132 , \NM/n34 , M_result2[9]);  // ../RTL/core/fpu_utils.v(253)
  not \NM/u370  (\NM/n11 , \NM/n373 );  // ../RTL/core/fpu_utils.v(181)
  or \NM/u371  (\NM/n375 , \NM/n8 , \NM/n374 );  // ../RTL/core/fpu_utils.v(175)
  not \NM/u372  (\NM/n9 , \NM/n375 );  // ../RTL/core/fpu_utils.v(175)
  not \NM/u373  (\NM/n7 , \NM/n376 );  // ../RTL/core/fpu_utils.v(169)
  not \NM/u38  (\NM/n38 , M_result2[6]);  // ../RTL/core/fpu_utils.v(265)
  or \NM/u39  (\NM/n176 , \NM/n36 , M_result2[8]);  // ../RTL/core/fpu_utils.v(259)
  not \NM/u40  (\NM/n40 , M_result2[5]);  // ../RTL/core/fpu_utils.v(271)
  or \NM/u41  (\NM/n193 , \NM/n38 , M_result2[7]);  // ../RTL/core/fpu_utils.v(265)
  not \NM/u42  (\NM/n42 , M_result2[4]);  // ../RTL/core/fpu_utils.v(277)
  or \NM/u44  (\NM/n257 , \NM/n40 , M_result2[6]);  // ../RTL/core/fpu_utils.v(271)
  not \NM/u45  (\NM/n45 , M_result2[3]);  // ../RTL/core/fpu_utils.v(283)
  or \NM/u46  (\NM/n214 , \NM/n42 , M_result2[5]);  // ../RTL/core/fpu_utils.v(277)
  not \NM/u47  (\NM/n47 , M_result2[2]);  // ../RTL/core/fpu_utils.v(289)
  or \NM/u48  (\NM/n248 , \NM/n45 , M_result2[4]);  // ../RTL/core/fpu_utils.v(283)
  not \NM/u49  (\NM/n49 , M_result2[1]);  // ../RTL/core/fpu_utils.v(295)
  and \NM/u5  (\NM/n2 , M_carry, \M04/M01/M01/invSL );  // ../RTL/core/fpu_utils.v(156)
  or \NM/u50  (\NM/n283 , \NM/n47 , M_result2[3]);  // ../RTL/core/fpu_utils.v(289)
  not \NM/u51  (\NM/n52 , M_result2[23]);  // ../RTL/core/fpu_utils.v(163)
  and \NM/u52  (\NM/n53 , \NM/n7 , \NM/n52 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u53  (\NM/n54 , M_result2[23], \NM/n7 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u54  (\NM/n55 , \NM/n54 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u55  (\NM/n56 , \NM/n9 , \NM/n55 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u56  (\NM/n57 , \NM/n54 , \NM/n9 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u57  (\NM/n58 , \NM/n57 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u58  (\NM/n59 , \NM/n11 , \NM/n58 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u59  (\NM/n60 , \NM/n57 , \NM/n11 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u60  (\NM/n61 , \NM/n60 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u61  (\NM/n62 , \NM/n13 , \NM/n61 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u62  (\NM/n63 , \NM/n60 , \NM/n13 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u63  (\NM/n64 , \NM/n63 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u64  (\NM/n65 , \NM/n15 , \NM/n64 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u65  (\NM/n66 , \NM/n63 , \NM/n15 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u66  (\NM/n67 , \NM/n66 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u67  (\NM/n68 , \NM/n17 , \NM/n67 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u68  (\NM/n69 , \NM/n66 , \NM/n17 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u69  (\NM/n70 , \NM/n69 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u7  (\NM/n6 , M_result2[22]);  // ../RTL/core/fpu_utils.v(169)
  and \NM/u70  (\NM/n71 , \NM/n19 , \NM/n70 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u71  (\NM/n72 , \NM/n69 , \NM/n19 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u72  (\NM/n73 , \NM/n72 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u73  (\NM/n74 , \NM/n21 , \NM/n73 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u74  (\NM/n75 , \NM/n72 , \NM/n21 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u75  (\NM/n76 , \NM/n75 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u76  (\NM/n77 , \NM/n23 , \NM/n76 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u77  (\NM/n78 , \NM/n75 , \NM/n23 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u78  (\NM/n79 , \NM/n78 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u79  (\NM/n80 , \NM/n25 , \NM/n79 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u8  (\NM/n8 , M_result2[21]);  // ../RTL/core/fpu_utils.v(175)
  or \NM/u80  (\NM/n81 , \NM/n78 , \NM/n25 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u81  (\NM/n82 , \NM/n81 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u82  (\NM/n83 , \NM/n27 , \NM/n82 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u83  (\NM/n84 , \NM/n81 , \NM/n27 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u84  (\NM/n85 , \NM/n84 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u85  (\NM/n86 , \NM/n29 , \NM/n85 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u86  (\NM/n87 , \NM/n84 , \NM/n29 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u87  (\NM/n88 , \NM/n87 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u88  (\NM/n89 , \NM/n31 , \NM/n88 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u89  (\NM/n90 , \NM/n87 , \NM/n31 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u9  (\NM/n376 , \NM/n6 , M_result2[23]);  // ../RTL/core/fpu_utils.v(169)
  not \NM/u90  (\NM/n91 , \NM/n90 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u91  (\NM/n92 , \NM/n33 , \NM/n91 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u92  (\NM/n93 , \NM/n90 , \NM/n33 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u93  (\NM/n94 , \NM/n93 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u94  (\NM/n95 , \NM/n35 , \NM/n94 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u95  (\NM/n96 , \NM/n93 , \NM/n35 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u96  (\NM/n97 , \NM/n96 );  // ../RTL/core/fpu_utils.v(163)
  and \NM/u97  (\NM/n98 , \NM/n37 , \NM/n97 );  // ../RTL/core/fpu_utils.v(163)
  or \NM/u98  (\NM/n99 , \NM/n96 , \NM/n37 );  // ../RTL/core/fpu_utils.v(163)
  not \NM/u99  (\NM/n100 , \NM/n99 );  // ../RTL/core/fpu_utils.v(163)
  or \RO01/u0  (\RO01/w1 , n1[24], n1[23]);  // ../RTL/core/fpu_utils.v(14)
  or \RO01/u1  (\RO01/w2 , n1[25], \RO01/w1 );  // ../RTL/core/fpu_utils.v(15)
  or \RO01/u2  (\RO01/w3 , n1[26], \RO01/w2 );  // ../RTL/core/fpu_utils.v(16)
  or \RO01/u3  (\RO01/w4 , n1[27], \RO01/w3 );  // ../RTL/core/fpu_utils.v(17)
  or \RO01/u4  (\RO01/w5 , n1[28], \RO01/w4 );  // ../RTL/core/fpu_utils.v(18)
  or \RO01/u5  (\RO01/w6 , n1[29], \RO01/w5 );  // ../RTL/core/fpu_utils.v(19)
  or \RO01/u6  (reduced_or_E1, n1[30], \RO01/w6 );  // ../RTL/core/fpu_utils.v(20)
  not \exp_diff[4]_inv  (\exp_diff[4]_neg , exp_diff[4]);
  binary_mux_s1_w1 mux0_b0 (
    .i0(n37[0]),
    .i1(n1[0]),
    .sel(isE1GreaterThanE2),
    .o(M1[0]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b1 (
    .i0(n37[1]),
    .i1(n1[1]),
    .sel(isE1GreaterThanE2),
    .o(M1[1]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b10 (
    .i0(n37[10]),
    .i1(n1[10]),
    .sel(isE1GreaterThanE2),
    .o(M1[10]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b11 (
    .i0(n37[11]),
    .i1(n1[11]),
    .sel(isE1GreaterThanE2),
    .o(M1[11]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b12 (
    .i0(n37[12]),
    .i1(n1[12]),
    .sel(isE1GreaterThanE2),
    .o(M1[12]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b13 (
    .i0(n37[13]),
    .i1(n1[13]),
    .sel(isE1GreaterThanE2),
    .o(M1[13]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b14 (
    .i0(n37[14]),
    .i1(n1[14]),
    .sel(isE1GreaterThanE2),
    .o(M1[14]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b15 (
    .i0(n37[15]),
    .i1(n1[15]),
    .sel(isE1GreaterThanE2),
    .o(M1[15]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b16 (
    .i0(n37[16]),
    .i1(n1[16]),
    .sel(isE1GreaterThanE2),
    .o(M1[16]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b17 (
    .i0(n37[17]),
    .i1(n1[17]),
    .sel(isE1GreaterThanE2),
    .o(M1[17]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b18 (
    .i0(n37[18]),
    .i1(n1[18]),
    .sel(isE1GreaterThanE2),
    .o(M1[18]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b19 (
    .i0(n37[19]),
    .i1(n1[19]),
    .sel(isE1GreaterThanE2),
    .o(M1[19]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b2 (
    .i0(n37[2]),
    .i1(n1[2]),
    .sel(isE1GreaterThanE2),
    .o(M1[2]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b20 (
    .i0(n37[20]),
    .i1(n1[20]),
    .sel(isE1GreaterThanE2),
    .o(M1[20]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b21 (
    .i0(n37[21]),
    .i1(n1[21]),
    .sel(isE1GreaterThanE2),
    .o(M1[21]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b22 (
    .i0(n37[22]),
    .i1(n1[22]),
    .sel(isE1GreaterThanE2),
    .o(M1[22]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b23 (
    .i0(n62[23]),
    .i1(reduced_or_E1),
    .sel(isE1GreaterThanE2),
    .o(M1[23]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b3 (
    .i0(n37[3]),
    .i1(n1[3]),
    .sel(isE1GreaterThanE2),
    .o(M1[3]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b4 (
    .i0(n37[4]),
    .i1(n1[4]),
    .sel(isE1GreaterThanE2),
    .o(M1[4]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b5 (
    .i0(n37[5]),
    .i1(n1[5]),
    .sel(isE1GreaterThanE2),
    .o(M1[5]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b6 (
    .i0(n37[6]),
    .i1(n1[6]),
    .sel(isE1GreaterThanE2),
    .o(M1[6]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b7 (
    .i0(n37[7]),
    .i1(n1[7]),
    .sel(isE1GreaterThanE2),
    .o(M1[7]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b8 (
    .i0(n37[8]),
    .i1(n1[8]),
    .sel(isE1GreaterThanE2),
    .o(M1[8]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux0_b9 (
    .i0(n37[9]),
    .i1(n1[9]),
    .sel(isE1GreaterThanE2),
    .o(M1[9]));  // ../RTL/core/fpu.v(127)
  binary_mux_s1_w1 mux1_b0 (
    .i0(n2[0]),
    .i1(n62[0]),
    .sel(isE1GreaterThanE2),
    .o(M2[0]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b1 (
    .i0(n2[1]),
    .i1(n62[1]),
    .sel(isE1GreaterThanE2),
    .o(M2[1]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b10 (
    .i0(n2[10]),
    .i1(n62[10]),
    .sel(isE1GreaterThanE2),
    .o(M2[10]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b11 (
    .i0(n2[11]),
    .i1(n62[11]),
    .sel(isE1GreaterThanE2),
    .o(M2[11]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b12 (
    .i0(n2[12]),
    .i1(n62[12]),
    .sel(isE1GreaterThanE2),
    .o(M2[12]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b13 (
    .i0(n2[13]),
    .i1(n62[13]),
    .sel(isE1GreaterThanE2),
    .o(M2[13]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b14 (
    .i0(n2[14]),
    .i1(n62[14]),
    .sel(isE1GreaterThanE2),
    .o(M2[14]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b15 (
    .i0(n2[15]),
    .i1(n62[15]),
    .sel(isE1GreaterThanE2),
    .o(M2[15]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b16 (
    .i0(n2[16]),
    .i1(n62[16]),
    .sel(isE1GreaterThanE2),
    .o(M2[16]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b17 (
    .i0(n2[17]),
    .i1(n62[17]),
    .sel(isE1GreaterThanE2),
    .o(M2[17]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b18 (
    .i0(n2[18]),
    .i1(n62[18]),
    .sel(isE1GreaterThanE2),
    .o(M2[18]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b19 (
    .i0(n2[19]),
    .i1(n62[19]),
    .sel(isE1GreaterThanE2),
    .o(M2[19]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b2 (
    .i0(n2[2]),
    .i1(n62[2]),
    .sel(isE1GreaterThanE2),
    .o(M2[2]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b20 (
    .i0(n2[20]),
    .i1(n62[20]),
    .sel(isE1GreaterThanE2),
    .o(M2[20]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b21 (
    .i0(n2[21]),
    .i1(n62[21]),
    .sel(isE1GreaterThanE2),
    .o(M2[21]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b22 (
    .i0(n2[22]),
    .i1(n62[22]),
    .sel(isE1GreaterThanE2),
    .o(M2[22]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b23 (
    .i0(reduced_or_E1),
    .i1(n62[23]),
    .sel(isE1GreaterThanE2),
    .o(M2[23]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b3 (
    .i0(n2[3]),
    .i1(n62[3]),
    .sel(isE1GreaterThanE2),
    .o(M2[3]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b4 (
    .i0(n2[4]),
    .i1(n62[4]),
    .sel(isE1GreaterThanE2),
    .o(M2[4]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b5 (
    .i0(n2[5]),
    .i1(n62[5]),
    .sel(isE1GreaterThanE2),
    .o(M2[5]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b6 (
    .i0(n2[6]),
    .i1(n62[6]),
    .sel(isE1GreaterThanE2),
    .o(M2[6]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b7 (
    .i0(n2[7]),
    .i1(n62[7]),
    .sel(isE1GreaterThanE2),
    .o(M2[7]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b8 (
    .i0(n2[8]),
    .i1(n62[8]),
    .sel(isE1GreaterThanE2),
    .o(M2[8]));  // ../RTL/core/fpu.v(128)
  binary_mux_s1_w1 mux1_b9 (
    .i0(n2[9]),
    .i1(n62[9]),
    .sel(isE1GreaterThanE2),
    .o(M2[9]));  // ../RTL/core/fpu.v(128)
  not n110_inv (n110_neg, n110);
  not \n1[31]_inv  (\n1[31]_neg , n1[31]);
  not \new_E[5]_inv  (\new_E[5]_neg , new_E[5]);
  not \new_E[6]_inv  (\new_E[6]_neg , new_E[6]);
  not \new_E[7]_inv  (\new_E[7]_neg , new_E[7]);
  AL_MUX u100 (
    .i0(n229),
    .i1(n227),
    .sel(exp_diff[1]),
    .o(n123));  // ../RTL/core/fpu.v(128)
  AL_MUX u101 (
    .i0(n228),
    .i1(n226),
    .sel(exp_diff[1]),
    .o(n122));  // ../RTL/core/fpu.v(128)
  AL_MUX u102 (
    .i0(n227),
    .i1(n225),
    .sel(exp_diff[1]),
    .o(n121));  // ../RTL/core/fpu.v(128)
  AL_MUX u103 (
    .i0(n226),
    .i1(n224),
    .sel(exp_diff[1]),
    .o(n120));  // ../RTL/core/fpu.v(128)
  AL_MUX u104 (
    .i0(n225),
    .i1(n223),
    .sel(exp_diff[1]),
    .o(n119));  // ../RTL/core/fpu.v(128)
  AL_MUX u105 (
    .i0(n224),
    .i1(n222),
    .sel(exp_diff[1]),
    .o(n118));  // ../RTL/core/fpu.v(128)
  AL_MUX u106 (
    .i0(n223),
    .i1(n221),
    .sel(exp_diff[1]),
    .o(n117));  // ../RTL/core/fpu.v(128)
  AL_MUX u107 (
    .i0(n222),
    .i1(n165),
    .sel(exp_diff[1]),
    .o(n116));  // ../RTL/core/fpu.v(128)
  AL_MUX u108 (
    .i0(n221),
    .i1(n164),
    .sel(exp_diff[1]),
    .o(n115));  // ../RTL/core/fpu.v(128)
  AL_MUX u109 (
    .i0(n165),
    .i1(n86),
    .sel(exp_diff[1]),
    .o(n114));  // ../RTL/core/fpu.v(128)
  AL_MUX u110 (
    .i0(n164),
    .i1(1'b0),
    .sel(exp_diff[1]),
    .o(n113));  // ../RTL/core/fpu.v(128)
  AL_MUX u111 (
    .i0(n86),
    .i1(1'b0),
    .sel(exp_diff[1]),
    .o(n112));  // ../RTL/core/fpu.v(128)
  AL_MUX u112 (
    .i0(n161),
    .i1(n131),
    .sel(exp_diff[2]),
    .o(n111));  // ../RTL/core/fpu.v(128)
  AL_MUX u113 (
    .i0(n134),
    .i1(n130),
    .sel(exp_diff[2]),
    .o(n220));  // ../RTL/core/fpu.v(128)
  AL_MUX u114 (
    .i0(n133),
    .i1(n129),
    .sel(exp_diff[2]),
    .o(n219));  // ../RTL/core/fpu.v(128)
  AL_MUX u115 (
    .i0(n132),
    .i1(n128),
    .sel(exp_diff[2]),
    .o(n218));  // ../RTL/core/fpu.v(128)
  AL_MUX u116 (
    .i0(n131),
    .i1(n127),
    .sel(exp_diff[2]),
    .o(n217));  // ../RTL/core/fpu.v(128)
  AL_MUX u117 (
    .i0(n130),
    .i1(n126),
    .sel(exp_diff[2]),
    .o(n216));  // ../RTL/core/fpu.v(128)
  AL_MUX u118 (
    .i0(n129),
    .i1(n125),
    .sel(exp_diff[2]),
    .o(n215));  // ../RTL/core/fpu.v(128)
  AL_MUX u119 (
    .i0(n128),
    .i1(n124),
    .sel(exp_diff[2]),
    .o(n214));  // ../RTL/core/fpu.v(128)
  and u12 (w2, \M04/M01/M01/invSL , n1[31]);  // ../RTL/core/fpu.v(141)
  AL_MUX u120 (
    .i0(n127),
    .i1(n123),
    .sel(exp_diff[2]),
    .o(n213));  // ../RTL/core/fpu.v(128)
  AL_MUX u121 (
    .i0(n126),
    .i1(n122),
    .sel(exp_diff[2]),
    .o(n212));  // ../RTL/core/fpu.v(128)
  AL_MUX u122 (
    .i0(n125),
    .i1(n121),
    .sel(exp_diff[2]),
    .o(n211));  // ../RTL/core/fpu.v(128)
  AL_MUX u123 (
    .i0(n124),
    .i1(n120),
    .sel(exp_diff[2]),
    .o(n210));  // ../RTL/core/fpu.v(128)
  AL_MUX u124 (
    .i0(n123),
    .i1(n119),
    .sel(exp_diff[2]),
    .o(n209));  // ../RTL/core/fpu.v(128)
  AL_MUX u125 (
    .i0(n122),
    .i1(n118),
    .sel(exp_diff[2]),
    .o(n208));  // ../RTL/core/fpu.v(128)
  AL_MUX u126 (
    .i0(n121),
    .i1(n117),
    .sel(exp_diff[2]),
    .o(n207));  // ../RTL/core/fpu.v(128)
  AL_MUX u127 (
    .i0(n120),
    .i1(n116),
    .sel(exp_diff[2]),
    .o(n206));  // ../RTL/core/fpu.v(128)
  AL_MUX u128 (
    .i0(n119),
    .i1(n115),
    .sel(exp_diff[2]),
    .o(n205));  // ../RTL/core/fpu.v(128)
  AL_MUX u129 (
    .i0(n118),
    .i1(n114),
    .sel(exp_diff[2]),
    .o(n204));  // ../RTL/core/fpu.v(128)
  and u13 (w3, M_carry, n1[31]);  // ../RTL/core/fpu.v(142)
  AL_MUX u130 (
    .i0(n117),
    .i1(n113),
    .sel(exp_diff[2]),
    .o(n203));  // ../RTL/core/fpu.v(128)
  AL_MUX u131 (
    .i0(n116),
    .i1(n112),
    .sel(exp_diff[2]),
    .o(n202));  // ../RTL/core/fpu.v(128)
  AL_MUX u132 (
    .i0(n115),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n201));  // ../RTL/core/fpu.v(128)
  AL_MUX u133 (
    .i0(n114),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n200));  // ../RTL/core/fpu.v(128)
  AL_MUX u134 (
    .i0(n113),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n199));  // ../RTL/core/fpu.v(128)
  AL_MUX u135 (
    .i0(n112),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n198));  // ../RTL/core/fpu.v(128)
  AL_MUX u136 (
    .i0(n111),
    .i1(n213),
    .sel(exp_diff[3]),
    .o(n197));  // ../RTL/core/fpu.v(128)
  AL_MUX u137 (
    .i0(n220),
    .i1(n212),
    .sel(exp_diff[3]),
    .o(n158));  // ../RTL/core/fpu.v(128)
  AL_MUX u138 (
    .i0(n219),
    .i1(n211),
    .sel(exp_diff[3]),
    .o(n157));  // ../RTL/core/fpu.v(128)
  AL_MUX u139 (
    .i0(n218),
    .i1(n210),
    .sel(exp_diff[3]),
    .o(n156));  // ../RTL/core/fpu.v(128)
  and u14 (n243, real_oper, \n1[31]_neg );  // ../RTL/core/fpu.v(140)
  AL_MUX u140 (
    .i0(n217),
    .i1(n209),
    .sel(exp_diff[3]),
    .o(n155));  // ../RTL/core/fpu.v(128)
  AL_MUX u141 (
    .i0(n216),
    .i1(n208),
    .sel(exp_diff[3]),
    .o(n154));  // ../RTL/core/fpu.v(128)
  AL_MUX u142 (
    .i0(n215),
    .i1(n207),
    .sel(exp_diff[3]),
    .o(n153));  // ../RTL/core/fpu.v(128)
  AL_MUX u143 (
    .i0(n214),
    .i1(n206),
    .sel(exp_diff[3]),
    .o(n152));  // ../RTL/core/fpu.v(128)
  AL_MUX u144 (
    .i0(n213),
    .i1(n205),
    .sel(exp_diff[3]),
    .o(n151));  // ../RTL/core/fpu.v(128)
  AL_MUX u145 (
    .i0(n212),
    .i1(n204),
    .sel(exp_diff[3]),
    .o(n150));  // ../RTL/core/fpu.v(128)
  AL_MUX u146 (
    .i0(n211),
    .i1(n203),
    .sel(exp_diff[3]),
    .o(n149));  // ../RTL/core/fpu.v(128)
  AL_MUX u147 (
    .i0(n210),
    .i1(n202),
    .sel(exp_diff[3]),
    .o(n148));  // ../RTL/core/fpu.v(128)
  AL_MUX u148 (
    .i0(n209),
    .i1(n201),
    .sel(exp_diff[3]),
    .o(n147));  // ../RTL/core/fpu.v(128)
  AL_MUX u149 (
    .i0(n208),
    .i1(n200),
    .sel(exp_diff[3]),
    .o(n146));  // ../RTL/core/fpu.v(128)
  AL_MUX u150 (
    .i0(n207),
    .i1(n199),
    .sel(exp_diff[3]),
    .o(n145));  // ../RTL/core/fpu.v(128)
  AL_MUX u151 (
    .i0(n206),
    .i1(n198),
    .sel(exp_diff[3]),
    .o(n144));  // ../RTL/core/fpu.v(128)
  AL_MUX u152 (
    .i0(n205),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n143));  // ../RTL/core/fpu.v(128)
  AL_MUX u153 (
    .i0(n204),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n142));  // ../RTL/core/fpu.v(128)
  AL_MUX u154 (
    .i0(n203),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n141));  // ../RTL/core/fpu.v(128)
  AL_MUX u155 (
    .i0(n202),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n140));  // ../RTL/core/fpu.v(128)
  AL_MUX u156 (
    .i0(n201),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n139));  // ../RTL/core/fpu.v(128)
  AL_MUX u157 (
    .i0(n200),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n138));  // ../RTL/core/fpu.v(128)
  AL_MUX u158 (
    .i0(n199),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n137));  // ../RTL/core/fpu.v(128)
  AL_MUX u159 (
    .i0(n198),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n136));  // ../RTL/core/fpu.v(128)
  AL_MUX u160 (
    .i0(n197),
    .i1(n143),
    .sel(exp_diff[4]),
    .o(n135));  // ../RTL/core/fpu.v(128)
  AL_MUX u161 (
    .i0(n158),
    .i1(n142),
    .sel(exp_diff[4]),
    .o(n194));  // ../RTL/core/fpu.v(128)
  AL_MUX u162 (
    .i0(n157),
    .i1(n141),
    .sel(exp_diff[4]),
    .o(n193));  // ../RTL/core/fpu.v(128)
  AL_MUX u163 (
    .i0(n156),
    .i1(n140),
    .sel(exp_diff[4]),
    .o(n192));  // ../RTL/core/fpu.v(128)
  AL_MUX u164 (
    .i0(n155),
    .i1(n139),
    .sel(exp_diff[4]),
    .o(n191));  // ../RTL/core/fpu.v(128)
  AL_MUX u165 (
    .i0(n154),
    .i1(n138),
    .sel(exp_diff[4]),
    .o(n190));  // ../RTL/core/fpu.v(128)
  AL_MUX u166 (
    .i0(n153),
    .i1(n137),
    .sel(exp_diff[4]),
    .o(n189));  // ../RTL/core/fpu.v(128)
  AL_MUX u167 (
    .i0(n152),
    .i1(n136),
    .sel(exp_diff[4]),
    .o(n188));  // ../RTL/core/fpu.v(128)
  and u18 (n196, real_oper, n160);  // ../RTL/core/fpu.v(151)
  or u184 (n171, exp_diff[6], exp_diff[7]);  // ../RTL/core/fpu.v(128)
  or u185 (n110, exp_diff[5], n171);  // ../RTL/core/fpu.v(128)
  AL_MUX u186 (
    .i0(n135),
    .i1(1'b0),
    .sel(n110),
    .o(n62[0]));  // ../RTL/core/fpu.v(128)
  AL_MUX u187 (
    .i0(n194),
    .i1(1'b0),
    .sel(n110),
    .o(n62[1]));  // ../RTL/core/fpu.v(128)
  AL_MUX u188 (
    .i0(n193),
    .i1(1'b0),
    .sel(n110),
    .o(n62[2]));  // ../RTL/core/fpu.v(128)
  AL_MUX u189 (
    .i0(n192),
    .i1(1'b0),
    .sel(n110),
    .o(n62[3]));  // ../RTL/core/fpu.v(128)
  or u19 (n244, w2, w1);  // ../RTL/core/fpu.v(143)
  AL_MUX u190 (
    .i0(n191),
    .i1(1'b0),
    .sel(n110),
    .o(n62[4]));  // ../RTL/core/fpu.v(128)
  AL_MUX u191 (
    .i0(n190),
    .i1(1'b0),
    .sel(n110),
    .o(n62[5]));  // ../RTL/core/fpu.v(128)
  AL_MUX u192 (
    .i0(n189),
    .i1(1'b0),
    .sel(n110),
    .o(n62[6]));  // ../RTL/core/fpu.v(128)
  AL_MUX u193 (
    .i0(n188),
    .i1(1'b0),
    .sel(n110),
    .o(n62[7]));  // ../RTL/core/fpu.v(128)
  AL_MUX u194 (
    .i0(1'b0),
    .i1(n151),
    .sel(u194_sel_is_0_o),
    .o(n62[8]));
  and u194_sel_is_0 (u194_sel_is_0_o, n110_neg, \exp_diff[4]_neg );
  AL_MUX u195 (
    .i0(1'b0),
    .i1(n150),
    .sel(u194_sel_is_0_o),
    .o(n62[9]));
  AL_MUX u196 (
    .i0(1'b0),
    .i1(n149),
    .sel(u194_sel_is_0_o),
    .o(n62[10]));
  AL_MUX u197 (
    .i0(1'b0),
    .i1(n148),
    .sel(u194_sel_is_0_o),
    .o(n62[11]));
  AL_MUX u198 (
    .i0(1'b0),
    .i1(n147),
    .sel(u194_sel_is_0_o),
    .o(n62[12]));
  AL_MUX u199 (
    .i0(1'b0),
    .i1(n146),
    .sel(u194_sel_is_0_o),
    .o(n62[13]));
  AL_MUX u200 (
    .i0(1'b0),
    .i1(n145),
    .sel(u194_sel_is_0_o),
    .o(n62[14]));
  AL_MUX u201 (
    .i0(1'b0),
    .i1(n144),
    .sel(u194_sel_is_0_o),
    .o(n62[15]));
  AL_MUX u202 (
    .i0(1'b0),
    .i1(n143),
    .sel(u194_sel_is_0_o),
    .o(n62[16]));
  AL_MUX u203 (
    .i0(1'b0),
    .i1(n142),
    .sel(u194_sel_is_0_o),
    .o(n62[17]));
  AL_MUX u204 (
    .i0(1'b0),
    .i1(n141),
    .sel(u194_sel_is_0_o),
    .o(n62[18]));
  AL_MUX u205 (
    .i0(1'b0),
    .i1(n140),
    .sel(u194_sel_is_0_o),
    .o(n62[19]));
  AL_MUX u206 (
    .i0(1'b0),
    .i1(n139),
    .sel(u194_sel_is_0_o),
    .o(n62[20]));
  AL_MUX u207 (
    .i0(1'b0),
    .i1(n138),
    .sel(u194_sel_is_0_o),
    .o(n62[21]));
  AL_MUX u208 (
    .i0(1'b0),
    .i1(n137),
    .sel(u194_sel_is_0_o),
    .o(n62[22]));
  AL_MUX u209 (
    .i0(1'b0),
    .i1(n136),
    .sel(u194_sel_is_0_o),
    .o(n62[23]));
  AL_MUX u210 (
    .i0(n1[1]),
    .i1(n1[2]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n108));  // ../RTL/core/fpu.v(127)
  AL_MUX u211 (
    .i0(n1[2]),
    .i1(n1[3]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n107));  // ../RTL/core/fpu.v(127)
  AL_MUX u212 (
    .i0(n1[3]),
    .i1(n1[4]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n106));  // ../RTL/core/fpu.v(127)
  AL_MUX u213 (
    .i0(n1[4]),
    .i1(n1[5]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n105));  // ../RTL/core/fpu.v(127)
  AL_MUX u214 (
    .i0(n1[5]),
    .i1(n1[6]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n104));  // ../RTL/core/fpu.v(127)
  AL_MUX u215 (
    .i0(n1[6]),
    .i1(n1[7]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n103));  // ../RTL/core/fpu.v(127)
  AL_MUX u216 (
    .i0(n1[7]),
    .i1(n1[8]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n102));  // ../RTL/core/fpu.v(127)
  AL_MUX u217 (
    .i0(n1[8]),
    .i1(n1[9]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n101));  // ../RTL/core/fpu.v(127)
  AL_MUX u218 (
    .i0(n1[9]),
    .i1(n1[10]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n100));  // ../RTL/core/fpu.v(127)
  AL_MUX u219 (
    .i0(n1[10]),
    .i1(n1[11]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n99));  // ../RTL/core/fpu.v(127)
  AL_MUX u220 (
    .i0(n1[11]),
    .i1(n1[12]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n98));  // ../RTL/core/fpu.v(127)
  AL_MUX u221 (
    .i0(n1[12]),
    .i1(n1[13]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n97));  // ../RTL/core/fpu.v(127)
  AL_MUX u222 (
    .i0(n1[13]),
    .i1(n1[14]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n96));  // ../RTL/core/fpu.v(127)
  AL_MUX u223 (
    .i0(n1[14]),
    .i1(n1[15]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n95));  // ../RTL/core/fpu.v(127)
  AL_MUX u224 (
    .i0(n1[15]),
    .i1(n1[16]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n94));  // ../RTL/core/fpu.v(127)
  AL_MUX u225 (
    .i0(n1[16]),
    .i1(n1[17]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n93));  // ../RTL/core/fpu.v(127)
  AL_MUX u226 (
    .i0(n1[17]),
    .i1(n1[18]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n92));  // ../RTL/core/fpu.v(127)
  AL_MUX u227 (
    .i0(n1[18]),
    .i1(n1[19]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n91));  // ../RTL/core/fpu.v(127)
  AL_MUX u228 (
    .i0(n1[19]),
    .i1(n1[20]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n90));  // ../RTL/core/fpu.v(127)
  AL_MUX u229 (
    .i0(n1[20]),
    .i1(n1[21]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n89));  // ../RTL/core/fpu.v(127)
  AL_MUX u230 (
    .i0(n1[21]),
    .i1(n1[22]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n88));  // ../RTL/core/fpu.v(127)
  AL_MUX u231 (
    .i0(n1[22]),
    .i1(reduced_or_E1),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n87));  // ../RTL/core/fpu.v(127)
  AL_MUX u232 (
    .i0(reduced_or_E1),
    .i1(1'b0),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n86));  // ../RTL/core/fpu.v(127)
  AL_MUX u233 (
    .i0(n109),
    .i1(n107),
    .sel(exp_diff[1]),
    .o(n85));  // ../RTL/core/fpu.v(127)
  AL_MUX u234 (
    .i0(n108),
    .i1(n106),
    .sel(exp_diff[1]),
    .o(n84));  // ../RTL/core/fpu.v(127)
  AL_MUX u235 (
    .i0(n107),
    .i1(n105),
    .sel(exp_diff[1]),
    .o(n83));  // ../RTL/core/fpu.v(127)
  AL_MUX u236 (
    .i0(n106),
    .i1(n104),
    .sel(exp_diff[1]),
    .o(n82));  // ../RTL/core/fpu.v(127)
  AL_MUX u237 (
    .i0(n105),
    .i1(n103),
    .sel(exp_diff[1]),
    .o(n81));  // ../RTL/core/fpu.v(127)
  AL_MUX u238 (
    .i0(n104),
    .i1(n102),
    .sel(exp_diff[1]),
    .o(n80));  // ../RTL/core/fpu.v(127)
  AL_MUX u239 (
    .i0(n103),
    .i1(n101),
    .sel(exp_diff[1]),
    .o(n79));  // ../RTL/core/fpu.v(127)
  AL_MUX u240 (
    .i0(n102),
    .i1(n100),
    .sel(exp_diff[1]),
    .o(n78));  // ../RTL/core/fpu.v(127)
  AL_MUX u241 (
    .i0(n101),
    .i1(n99),
    .sel(exp_diff[1]),
    .o(n77));  // ../RTL/core/fpu.v(127)
  AL_MUX u242 (
    .i0(n100),
    .i1(n98),
    .sel(exp_diff[1]),
    .o(n76));  // ../RTL/core/fpu.v(127)
  AL_MUX u243 (
    .i0(n99),
    .i1(n97),
    .sel(exp_diff[1]),
    .o(n75));  // ../RTL/core/fpu.v(127)
  AL_MUX u244 (
    .i0(n98),
    .i1(n96),
    .sel(exp_diff[1]),
    .o(n74));  // ../RTL/core/fpu.v(127)
  AL_MUX u245 (
    .i0(n97),
    .i1(n95),
    .sel(exp_diff[1]),
    .o(n73));  // ../RTL/core/fpu.v(127)
  AL_MUX u246 (
    .i0(n96),
    .i1(n94),
    .sel(exp_diff[1]),
    .o(n72));  // ../RTL/core/fpu.v(127)
  AL_MUX u247 (
    .i0(n95),
    .i1(n93),
    .sel(exp_diff[1]),
    .o(n71));  // ../RTL/core/fpu.v(127)
  AL_MUX u248 (
    .i0(n94),
    .i1(n92),
    .sel(exp_diff[1]),
    .o(n70));  // ../RTL/core/fpu.v(127)
  AL_MUX u249 (
    .i0(n93),
    .i1(n91),
    .sel(exp_diff[1]),
    .o(n69));  // ../RTL/core/fpu.v(127)
  AL_MUX u250 (
    .i0(n92),
    .i1(n90),
    .sel(exp_diff[1]),
    .o(n68));  // ../RTL/core/fpu.v(127)
  AL_MUX u251 (
    .i0(n91),
    .i1(n89),
    .sel(exp_diff[1]),
    .o(n67));  // ../RTL/core/fpu.v(127)
  AL_MUX u252 (
    .i0(n90),
    .i1(n88),
    .sel(exp_diff[1]),
    .o(n66));  // ../RTL/core/fpu.v(127)
  AL_MUX u253 (
    .i0(n89),
    .i1(n87),
    .sel(exp_diff[1]),
    .o(n65));  // ../RTL/core/fpu.v(127)
  AL_MUX u254 (
    .i0(n88),
    .i1(n86),
    .sel(exp_diff[1]),
    .o(n64));  // ../RTL/core/fpu.v(127)
  AL_MUX u255 (
    .i0(n87),
    .i1(1'b0),
    .sel(exp_diff[1]),
    .o(n63));  // ../RTL/core/fpu.v(127)
  AL_MUX u257 (
    .i0(n85),
    .i1(n81),
    .sel(exp_diff[2]),
    .o(n60));  // ../RTL/core/fpu.v(127)
  AL_MUX u258 (
    .i0(n84),
    .i1(n80),
    .sel(exp_diff[2]),
    .o(n59));  // ../RTL/core/fpu.v(127)
  AL_MUX u259 (
    .i0(n83),
    .i1(n79),
    .sel(exp_diff[2]),
    .o(n58));  // ../RTL/core/fpu.v(127)
  AL_MUX u260 (
    .i0(n82),
    .i1(n78),
    .sel(exp_diff[2]),
    .o(n57));  // ../RTL/core/fpu.v(127)
  AL_MUX u261 (
    .i0(n81),
    .i1(n77),
    .sel(exp_diff[2]),
    .o(n56));  // ../RTL/core/fpu.v(127)
  AL_MUX u262 (
    .i0(n80),
    .i1(n76),
    .sel(exp_diff[2]),
    .o(n55));  // ../RTL/core/fpu.v(127)
  AL_MUX u263 (
    .i0(n79),
    .i1(n75),
    .sel(exp_diff[2]),
    .o(n54));  // ../RTL/core/fpu.v(127)
  AL_MUX u264 (
    .i0(n78),
    .i1(n74),
    .sel(exp_diff[2]),
    .o(n53));  // ../RTL/core/fpu.v(127)
  AL_MUX u265 (
    .i0(n77),
    .i1(n73),
    .sel(exp_diff[2]),
    .o(n52));  // ../RTL/core/fpu.v(127)
  AL_MUX u266 (
    .i0(n76),
    .i1(n72),
    .sel(exp_diff[2]),
    .o(n51));  // ../RTL/core/fpu.v(127)
  AL_MUX u267 (
    .i0(n75),
    .i1(n71),
    .sel(exp_diff[2]),
    .o(n50));  // ../RTL/core/fpu.v(127)
  AL_MUX u268 (
    .i0(n74),
    .i1(n70),
    .sel(exp_diff[2]),
    .o(n49));  // ../RTL/core/fpu.v(127)
  AL_MUX u269 (
    .i0(n73),
    .i1(n69),
    .sel(exp_diff[2]),
    .o(n48));  // ../RTL/core/fpu.v(127)
  AL_MUX u270 (
    .i0(n72),
    .i1(n68),
    .sel(exp_diff[2]),
    .o(n47));  // ../RTL/core/fpu.v(127)
  AL_MUX u271 (
    .i0(n71),
    .i1(n67),
    .sel(exp_diff[2]),
    .o(n46));  // ../RTL/core/fpu.v(127)
  AL_MUX u272 (
    .i0(n70),
    .i1(n66),
    .sel(exp_diff[2]),
    .o(n45));  // ../RTL/core/fpu.v(127)
  AL_MUX u273 (
    .i0(n69),
    .i1(n65),
    .sel(exp_diff[2]),
    .o(n44));  // ../RTL/core/fpu.v(127)
  AL_MUX u274 (
    .i0(n68),
    .i1(n64),
    .sel(exp_diff[2]),
    .o(n43));  // ../RTL/core/fpu.v(127)
  AL_MUX u275 (
    .i0(n67),
    .i1(n63),
    .sel(exp_diff[2]),
    .o(n42));  // ../RTL/core/fpu.v(127)
  AL_MUX u276 (
    .i0(n66),
    .i1(n112),
    .sel(exp_diff[2]),
    .o(n41));  // ../RTL/core/fpu.v(127)
  AL_MUX u277 (
    .i0(n65),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n40));  // ../RTL/core/fpu.v(127)
  AL_MUX u278 (
    .i0(n64),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n39));  // ../RTL/core/fpu.v(127)
  AL_MUX u279 (
    .i0(n63),
    .i1(1'b0),
    .sel(exp_diff[2]),
    .o(n38));  // ../RTL/core/fpu.v(127)
  AL_MUX u281 (
    .i0(n60),
    .i1(n52),
    .sel(exp_diff[3]),
    .o(n263));  // ../RTL/core/fpu.v(127)
  AL_MUX u282 (
    .i0(n59),
    .i1(n51),
    .sel(exp_diff[3]),
    .o(n262));  // ../RTL/core/fpu.v(127)
  AL_MUX u283 (
    .i0(n58),
    .i1(n50),
    .sel(exp_diff[3]),
    .o(n261));  // ../RTL/core/fpu.v(127)
  AL_MUX u284 (
    .i0(n57),
    .i1(n49),
    .sel(exp_diff[3]),
    .o(n260));  // ../RTL/core/fpu.v(127)
  AL_MUX u285 (
    .i0(n56),
    .i1(n48),
    .sel(exp_diff[3]),
    .o(n259));  // ../RTL/core/fpu.v(127)
  AL_MUX u286 (
    .i0(n55),
    .i1(n47),
    .sel(exp_diff[3]),
    .o(n258));  // ../RTL/core/fpu.v(127)
  AL_MUX u287 (
    .i0(n54),
    .i1(n46),
    .sel(exp_diff[3]),
    .o(n257));  // ../RTL/core/fpu.v(127)
  AL_MUX u288 (
    .i0(n53),
    .i1(n45),
    .sel(exp_diff[3]),
    .o(n265));  // ../RTL/core/fpu.v(127)
  AL_MUX u289 (
    .i0(n52),
    .i1(n44),
    .sel(exp_diff[3]),
    .o(n256));  // ../RTL/core/fpu.v(127)
  AL_MUX u290 (
    .i0(n51),
    .i1(n43),
    .sel(exp_diff[3]),
    .o(n255));  // ../RTL/core/fpu.v(127)
  AL_MUX u291 (
    .i0(n50),
    .i1(n42),
    .sel(exp_diff[3]),
    .o(n254));  // ../RTL/core/fpu.v(127)
  AL_MUX u292 (
    .i0(n49),
    .i1(n41),
    .sel(exp_diff[3]),
    .o(n253));  // ../RTL/core/fpu.v(127)
  AL_MUX u293 (
    .i0(n48),
    .i1(n40),
    .sel(exp_diff[3]),
    .o(n252));  // ../RTL/core/fpu.v(127)
  AL_MUX u294 (
    .i0(n47),
    .i1(n39),
    .sel(exp_diff[3]),
    .o(n251));  // ../RTL/core/fpu.v(127)
  AL_MUX u295 (
    .i0(n46),
    .i1(n38),
    .sel(exp_diff[3]),
    .o(n250));  // ../RTL/core/fpu.v(127)
  AL_MUX u296 (
    .i0(n45),
    .i1(n198),
    .sel(exp_diff[3]),
    .o(n249));  // ../RTL/core/fpu.v(127)
  AL_MUX u297 (
    .i0(n44),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n11));  // ../RTL/core/fpu.v(127)
  AL_MUX u298 (
    .i0(n43),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n10));  // ../RTL/core/fpu.v(127)
  AL_MUX u299 (
    .i0(n42),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n9));  // ../RTL/core/fpu.v(127)
  AL_MUX u300 (
    .i0(n41),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n8));  // ../RTL/core/fpu.v(127)
  AL_MUX u301 (
    .i0(n40),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n7));  // ../RTL/core/fpu.v(127)
  AL_MUX u302 (
    .i0(n39),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n6));  // ../RTL/core/fpu.v(127)
  AL_MUX u303 (
    .i0(n38),
    .i1(1'b0),
    .sel(exp_diff[3]),
    .o(n5));  // ../RTL/core/fpu.v(127)
  AL_MUX u305 (
    .i0(n263),
    .i1(n11),
    .sel(exp_diff[4]),
    .o(n36));  // ../RTL/core/fpu.v(127)
  AL_MUX u306 (
    .i0(n262),
    .i1(n10),
    .sel(exp_diff[4]),
    .o(n35));  // ../RTL/core/fpu.v(127)
  AL_MUX u307 (
    .i0(n261),
    .i1(n9),
    .sel(exp_diff[4]),
    .o(n34));  // ../RTL/core/fpu.v(127)
  AL_MUX u308 (
    .i0(n260),
    .i1(n8),
    .sel(exp_diff[4]),
    .o(n33));  // ../RTL/core/fpu.v(127)
  AL_MUX u309 (
    .i0(n259),
    .i1(n7),
    .sel(exp_diff[4]),
    .o(n32));  // ../RTL/core/fpu.v(127)
  AL_MUX u310 (
    .i0(n258),
    .i1(n6),
    .sel(exp_diff[4]),
    .o(n31));  // ../RTL/core/fpu.v(127)
  AL_MUX u311 (
    .i0(n257),
    .i1(n5),
    .sel(exp_diff[4]),
    .o(n30));  // ../RTL/core/fpu.v(127)
  AL_MUX u312 (
    .i0(n265),
    .i1(n136),
    .sel(exp_diff[4]),
    .o(n29));  // ../RTL/core/fpu.v(127)
  AL_MUX u331 (
    .i0(n36),
    .i1(1'b0),
    .sel(n110),
    .o(n37[0]));  // ../RTL/core/fpu.v(127)
  AL_MUX u332 (
    .i0(n35),
    .i1(1'b0),
    .sel(n110),
    .o(n37[1]));  // ../RTL/core/fpu.v(127)
  AL_MUX u333 (
    .i0(n34),
    .i1(1'b0),
    .sel(n110),
    .o(n37[2]));  // ../RTL/core/fpu.v(127)
  AL_MUX u334 (
    .i0(n33),
    .i1(1'b0),
    .sel(n110),
    .o(n37[3]));  // ../RTL/core/fpu.v(127)
  AL_MUX u335 (
    .i0(n32),
    .i1(1'b0),
    .sel(n110),
    .o(n37[4]));  // ../RTL/core/fpu.v(127)
  AL_MUX u336 (
    .i0(n31),
    .i1(1'b0),
    .sel(n110),
    .o(n37[5]));  // ../RTL/core/fpu.v(127)
  AL_MUX u337 (
    .i0(n30),
    .i1(1'b0),
    .sel(n110),
    .o(n37[6]));  // ../RTL/core/fpu.v(127)
  AL_MUX u338 (
    .i0(n29),
    .i1(1'b0),
    .sel(n110),
    .o(n37[7]));  // ../RTL/core/fpu.v(127)
  AL_MUX u339 (
    .i0(1'b0),
    .i1(n256),
    .sel(u194_sel_is_0_o),
    .o(n37[8]));
  AL_MUX u340 (
    .i0(1'b0),
    .i1(n255),
    .sel(u194_sel_is_0_o),
    .o(n37[9]));
  AL_MUX u341 (
    .i0(1'b0),
    .i1(n254),
    .sel(u194_sel_is_0_o),
    .o(n37[10]));
  AL_MUX u342 (
    .i0(1'b0),
    .i1(n253),
    .sel(u194_sel_is_0_o),
    .o(n37[11]));
  AL_MUX u343 (
    .i0(1'b0),
    .i1(n252),
    .sel(u194_sel_is_0_o),
    .o(n37[12]));
  AL_MUX u344 (
    .i0(1'b0),
    .i1(n251),
    .sel(u194_sel_is_0_o),
    .o(n37[13]));
  AL_MUX u345 (
    .i0(1'b0),
    .i1(n250),
    .sel(u194_sel_is_0_o),
    .o(n37[14]));
  AL_MUX u346 (
    .i0(1'b0),
    .i1(n249),
    .sel(u194_sel_is_0_o),
    .o(n37[15]));
  AL_MUX u347 (
    .i0(1'b0),
    .i1(n11),
    .sel(u194_sel_is_0_o),
    .o(n37[16]));
  AL_MUX u348 (
    .i0(1'b0),
    .i1(n10),
    .sel(u194_sel_is_0_o),
    .o(n37[17]));
  AL_MUX u349 (
    .i0(1'b0),
    .i1(n9),
    .sel(u194_sel_is_0_o),
    .o(n37[18]));
  AL_MUX u350 (
    .i0(1'b0),
    .i1(n8),
    .sel(u194_sel_is_0_o),
    .o(n37[19]));
  AL_MUX u351 (
    .i0(1'b0),
    .i1(n7),
    .sel(u194_sel_is_0_o),
    .o(n37[20]));
  AL_MUX u352 (
    .i0(1'b0),
    .i1(n6),
    .sel(u194_sel_is_0_o),
    .o(n37[21]));
  AL_MUX u353 (
    .i0(1'b0),
    .i1(n5),
    .sel(u194_sel_is_0_o),
    .o(n37[22]));
  AL_MUX u5 (
    .i0(n1[0]),
    .i1(n1[1]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n109));  // ../RTL/core/fpu.v(127)
  AL_MUX u6 (
    .i0(n2[0]),
    .i1(n2[1]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n241));  // ../RTL/core/fpu.v(128)
  or u62 (result[31], w3, n244);  // ../RTL/core/fpu.v(143)
  and u63 (w1, n160, n243);  // ../RTL/core/fpu.v(140)
  xor u64 (real_oper, n2[31], \n1[31]_neg );  // ../RTL/core/fpu.v(131)
  AL_MUX u65 (
    .i0(n2[1]),
    .i1(n2[2]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n240));  // ../RTL/core/fpu.v(128)
  AL_MUX u66 (
    .i0(n2[2]),
    .i1(n2[3]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n239));  // ../RTL/core/fpu.v(128)
  AL_MUX u67 (
    .i0(n2[3]),
    .i1(n2[4]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n238));  // ../RTL/core/fpu.v(128)
  AL_MUX u68 (
    .i0(n2[4]),
    .i1(n2[5]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n237));  // ../RTL/core/fpu.v(128)
  AL_MUX u69 (
    .i0(n2[5]),
    .i1(n2[6]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n236));  // ../RTL/core/fpu.v(128)
  AL_MUX u70 (
    .i0(n2[6]),
    .i1(n2[7]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n235));  // ../RTL/core/fpu.v(128)
  AL_MUX u71 (
    .i0(n2[7]),
    .i1(n2[8]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n234));  // ../RTL/core/fpu.v(128)
  AL_MUX u72 (
    .i0(n2[8]),
    .i1(n2[9]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n233));  // ../RTL/core/fpu.v(128)
  AL_MUX u73 (
    .i0(n2[9]),
    .i1(n2[10]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n232));  // ../RTL/core/fpu.v(128)
  AL_MUX u74 (
    .i0(n2[10]),
    .i1(n2[11]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n231));  // ../RTL/core/fpu.v(128)
  AL_MUX u75 (
    .i0(n2[11]),
    .i1(n2[12]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n230));  // ../RTL/core/fpu.v(128)
  AL_MUX u76 (
    .i0(n2[12]),
    .i1(n2[13]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n229));  // ../RTL/core/fpu.v(128)
  AL_MUX u77 (
    .i0(n2[13]),
    .i1(n2[14]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n228));  // ../RTL/core/fpu.v(128)
  AL_MUX u78 (
    .i0(n2[14]),
    .i1(n2[15]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n227));  // ../RTL/core/fpu.v(128)
  AL_MUX u79 (
    .i0(n2[15]),
    .i1(n2[16]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n226));  // ../RTL/core/fpu.v(128)
  AL_MUX u80 (
    .i0(n2[16]),
    .i1(n2[17]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n225));  // ../RTL/core/fpu.v(128)
  AL_MUX u81 (
    .i0(n2[17]),
    .i1(n2[18]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n224));  // ../RTL/core/fpu.v(128)
  AL_MUX u82 (
    .i0(n2[18]),
    .i1(n2[19]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n223));  // ../RTL/core/fpu.v(128)
  AL_MUX u83 (
    .i0(n2[19]),
    .i1(n2[20]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n222));  // ../RTL/core/fpu.v(128)
  AL_MUX u84 (
    .i0(n2[20]),
    .i1(n2[21]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n221));  // ../RTL/core/fpu.v(128)
  AL_MUX u85 (
    .i0(n2[21]),
    .i1(n2[22]),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n165));  // ../RTL/core/fpu.v(128)
  AL_MUX u86 (
    .i0(n2[22]),
    .i1(reduced_or_E1),
    .sel(\ADD01/ADD01/p0_neg ),
    .o(n164));  // ../RTL/core/fpu.v(128)
  AL_MUX u88 (
    .i0(n241),
    .i1(n239),
    .sel(exp_diff[1]),
    .o(n161));  // ../RTL/core/fpu.v(128)
  AL_MUX u89 (
    .i0(n240),
    .i1(n238),
    .sel(exp_diff[1]),
    .o(n134));  // ../RTL/core/fpu.v(128)
  not u9 (n160, M_carry);  // ../RTL/core/fpu.v(140)
  AL_MUX u90 (
    .i0(n239),
    .i1(n237),
    .sel(exp_diff[1]),
    .o(n133));  // ../RTL/core/fpu.v(128)
  AL_MUX u91 (
    .i0(n238),
    .i1(n236),
    .sel(exp_diff[1]),
    .o(n132));  // ../RTL/core/fpu.v(128)
  AL_MUX u92 (
    .i0(n237),
    .i1(n235),
    .sel(exp_diff[1]),
    .o(n131));  // ../RTL/core/fpu.v(128)
  AL_MUX u93 (
    .i0(n236),
    .i1(n234),
    .sel(exp_diff[1]),
    .o(n130));  // ../RTL/core/fpu.v(128)
  AL_MUX u94 (
    .i0(n235),
    .i1(n233),
    .sel(exp_diff[1]),
    .o(n129));  // ../RTL/core/fpu.v(128)
  AL_MUX u95 (
    .i0(n234),
    .i1(n232),
    .sel(exp_diff[1]),
    .o(n128));  // ../RTL/core/fpu.v(128)
  AL_MUX u96 (
    .i0(n233),
    .i1(n231),
    .sel(exp_diff[1]),
    .o(n127));  // ../RTL/core/fpu.v(128)
  AL_MUX u97 (
    .i0(n232),
    .i1(n230),
    .sel(exp_diff[1]),
    .o(n126));  // ../RTL/core/fpu.v(128)
  AL_MUX u98 (
    .i0(n231),
    .i1(n229),
    .sel(exp_diff[1]),
    .o(n125));  // ../RTL/core/fpu.v(128)
  AL_MUX u99 (
    .i0(n230),
    .i1(n228),
    .sel(exp_diff[1]),
    .o(n124));  // ../RTL/core/fpu.v(128)

endmodule 

module add_pu8_pu8_o8
  (
  i0,
  i1,
  o
  );

  input [7:0] i0;
  input [7:0] i1;
  output [7:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a2;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_b0;
  wire net_b1;
  wire net_b2;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_cout0;
  wire net_cout1;
  wire net_cout2;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_sum0;
  wire net_sum1;
  wire net_sum2;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;

  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));

endmodule 

module mult_s32_s32_o64
  (
  i0,
  i1,
  o
  );

  input signed [31:0] i0;
  input signed [31:0] i1;
  output [63:0] o;

  wire [31:0] and_0;
  wire [31:0] and_1;
  wire [31:0] and_10;
  wire [31:0] and_11;
  wire [31:0] and_12;
  wire [31:0] and_13;
  wire [31:0] and_14;
  wire [31:0] and_15;
  wire [31:0] and_16;
  wire [31:0] and_17;
  wire [31:0] and_18;
  wire [31:0] and_19;
  wire [31:0] and_2;
  wire [31:0] and_20;
  wire [31:0] and_21;
  wire [31:0] and_22;
  wire [31:0] and_23;
  wire [31:0] and_24;
  wire [31:0] and_25;
  wire [31:0] and_26;
  wire [31:0] and_27;
  wire [31:0] and_28;
  wire [31:0] and_29;
  wire [31:0] and_3;
  wire [31:0] and_30;
  wire [31:0] and_31;
  wire [31:0] and_4;
  wire [31:0] and_5;
  wire [31:0] and_6;
  wire [31:0] and_7;
  wire [31:0] and_8;
  wire [31:0] and_9;
  wire [31:0] nand_0;
  wire [31:0] nand_1;
  wire [31:0] nand_10;
  wire [31:0] nand_11;
  wire [31:0] nand_12;
  wire [31:0] nand_13;
  wire [31:0] nand_14;
  wire [31:0] nand_15;
  wire [31:0] nand_16;
  wire [31:0] nand_17;
  wire [31:0] nand_18;
  wire [31:0] nand_19;
  wire [31:0] nand_2;
  wire [31:0] nand_20;
  wire [31:0] nand_21;
  wire [31:0] nand_22;
  wire [31:0] nand_23;
  wire [31:0] nand_24;
  wire [31:0] nand_25;
  wire [31:0] nand_26;
  wire [31:0] nand_27;
  wire [31:0] nand_28;
  wire [31:0] nand_29;
  wire [31:0] nand_3;
  wire [31:0] nand_30;
  wire [31:0] nand_31;
  wire [31:0] nand_4;
  wire [31:0] nand_5;
  wire [31:0] nand_6;
  wire [31:0] nand_7;
  wire [31:0] nand_8;
  wire [31:0] nand_9;

  and and_a0_b0 (and_0[0], i0[0], i1[0]);
  and and_a0_b1 (and_1[0], i0[0], i1[1]);
  and and_a0_b10 (and_10[0], i0[0], i1[10]);
  and and_a0_b11 (and_11[0], i0[0], i1[11]);
  and and_a0_b12 (and_12[0], i0[0], i1[12]);
  and and_a0_b13 (and_13[0], i0[0], i1[13]);
  and and_a0_b14 (and_14[0], i0[0], i1[14]);
  and and_a0_b15 (and_15[0], i0[0], i1[15]);
  and and_a0_b16 (and_16[0], i0[0], i1[16]);
  and and_a0_b17 (and_17[0], i0[0], i1[17]);
  and and_a0_b18 (and_18[0], i0[0], i1[18]);
  and and_a0_b19 (and_19[0], i0[0], i1[19]);
  and and_a0_b2 (and_2[0], i0[0], i1[2]);
  and and_a0_b20 (and_20[0], i0[0], i1[20]);
  and and_a0_b21 (and_21[0], i0[0], i1[21]);
  and and_a0_b22 (and_22[0], i0[0], i1[22]);
  and and_a0_b23 (and_23[0], i0[0], i1[23]);
  and and_a0_b24 (and_24[0], i0[0], i1[24]);
  and and_a0_b25 (and_25[0], i0[0], i1[25]);
  and and_a0_b26 (and_26[0], i0[0], i1[26]);
  and and_a0_b27 (and_27[0], i0[0], i1[27]);
  and and_a0_b28 (and_28[0], i0[0], i1[28]);
  and and_a0_b29 (and_29[0], i0[0], i1[29]);
  and and_a0_b3 (and_3[0], i0[0], i1[3]);
  and and_a0_b30 (and_30[0], i0[0], i1[30]);
  and and_a0_b31 (nand_31[0], i0[0], i1[31]);
  and and_a0_b4 (and_4[0], i0[0], i1[4]);
  and and_a0_b5 (and_5[0], i0[0], i1[5]);
  and and_a0_b6 (and_6[0], i0[0], i1[6]);
  and and_a0_b7 (and_7[0], i0[0], i1[7]);
  and and_a0_b8 (and_8[0], i0[0], i1[8]);
  and and_a0_b9 (and_9[0], i0[0], i1[9]);
  and and_a10_b0 (and_0[10], i0[10], i1[0]);
  and and_a10_b1 (and_1[10], i0[10], i1[1]);
  and and_a10_b10 (and_10[10], i0[10], i1[10]);
  and and_a10_b11 (and_11[10], i0[10], i1[11]);
  and and_a10_b12 (and_12[10], i0[10], i1[12]);
  and and_a10_b13 (and_13[10], i0[10], i1[13]);
  and and_a10_b14 (and_14[10], i0[10], i1[14]);
  and and_a10_b15 (and_15[10], i0[10], i1[15]);
  and and_a10_b16 (and_16[10], i0[10], i1[16]);
  and and_a10_b17 (and_17[10], i0[10], i1[17]);
  and and_a10_b18 (and_18[10], i0[10], i1[18]);
  and and_a10_b19 (and_19[10], i0[10], i1[19]);
  and and_a10_b2 (and_2[10], i0[10], i1[2]);
  and and_a10_b20 (and_20[10], i0[10], i1[20]);
  and and_a10_b21 (and_21[10], i0[10], i1[21]);
  and and_a10_b22 (and_22[10], i0[10], i1[22]);
  and and_a10_b23 (and_23[10], i0[10], i1[23]);
  and and_a10_b24 (and_24[10], i0[10], i1[24]);
  and and_a10_b25 (and_25[10], i0[10], i1[25]);
  and and_a10_b26 (and_26[10], i0[10], i1[26]);
  and and_a10_b27 (and_27[10], i0[10], i1[27]);
  and and_a10_b28 (and_28[10], i0[10], i1[28]);
  and and_a10_b29 (and_29[10], i0[10], i1[29]);
  and and_a10_b3 (and_3[10], i0[10], i1[3]);
  and and_a10_b30 (and_30[10], i0[10], i1[30]);
  and and_a10_b31 (nand_31[10], i0[10], i1[31]);
  and and_a10_b4 (and_4[10], i0[10], i1[4]);
  and and_a10_b5 (and_5[10], i0[10], i1[5]);
  and and_a10_b6 (and_6[10], i0[10], i1[6]);
  and and_a10_b7 (and_7[10], i0[10], i1[7]);
  and and_a10_b8 (and_8[10], i0[10], i1[8]);
  and and_a10_b9 (and_9[10], i0[10], i1[9]);
  and and_a11_b0 (and_0[11], i0[11], i1[0]);
  and and_a11_b1 (and_1[11], i0[11], i1[1]);
  and and_a11_b10 (and_10[11], i0[11], i1[10]);
  and and_a11_b11 (and_11[11], i0[11], i1[11]);
  and and_a11_b12 (and_12[11], i0[11], i1[12]);
  and and_a11_b13 (and_13[11], i0[11], i1[13]);
  and and_a11_b14 (and_14[11], i0[11], i1[14]);
  and and_a11_b15 (and_15[11], i0[11], i1[15]);
  and and_a11_b16 (and_16[11], i0[11], i1[16]);
  and and_a11_b17 (and_17[11], i0[11], i1[17]);
  and and_a11_b18 (and_18[11], i0[11], i1[18]);
  and and_a11_b19 (and_19[11], i0[11], i1[19]);
  and and_a11_b2 (and_2[11], i0[11], i1[2]);
  and and_a11_b20 (and_20[11], i0[11], i1[20]);
  and and_a11_b21 (and_21[11], i0[11], i1[21]);
  and and_a11_b22 (and_22[11], i0[11], i1[22]);
  and and_a11_b23 (and_23[11], i0[11], i1[23]);
  and and_a11_b24 (and_24[11], i0[11], i1[24]);
  and and_a11_b25 (and_25[11], i0[11], i1[25]);
  and and_a11_b26 (and_26[11], i0[11], i1[26]);
  and and_a11_b27 (and_27[11], i0[11], i1[27]);
  and and_a11_b28 (and_28[11], i0[11], i1[28]);
  and and_a11_b29 (and_29[11], i0[11], i1[29]);
  and and_a11_b3 (and_3[11], i0[11], i1[3]);
  and and_a11_b30 (and_30[11], i0[11], i1[30]);
  and and_a11_b31 (nand_31[11], i0[11], i1[31]);
  and and_a11_b4 (and_4[11], i0[11], i1[4]);
  and and_a11_b5 (and_5[11], i0[11], i1[5]);
  and and_a11_b6 (and_6[11], i0[11], i1[6]);
  and and_a11_b7 (and_7[11], i0[11], i1[7]);
  and and_a11_b8 (and_8[11], i0[11], i1[8]);
  and and_a11_b9 (and_9[11], i0[11], i1[9]);
  and and_a12_b0 (and_0[12], i0[12], i1[0]);
  and and_a12_b1 (and_1[12], i0[12], i1[1]);
  and and_a12_b10 (and_10[12], i0[12], i1[10]);
  and and_a12_b11 (and_11[12], i0[12], i1[11]);
  and and_a12_b12 (and_12[12], i0[12], i1[12]);
  and and_a12_b13 (and_13[12], i0[12], i1[13]);
  and and_a12_b14 (and_14[12], i0[12], i1[14]);
  and and_a12_b15 (and_15[12], i0[12], i1[15]);
  and and_a12_b16 (and_16[12], i0[12], i1[16]);
  and and_a12_b17 (and_17[12], i0[12], i1[17]);
  and and_a12_b18 (and_18[12], i0[12], i1[18]);
  and and_a12_b19 (and_19[12], i0[12], i1[19]);
  and and_a12_b2 (and_2[12], i0[12], i1[2]);
  and and_a12_b20 (and_20[12], i0[12], i1[20]);
  and and_a12_b21 (and_21[12], i0[12], i1[21]);
  and and_a12_b22 (and_22[12], i0[12], i1[22]);
  and and_a12_b23 (and_23[12], i0[12], i1[23]);
  and and_a12_b24 (and_24[12], i0[12], i1[24]);
  and and_a12_b25 (and_25[12], i0[12], i1[25]);
  and and_a12_b26 (and_26[12], i0[12], i1[26]);
  and and_a12_b27 (and_27[12], i0[12], i1[27]);
  and and_a12_b28 (and_28[12], i0[12], i1[28]);
  and and_a12_b29 (and_29[12], i0[12], i1[29]);
  and and_a12_b3 (and_3[12], i0[12], i1[3]);
  and and_a12_b30 (and_30[12], i0[12], i1[30]);
  and and_a12_b31 (nand_31[12], i0[12], i1[31]);
  and and_a12_b4 (and_4[12], i0[12], i1[4]);
  and and_a12_b5 (and_5[12], i0[12], i1[5]);
  and and_a12_b6 (and_6[12], i0[12], i1[6]);
  and and_a12_b7 (and_7[12], i0[12], i1[7]);
  and and_a12_b8 (and_8[12], i0[12], i1[8]);
  and and_a12_b9 (and_9[12], i0[12], i1[9]);
  and and_a13_b0 (and_0[13], i0[13], i1[0]);
  and and_a13_b1 (and_1[13], i0[13], i1[1]);
  and and_a13_b10 (and_10[13], i0[13], i1[10]);
  and and_a13_b11 (and_11[13], i0[13], i1[11]);
  and and_a13_b12 (and_12[13], i0[13], i1[12]);
  and and_a13_b13 (and_13[13], i0[13], i1[13]);
  and and_a13_b14 (and_14[13], i0[13], i1[14]);
  and and_a13_b15 (and_15[13], i0[13], i1[15]);
  and and_a13_b16 (and_16[13], i0[13], i1[16]);
  and and_a13_b17 (and_17[13], i0[13], i1[17]);
  and and_a13_b18 (and_18[13], i0[13], i1[18]);
  and and_a13_b19 (and_19[13], i0[13], i1[19]);
  and and_a13_b2 (and_2[13], i0[13], i1[2]);
  and and_a13_b20 (and_20[13], i0[13], i1[20]);
  and and_a13_b21 (and_21[13], i0[13], i1[21]);
  and and_a13_b22 (and_22[13], i0[13], i1[22]);
  and and_a13_b23 (and_23[13], i0[13], i1[23]);
  and and_a13_b24 (and_24[13], i0[13], i1[24]);
  and and_a13_b25 (and_25[13], i0[13], i1[25]);
  and and_a13_b26 (and_26[13], i0[13], i1[26]);
  and and_a13_b27 (and_27[13], i0[13], i1[27]);
  and and_a13_b28 (and_28[13], i0[13], i1[28]);
  and and_a13_b29 (and_29[13], i0[13], i1[29]);
  and and_a13_b3 (and_3[13], i0[13], i1[3]);
  and and_a13_b30 (and_30[13], i0[13], i1[30]);
  and and_a13_b31 (nand_31[13], i0[13], i1[31]);
  and and_a13_b4 (and_4[13], i0[13], i1[4]);
  and and_a13_b5 (and_5[13], i0[13], i1[5]);
  and and_a13_b6 (and_6[13], i0[13], i1[6]);
  and and_a13_b7 (and_7[13], i0[13], i1[7]);
  and and_a13_b8 (and_8[13], i0[13], i1[8]);
  and and_a13_b9 (and_9[13], i0[13], i1[9]);
  and and_a14_b0 (and_0[14], i0[14], i1[0]);
  and and_a14_b1 (and_1[14], i0[14], i1[1]);
  and and_a14_b10 (and_10[14], i0[14], i1[10]);
  and and_a14_b11 (and_11[14], i0[14], i1[11]);
  and and_a14_b12 (and_12[14], i0[14], i1[12]);
  and and_a14_b13 (and_13[14], i0[14], i1[13]);
  and and_a14_b14 (and_14[14], i0[14], i1[14]);
  and and_a14_b15 (and_15[14], i0[14], i1[15]);
  and and_a14_b16 (and_16[14], i0[14], i1[16]);
  and and_a14_b17 (and_17[14], i0[14], i1[17]);
  and and_a14_b18 (and_18[14], i0[14], i1[18]);
  and and_a14_b19 (and_19[14], i0[14], i1[19]);
  and and_a14_b2 (and_2[14], i0[14], i1[2]);
  and and_a14_b20 (and_20[14], i0[14], i1[20]);
  and and_a14_b21 (and_21[14], i0[14], i1[21]);
  and and_a14_b22 (and_22[14], i0[14], i1[22]);
  and and_a14_b23 (and_23[14], i0[14], i1[23]);
  and and_a14_b24 (and_24[14], i0[14], i1[24]);
  and and_a14_b25 (and_25[14], i0[14], i1[25]);
  and and_a14_b26 (and_26[14], i0[14], i1[26]);
  and and_a14_b27 (and_27[14], i0[14], i1[27]);
  and and_a14_b28 (and_28[14], i0[14], i1[28]);
  and and_a14_b29 (and_29[14], i0[14], i1[29]);
  and and_a14_b3 (and_3[14], i0[14], i1[3]);
  and and_a14_b30 (and_30[14], i0[14], i1[30]);
  and and_a14_b31 (nand_31[14], i0[14], i1[31]);
  and and_a14_b4 (and_4[14], i0[14], i1[4]);
  and and_a14_b5 (and_5[14], i0[14], i1[5]);
  and and_a14_b6 (and_6[14], i0[14], i1[6]);
  and and_a14_b7 (and_7[14], i0[14], i1[7]);
  and and_a14_b8 (and_8[14], i0[14], i1[8]);
  and and_a14_b9 (and_9[14], i0[14], i1[9]);
  and and_a15_b0 (and_0[15], i0[15], i1[0]);
  and and_a15_b1 (and_1[15], i0[15], i1[1]);
  and and_a15_b10 (and_10[15], i0[15], i1[10]);
  and and_a15_b11 (and_11[15], i0[15], i1[11]);
  and and_a15_b12 (and_12[15], i0[15], i1[12]);
  and and_a15_b13 (and_13[15], i0[15], i1[13]);
  and and_a15_b14 (and_14[15], i0[15], i1[14]);
  and and_a15_b15 (and_15[15], i0[15], i1[15]);
  and and_a15_b16 (and_16[15], i0[15], i1[16]);
  and and_a15_b17 (and_17[15], i0[15], i1[17]);
  and and_a15_b18 (and_18[15], i0[15], i1[18]);
  and and_a15_b19 (and_19[15], i0[15], i1[19]);
  and and_a15_b2 (and_2[15], i0[15], i1[2]);
  and and_a15_b20 (and_20[15], i0[15], i1[20]);
  and and_a15_b21 (and_21[15], i0[15], i1[21]);
  and and_a15_b22 (and_22[15], i0[15], i1[22]);
  and and_a15_b23 (and_23[15], i0[15], i1[23]);
  and and_a15_b24 (and_24[15], i0[15], i1[24]);
  and and_a15_b25 (and_25[15], i0[15], i1[25]);
  and and_a15_b26 (and_26[15], i0[15], i1[26]);
  and and_a15_b27 (and_27[15], i0[15], i1[27]);
  and and_a15_b28 (and_28[15], i0[15], i1[28]);
  and and_a15_b29 (and_29[15], i0[15], i1[29]);
  and and_a15_b3 (and_3[15], i0[15], i1[3]);
  and and_a15_b30 (and_30[15], i0[15], i1[30]);
  and and_a15_b31 (nand_31[15], i0[15], i1[31]);
  and and_a15_b4 (and_4[15], i0[15], i1[4]);
  and and_a15_b5 (and_5[15], i0[15], i1[5]);
  and and_a15_b6 (and_6[15], i0[15], i1[6]);
  and and_a15_b7 (and_7[15], i0[15], i1[7]);
  and and_a15_b8 (and_8[15], i0[15], i1[8]);
  and and_a15_b9 (and_9[15], i0[15], i1[9]);
  and and_a16_b0 (and_0[16], i0[16], i1[0]);
  and and_a16_b1 (and_1[16], i0[16], i1[1]);
  and and_a16_b10 (and_10[16], i0[16], i1[10]);
  and and_a16_b11 (and_11[16], i0[16], i1[11]);
  and and_a16_b12 (and_12[16], i0[16], i1[12]);
  and and_a16_b13 (and_13[16], i0[16], i1[13]);
  and and_a16_b14 (and_14[16], i0[16], i1[14]);
  and and_a16_b15 (and_15[16], i0[16], i1[15]);
  and and_a16_b16 (and_16[16], i0[16], i1[16]);
  and and_a16_b17 (and_17[16], i0[16], i1[17]);
  and and_a16_b18 (and_18[16], i0[16], i1[18]);
  and and_a16_b19 (and_19[16], i0[16], i1[19]);
  and and_a16_b2 (and_2[16], i0[16], i1[2]);
  and and_a16_b20 (and_20[16], i0[16], i1[20]);
  and and_a16_b21 (and_21[16], i0[16], i1[21]);
  and and_a16_b22 (and_22[16], i0[16], i1[22]);
  and and_a16_b23 (and_23[16], i0[16], i1[23]);
  and and_a16_b24 (and_24[16], i0[16], i1[24]);
  and and_a16_b25 (and_25[16], i0[16], i1[25]);
  and and_a16_b26 (and_26[16], i0[16], i1[26]);
  and and_a16_b27 (and_27[16], i0[16], i1[27]);
  and and_a16_b28 (and_28[16], i0[16], i1[28]);
  and and_a16_b29 (and_29[16], i0[16], i1[29]);
  and and_a16_b3 (and_3[16], i0[16], i1[3]);
  and and_a16_b30 (and_30[16], i0[16], i1[30]);
  and and_a16_b31 (nand_31[16], i0[16], i1[31]);
  and and_a16_b4 (and_4[16], i0[16], i1[4]);
  and and_a16_b5 (and_5[16], i0[16], i1[5]);
  and and_a16_b6 (and_6[16], i0[16], i1[6]);
  and and_a16_b7 (and_7[16], i0[16], i1[7]);
  and and_a16_b8 (and_8[16], i0[16], i1[8]);
  and and_a16_b9 (and_9[16], i0[16], i1[9]);
  and and_a17_b0 (and_0[17], i0[17], i1[0]);
  and and_a17_b1 (and_1[17], i0[17], i1[1]);
  and and_a17_b10 (and_10[17], i0[17], i1[10]);
  and and_a17_b11 (and_11[17], i0[17], i1[11]);
  and and_a17_b12 (and_12[17], i0[17], i1[12]);
  and and_a17_b13 (and_13[17], i0[17], i1[13]);
  and and_a17_b14 (and_14[17], i0[17], i1[14]);
  and and_a17_b15 (and_15[17], i0[17], i1[15]);
  and and_a17_b16 (and_16[17], i0[17], i1[16]);
  and and_a17_b17 (and_17[17], i0[17], i1[17]);
  and and_a17_b18 (and_18[17], i0[17], i1[18]);
  and and_a17_b19 (and_19[17], i0[17], i1[19]);
  and and_a17_b2 (and_2[17], i0[17], i1[2]);
  and and_a17_b20 (and_20[17], i0[17], i1[20]);
  and and_a17_b21 (and_21[17], i0[17], i1[21]);
  and and_a17_b22 (and_22[17], i0[17], i1[22]);
  and and_a17_b23 (and_23[17], i0[17], i1[23]);
  and and_a17_b24 (and_24[17], i0[17], i1[24]);
  and and_a17_b25 (and_25[17], i0[17], i1[25]);
  and and_a17_b26 (and_26[17], i0[17], i1[26]);
  and and_a17_b27 (and_27[17], i0[17], i1[27]);
  and and_a17_b28 (and_28[17], i0[17], i1[28]);
  and and_a17_b29 (and_29[17], i0[17], i1[29]);
  and and_a17_b3 (and_3[17], i0[17], i1[3]);
  and and_a17_b30 (and_30[17], i0[17], i1[30]);
  and and_a17_b31 (nand_31[17], i0[17], i1[31]);
  and and_a17_b4 (and_4[17], i0[17], i1[4]);
  and and_a17_b5 (and_5[17], i0[17], i1[5]);
  and and_a17_b6 (and_6[17], i0[17], i1[6]);
  and and_a17_b7 (and_7[17], i0[17], i1[7]);
  and and_a17_b8 (and_8[17], i0[17], i1[8]);
  and and_a17_b9 (and_9[17], i0[17], i1[9]);
  and and_a18_b0 (and_0[18], i0[18], i1[0]);
  and and_a18_b1 (and_1[18], i0[18], i1[1]);
  and and_a18_b10 (and_10[18], i0[18], i1[10]);
  and and_a18_b11 (and_11[18], i0[18], i1[11]);
  and and_a18_b12 (and_12[18], i0[18], i1[12]);
  and and_a18_b13 (and_13[18], i0[18], i1[13]);
  and and_a18_b14 (and_14[18], i0[18], i1[14]);
  and and_a18_b15 (and_15[18], i0[18], i1[15]);
  and and_a18_b16 (and_16[18], i0[18], i1[16]);
  and and_a18_b17 (and_17[18], i0[18], i1[17]);
  and and_a18_b18 (and_18[18], i0[18], i1[18]);
  and and_a18_b19 (and_19[18], i0[18], i1[19]);
  and and_a18_b2 (and_2[18], i0[18], i1[2]);
  and and_a18_b20 (and_20[18], i0[18], i1[20]);
  and and_a18_b21 (and_21[18], i0[18], i1[21]);
  and and_a18_b22 (and_22[18], i0[18], i1[22]);
  and and_a18_b23 (and_23[18], i0[18], i1[23]);
  and and_a18_b24 (and_24[18], i0[18], i1[24]);
  and and_a18_b25 (and_25[18], i0[18], i1[25]);
  and and_a18_b26 (and_26[18], i0[18], i1[26]);
  and and_a18_b27 (and_27[18], i0[18], i1[27]);
  and and_a18_b28 (and_28[18], i0[18], i1[28]);
  and and_a18_b29 (and_29[18], i0[18], i1[29]);
  and and_a18_b3 (and_3[18], i0[18], i1[3]);
  and and_a18_b30 (and_30[18], i0[18], i1[30]);
  and and_a18_b31 (nand_31[18], i0[18], i1[31]);
  and and_a18_b4 (and_4[18], i0[18], i1[4]);
  and and_a18_b5 (and_5[18], i0[18], i1[5]);
  and and_a18_b6 (and_6[18], i0[18], i1[6]);
  and and_a18_b7 (and_7[18], i0[18], i1[7]);
  and and_a18_b8 (and_8[18], i0[18], i1[8]);
  and and_a18_b9 (and_9[18], i0[18], i1[9]);
  and and_a19_b0 (and_0[19], i0[19], i1[0]);
  and and_a19_b1 (and_1[19], i0[19], i1[1]);
  and and_a19_b10 (and_10[19], i0[19], i1[10]);
  and and_a19_b11 (and_11[19], i0[19], i1[11]);
  and and_a19_b12 (and_12[19], i0[19], i1[12]);
  and and_a19_b13 (and_13[19], i0[19], i1[13]);
  and and_a19_b14 (and_14[19], i0[19], i1[14]);
  and and_a19_b15 (and_15[19], i0[19], i1[15]);
  and and_a19_b16 (and_16[19], i0[19], i1[16]);
  and and_a19_b17 (and_17[19], i0[19], i1[17]);
  and and_a19_b18 (and_18[19], i0[19], i1[18]);
  and and_a19_b19 (and_19[19], i0[19], i1[19]);
  and and_a19_b2 (and_2[19], i0[19], i1[2]);
  and and_a19_b20 (and_20[19], i0[19], i1[20]);
  and and_a19_b21 (and_21[19], i0[19], i1[21]);
  and and_a19_b22 (and_22[19], i0[19], i1[22]);
  and and_a19_b23 (and_23[19], i0[19], i1[23]);
  and and_a19_b24 (and_24[19], i0[19], i1[24]);
  and and_a19_b25 (and_25[19], i0[19], i1[25]);
  and and_a19_b26 (and_26[19], i0[19], i1[26]);
  and and_a19_b27 (and_27[19], i0[19], i1[27]);
  and and_a19_b28 (and_28[19], i0[19], i1[28]);
  and and_a19_b29 (and_29[19], i0[19], i1[29]);
  and and_a19_b3 (and_3[19], i0[19], i1[3]);
  and and_a19_b30 (and_30[19], i0[19], i1[30]);
  and and_a19_b31 (nand_31[19], i0[19], i1[31]);
  and and_a19_b4 (and_4[19], i0[19], i1[4]);
  and and_a19_b5 (and_5[19], i0[19], i1[5]);
  and and_a19_b6 (and_6[19], i0[19], i1[6]);
  and and_a19_b7 (and_7[19], i0[19], i1[7]);
  and and_a19_b8 (and_8[19], i0[19], i1[8]);
  and and_a19_b9 (and_9[19], i0[19], i1[9]);
  and and_a1_b0 (and_0[1], i0[1], i1[0]);
  and and_a1_b1 (and_1[1], i0[1], i1[1]);
  and and_a1_b10 (and_10[1], i0[1], i1[10]);
  and and_a1_b11 (and_11[1], i0[1], i1[11]);
  and and_a1_b12 (and_12[1], i0[1], i1[12]);
  and and_a1_b13 (and_13[1], i0[1], i1[13]);
  and and_a1_b14 (and_14[1], i0[1], i1[14]);
  and and_a1_b15 (and_15[1], i0[1], i1[15]);
  and and_a1_b16 (and_16[1], i0[1], i1[16]);
  and and_a1_b17 (and_17[1], i0[1], i1[17]);
  and and_a1_b18 (and_18[1], i0[1], i1[18]);
  and and_a1_b19 (and_19[1], i0[1], i1[19]);
  and and_a1_b2 (and_2[1], i0[1], i1[2]);
  and and_a1_b20 (and_20[1], i0[1], i1[20]);
  and and_a1_b21 (and_21[1], i0[1], i1[21]);
  and and_a1_b22 (and_22[1], i0[1], i1[22]);
  and and_a1_b23 (and_23[1], i0[1], i1[23]);
  and and_a1_b24 (and_24[1], i0[1], i1[24]);
  and and_a1_b25 (and_25[1], i0[1], i1[25]);
  and and_a1_b26 (and_26[1], i0[1], i1[26]);
  and and_a1_b27 (and_27[1], i0[1], i1[27]);
  and and_a1_b28 (and_28[1], i0[1], i1[28]);
  and and_a1_b29 (and_29[1], i0[1], i1[29]);
  and and_a1_b3 (and_3[1], i0[1], i1[3]);
  and and_a1_b30 (and_30[1], i0[1], i1[30]);
  and and_a1_b31 (nand_31[1], i0[1], i1[31]);
  and and_a1_b4 (and_4[1], i0[1], i1[4]);
  and and_a1_b5 (and_5[1], i0[1], i1[5]);
  and and_a1_b6 (and_6[1], i0[1], i1[6]);
  and and_a1_b7 (and_7[1], i0[1], i1[7]);
  and and_a1_b8 (and_8[1], i0[1], i1[8]);
  and and_a1_b9 (and_9[1], i0[1], i1[9]);
  and and_a20_b0 (and_0[20], i0[20], i1[0]);
  and and_a20_b1 (and_1[20], i0[20], i1[1]);
  and and_a20_b10 (and_10[20], i0[20], i1[10]);
  and and_a20_b11 (and_11[20], i0[20], i1[11]);
  and and_a20_b12 (and_12[20], i0[20], i1[12]);
  and and_a20_b13 (and_13[20], i0[20], i1[13]);
  and and_a20_b14 (and_14[20], i0[20], i1[14]);
  and and_a20_b15 (and_15[20], i0[20], i1[15]);
  and and_a20_b16 (and_16[20], i0[20], i1[16]);
  and and_a20_b17 (and_17[20], i0[20], i1[17]);
  and and_a20_b18 (and_18[20], i0[20], i1[18]);
  and and_a20_b19 (and_19[20], i0[20], i1[19]);
  and and_a20_b2 (and_2[20], i0[20], i1[2]);
  and and_a20_b20 (and_20[20], i0[20], i1[20]);
  and and_a20_b21 (and_21[20], i0[20], i1[21]);
  and and_a20_b22 (and_22[20], i0[20], i1[22]);
  and and_a20_b23 (and_23[20], i0[20], i1[23]);
  and and_a20_b24 (and_24[20], i0[20], i1[24]);
  and and_a20_b25 (and_25[20], i0[20], i1[25]);
  and and_a20_b26 (and_26[20], i0[20], i1[26]);
  and and_a20_b27 (and_27[20], i0[20], i1[27]);
  and and_a20_b28 (and_28[20], i0[20], i1[28]);
  and and_a20_b29 (and_29[20], i0[20], i1[29]);
  and and_a20_b3 (and_3[20], i0[20], i1[3]);
  and and_a20_b30 (and_30[20], i0[20], i1[30]);
  and and_a20_b31 (nand_31[20], i0[20], i1[31]);
  and and_a20_b4 (and_4[20], i0[20], i1[4]);
  and and_a20_b5 (and_5[20], i0[20], i1[5]);
  and and_a20_b6 (and_6[20], i0[20], i1[6]);
  and and_a20_b7 (and_7[20], i0[20], i1[7]);
  and and_a20_b8 (and_8[20], i0[20], i1[8]);
  and and_a20_b9 (and_9[20], i0[20], i1[9]);
  and and_a21_b0 (and_0[21], i0[21], i1[0]);
  and and_a21_b1 (and_1[21], i0[21], i1[1]);
  and and_a21_b10 (and_10[21], i0[21], i1[10]);
  and and_a21_b11 (and_11[21], i0[21], i1[11]);
  and and_a21_b12 (and_12[21], i0[21], i1[12]);
  and and_a21_b13 (and_13[21], i0[21], i1[13]);
  and and_a21_b14 (and_14[21], i0[21], i1[14]);
  and and_a21_b15 (and_15[21], i0[21], i1[15]);
  and and_a21_b16 (and_16[21], i0[21], i1[16]);
  and and_a21_b17 (and_17[21], i0[21], i1[17]);
  and and_a21_b18 (and_18[21], i0[21], i1[18]);
  and and_a21_b19 (and_19[21], i0[21], i1[19]);
  and and_a21_b2 (and_2[21], i0[21], i1[2]);
  and and_a21_b20 (and_20[21], i0[21], i1[20]);
  and and_a21_b21 (and_21[21], i0[21], i1[21]);
  and and_a21_b22 (and_22[21], i0[21], i1[22]);
  and and_a21_b23 (and_23[21], i0[21], i1[23]);
  and and_a21_b24 (and_24[21], i0[21], i1[24]);
  and and_a21_b25 (and_25[21], i0[21], i1[25]);
  and and_a21_b26 (and_26[21], i0[21], i1[26]);
  and and_a21_b27 (and_27[21], i0[21], i1[27]);
  and and_a21_b28 (and_28[21], i0[21], i1[28]);
  and and_a21_b29 (and_29[21], i0[21], i1[29]);
  and and_a21_b3 (and_3[21], i0[21], i1[3]);
  and and_a21_b30 (and_30[21], i0[21], i1[30]);
  and and_a21_b31 (nand_31[21], i0[21], i1[31]);
  and and_a21_b4 (and_4[21], i0[21], i1[4]);
  and and_a21_b5 (and_5[21], i0[21], i1[5]);
  and and_a21_b6 (and_6[21], i0[21], i1[6]);
  and and_a21_b7 (and_7[21], i0[21], i1[7]);
  and and_a21_b8 (and_8[21], i0[21], i1[8]);
  and and_a21_b9 (and_9[21], i0[21], i1[9]);
  and and_a22_b0 (and_0[22], i0[22], i1[0]);
  and and_a22_b1 (and_1[22], i0[22], i1[1]);
  and and_a22_b10 (and_10[22], i0[22], i1[10]);
  and and_a22_b11 (and_11[22], i0[22], i1[11]);
  and and_a22_b12 (and_12[22], i0[22], i1[12]);
  and and_a22_b13 (and_13[22], i0[22], i1[13]);
  and and_a22_b14 (and_14[22], i0[22], i1[14]);
  and and_a22_b15 (and_15[22], i0[22], i1[15]);
  and and_a22_b16 (and_16[22], i0[22], i1[16]);
  and and_a22_b17 (and_17[22], i0[22], i1[17]);
  and and_a22_b18 (and_18[22], i0[22], i1[18]);
  and and_a22_b19 (and_19[22], i0[22], i1[19]);
  and and_a22_b2 (and_2[22], i0[22], i1[2]);
  and and_a22_b20 (and_20[22], i0[22], i1[20]);
  and and_a22_b21 (and_21[22], i0[22], i1[21]);
  and and_a22_b22 (and_22[22], i0[22], i1[22]);
  and and_a22_b23 (and_23[22], i0[22], i1[23]);
  and and_a22_b24 (and_24[22], i0[22], i1[24]);
  and and_a22_b25 (and_25[22], i0[22], i1[25]);
  and and_a22_b26 (and_26[22], i0[22], i1[26]);
  and and_a22_b27 (and_27[22], i0[22], i1[27]);
  and and_a22_b28 (and_28[22], i0[22], i1[28]);
  and and_a22_b29 (and_29[22], i0[22], i1[29]);
  and and_a22_b3 (and_3[22], i0[22], i1[3]);
  and and_a22_b30 (and_30[22], i0[22], i1[30]);
  and and_a22_b31 (nand_31[22], i0[22], i1[31]);
  and and_a22_b4 (and_4[22], i0[22], i1[4]);
  and and_a22_b5 (and_5[22], i0[22], i1[5]);
  and and_a22_b6 (and_6[22], i0[22], i1[6]);
  and and_a22_b7 (and_7[22], i0[22], i1[7]);
  and and_a22_b8 (and_8[22], i0[22], i1[8]);
  and and_a22_b9 (and_9[22], i0[22], i1[9]);
  and and_a23_b0 (and_0[23], i0[23], i1[0]);
  and and_a23_b1 (and_1[23], i0[23], i1[1]);
  and and_a23_b10 (and_10[23], i0[23], i1[10]);
  and and_a23_b11 (and_11[23], i0[23], i1[11]);
  and and_a23_b12 (and_12[23], i0[23], i1[12]);
  and and_a23_b13 (and_13[23], i0[23], i1[13]);
  and and_a23_b14 (and_14[23], i0[23], i1[14]);
  and and_a23_b15 (and_15[23], i0[23], i1[15]);
  and and_a23_b16 (and_16[23], i0[23], i1[16]);
  and and_a23_b17 (and_17[23], i0[23], i1[17]);
  and and_a23_b18 (and_18[23], i0[23], i1[18]);
  and and_a23_b19 (and_19[23], i0[23], i1[19]);
  and and_a23_b2 (and_2[23], i0[23], i1[2]);
  and and_a23_b20 (and_20[23], i0[23], i1[20]);
  and and_a23_b21 (and_21[23], i0[23], i1[21]);
  and and_a23_b22 (and_22[23], i0[23], i1[22]);
  and and_a23_b23 (and_23[23], i0[23], i1[23]);
  and and_a23_b24 (and_24[23], i0[23], i1[24]);
  and and_a23_b25 (and_25[23], i0[23], i1[25]);
  and and_a23_b26 (and_26[23], i0[23], i1[26]);
  and and_a23_b27 (and_27[23], i0[23], i1[27]);
  and and_a23_b28 (and_28[23], i0[23], i1[28]);
  and and_a23_b29 (and_29[23], i0[23], i1[29]);
  and and_a23_b3 (and_3[23], i0[23], i1[3]);
  and and_a23_b30 (and_30[23], i0[23], i1[30]);
  and and_a23_b31 (nand_31[23], i0[23], i1[31]);
  and and_a23_b4 (and_4[23], i0[23], i1[4]);
  and and_a23_b5 (and_5[23], i0[23], i1[5]);
  and and_a23_b6 (and_6[23], i0[23], i1[6]);
  and and_a23_b7 (and_7[23], i0[23], i1[7]);
  and and_a23_b8 (and_8[23], i0[23], i1[8]);
  and and_a23_b9 (and_9[23], i0[23], i1[9]);
  and and_a24_b0 (and_0[24], i0[24], i1[0]);
  and and_a24_b1 (and_1[24], i0[24], i1[1]);
  and and_a24_b10 (and_10[24], i0[24], i1[10]);
  and and_a24_b11 (and_11[24], i0[24], i1[11]);
  and and_a24_b12 (and_12[24], i0[24], i1[12]);
  and and_a24_b13 (and_13[24], i0[24], i1[13]);
  and and_a24_b14 (and_14[24], i0[24], i1[14]);
  and and_a24_b15 (and_15[24], i0[24], i1[15]);
  and and_a24_b16 (and_16[24], i0[24], i1[16]);
  and and_a24_b17 (and_17[24], i0[24], i1[17]);
  and and_a24_b18 (and_18[24], i0[24], i1[18]);
  and and_a24_b19 (and_19[24], i0[24], i1[19]);
  and and_a24_b2 (and_2[24], i0[24], i1[2]);
  and and_a24_b20 (and_20[24], i0[24], i1[20]);
  and and_a24_b21 (and_21[24], i0[24], i1[21]);
  and and_a24_b22 (and_22[24], i0[24], i1[22]);
  and and_a24_b23 (and_23[24], i0[24], i1[23]);
  and and_a24_b24 (and_24[24], i0[24], i1[24]);
  and and_a24_b25 (and_25[24], i0[24], i1[25]);
  and and_a24_b26 (and_26[24], i0[24], i1[26]);
  and and_a24_b27 (and_27[24], i0[24], i1[27]);
  and and_a24_b28 (and_28[24], i0[24], i1[28]);
  and and_a24_b29 (and_29[24], i0[24], i1[29]);
  and and_a24_b3 (and_3[24], i0[24], i1[3]);
  and and_a24_b30 (and_30[24], i0[24], i1[30]);
  and and_a24_b31 (nand_31[24], i0[24], i1[31]);
  and and_a24_b4 (and_4[24], i0[24], i1[4]);
  and and_a24_b5 (and_5[24], i0[24], i1[5]);
  and and_a24_b6 (and_6[24], i0[24], i1[6]);
  and and_a24_b7 (and_7[24], i0[24], i1[7]);
  and and_a24_b8 (and_8[24], i0[24], i1[8]);
  and and_a24_b9 (and_9[24], i0[24], i1[9]);
  and and_a25_b0 (and_0[25], i0[25], i1[0]);
  and and_a25_b1 (and_1[25], i0[25], i1[1]);
  and and_a25_b10 (and_10[25], i0[25], i1[10]);
  and and_a25_b11 (and_11[25], i0[25], i1[11]);
  and and_a25_b12 (and_12[25], i0[25], i1[12]);
  and and_a25_b13 (and_13[25], i0[25], i1[13]);
  and and_a25_b14 (and_14[25], i0[25], i1[14]);
  and and_a25_b15 (and_15[25], i0[25], i1[15]);
  and and_a25_b16 (and_16[25], i0[25], i1[16]);
  and and_a25_b17 (and_17[25], i0[25], i1[17]);
  and and_a25_b18 (and_18[25], i0[25], i1[18]);
  and and_a25_b19 (and_19[25], i0[25], i1[19]);
  and and_a25_b2 (and_2[25], i0[25], i1[2]);
  and and_a25_b20 (and_20[25], i0[25], i1[20]);
  and and_a25_b21 (and_21[25], i0[25], i1[21]);
  and and_a25_b22 (and_22[25], i0[25], i1[22]);
  and and_a25_b23 (and_23[25], i0[25], i1[23]);
  and and_a25_b24 (and_24[25], i0[25], i1[24]);
  and and_a25_b25 (and_25[25], i0[25], i1[25]);
  and and_a25_b26 (and_26[25], i0[25], i1[26]);
  and and_a25_b27 (and_27[25], i0[25], i1[27]);
  and and_a25_b28 (and_28[25], i0[25], i1[28]);
  and and_a25_b29 (and_29[25], i0[25], i1[29]);
  and and_a25_b3 (and_3[25], i0[25], i1[3]);
  and and_a25_b30 (and_30[25], i0[25], i1[30]);
  and and_a25_b31 (nand_31[25], i0[25], i1[31]);
  and and_a25_b4 (and_4[25], i0[25], i1[4]);
  and and_a25_b5 (and_5[25], i0[25], i1[5]);
  and and_a25_b6 (and_6[25], i0[25], i1[6]);
  and and_a25_b7 (and_7[25], i0[25], i1[7]);
  and and_a25_b8 (and_8[25], i0[25], i1[8]);
  and and_a25_b9 (and_9[25], i0[25], i1[9]);
  and and_a26_b0 (and_0[26], i0[26], i1[0]);
  and and_a26_b1 (and_1[26], i0[26], i1[1]);
  and and_a26_b10 (and_10[26], i0[26], i1[10]);
  and and_a26_b11 (and_11[26], i0[26], i1[11]);
  and and_a26_b12 (and_12[26], i0[26], i1[12]);
  and and_a26_b13 (and_13[26], i0[26], i1[13]);
  and and_a26_b14 (and_14[26], i0[26], i1[14]);
  and and_a26_b15 (and_15[26], i0[26], i1[15]);
  and and_a26_b16 (and_16[26], i0[26], i1[16]);
  and and_a26_b17 (and_17[26], i0[26], i1[17]);
  and and_a26_b18 (and_18[26], i0[26], i1[18]);
  and and_a26_b19 (and_19[26], i0[26], i1[19]);
  and and_a26_b2 (and_2[26], i0[26], i1[2]);
  and and_a26_b20 (and_20[26], i0[26], i1[20]);
  and and_a26_b21 (and_21[26], i0[26], i1[21]);
  and and_a26_b22 (and_22[26], i0[26], i1[22]);
  and and_a26_b23 (and_23[26], i0[26], i1[23]);
  and and_a26_b24 (and_24[26], i0[26], i1[24]);
  and and_a26_b25 (and_25[26], i0[26], i1[25]);
  and and_a26_b26 (and_26[26], i0[26], i1[26]);
  and and_a26_b27 (and_27[26], i0[26], i1[27]);
  and and_a26_b28 (and_28[26], i0[26], i1[28]);
  and and_a26_b29 (and_29[26], i0[26], i1[29]);
  and and_a26_b3 (and_3[26], i0[26], i1[3]);
  and and_a26_b30 (and_30[26], i0[26], i1[30]);
  and and_a26_b31 (nand_31[26], i0[26], i1[31]);
  and and_a26_b4 (and_4[26], i0[26], i1[4]);
  and and_a26_b5 (and_5[26], i0[26], i1[5]);
  and and_a26_b6 (and_6[26], i0[26], i1[6]);
  and and_a26_b7 (and_7[26], i0[26], i1[7]);
  and and_a26_b8 (and_8[26], i0[26], i1[8]);
  and and_a26_b9 (and_9[26], i0[26], i1[9]);
  and and_a27_b0 (and_0[27], i0[27], i1[0]);
  and and_a27_b1 (and_1[27], i0[27], i1[1]);
  and and_a27_b10 (and_10[27], i0[27], i1[10]);
  and and_a27_b11 (and_11[27], i0[27], i1[11]);
  and and_a27_b12 (and_12[27], i0[27], i1[12]);
  and and_a27_b13 (and_13[27], i0[27], i1[13]);
  and and_a27_b14 (and_14[27], i0[27], i1[14]);
  and and_a27_b15 (and_15[27], i0[27], i1[15]);
  and and_a27_b16 (and_16[27], i0[27], i1[16]);
  and and_a27_b17 (and_17[27], i0[27], i1[17]);
  and and_a27_b18 (and_18[27], i0[27], i1[18]);
  and and_a27_b19 (and_19[27], i0[27], i1[19]);
  and and_a27_b2 (and_2[27], i0[27], i1[2]);
  and and_a27_b20 (and_20[27], i0[27], i1[20]);
  and and_a27_b21 (and_21[27], i0[27], i1[21]);
  and and_a27_b22 (and_22[27], i0[27], i1[22]);
  and and_a27_b23 (and_23[27], i0[27], i1[23]);
  and and_a27_b24 (and_24[27], i0[27], i1[24]);
  and and_a27_b25 (and_25[27], i0[27], i1[25]);
  and and_a27_b26 (and_26[27], i0[27], i1[26]);
  and and_a27_b27 (and_27[27], i0[27], i1[27]);
  and and_a27_b28 (and_28[27], i0[27], i1[28]);
  and and_a27_b29 (and_29[27], i0[27], i1[29]);
  and and_a27_b3 (and_3[27], i0[27], i1[3]);
  and and_a27_b30 (and_30[27], i0[27], i1[30]);
  and and_a27_b31 (nand_31[27], i0[27], i1[31]);
  and and_a27_b4 (and_4[27], i0[27], i1[4]);
  and and_a27_b5 (and_5[27], i0[27], i1[5]);
  and and_a27_b6 (and_6[27], i0[27], i1[6]);
  and and_a27_b7 (and_7[27], i0[27], i1[7]);
  and and_a27_b8 (and_8[27], i0[27], i1[8]);
  and and_a27_b9 (and_9[27], i0[27], i1[9]);
  and and_a28_b0 (and_0[28], i0[28], i1[0]);
  and and_a28_b1 (and_1[28], i0[28], i1[1]);
  and and_a28_b10 (and_10[28], i0[28], i1[10]);
  and and_a28_b11 (and_11[28], i0[28], i1[11]);
  and and_a28_b12 (and_12[28], i0[28], i1[12]);
  and and_a28_b13 (and_13[28], i0[28], i1[13]);
  and and_a28_b14 (and_14[28], i0[28], i1[14]);
  and and_a28_b15 (and_15[28], i0[28], i1[15]);
  and and_a28_b16 (and_16[28], i0[28], i1[16]);
  and and_a28_b17 (and_17[28], i0[28], i1[17]);
  and and_a28_b18 (and_18[28], i0[28], i1[18]);
  and and_a28_b19 (and_19[28], i0[28], i1[19]);
  and and_a28_b2 (and_2[28], i0[28], i1[2]);
  and and_a28_b20 (and_20[28], i0[28], i1[20]);
  and and_a28_b21 (and_21[28], i0[28], i1[21]);
  and and_a28_b22 (and_22[28], i0[28], i1[22]);
  and and_a28_b23 (and_23[28], i0[28], i1[23]);
  and and_a28_b24 (and_24[28], i0[28], i1[24]);
  and and_a28_b25 (and_25[28], i0[28], i1[25]);
  and and_a28_b26 (and_26[28], i0[28], i1[26]);
  and and_a28_b27 (and_27[28], i0[28], i1[27]);
  and and_a28_b28 (and_28[28], i0[28], i1[28]);
  and and_a28_b29 (and_29[28], i0[28], i1[29]);
  and and_a28_b3 (and_3[28], i0[28], i1[3]);
  and and_a28_b30 (and_30[28], i0[28], i1[30]);
  and and_a28_b31 (nand_31[28], i0[28], i1[31]);
  and and_a28_b4 (and_4[28], i0[28], i1[4]);
  and and_a28_b5 (and_5[28], i0[28], i1[5]);
  and and_a28_b6 (and_6[28], i0[28], i1[6]);
  and and_a28_b7 (and_7[28], i0[28], i1[7]);
  and and_a28_b8 (and_8[28], i0[28], i1[8]);
  and and_a28_b9 (and_9[28], i0[28], i1[9]);
  and and_a29_b0 (and_0[29], i0[29], i1[0]);
  and and_a29_b1 (and_1[29], i0[29], i1[1]);
  and and_a29_b10 (and_10[29], i0[29], i1[10]);
  and and_a29_b11 (and_11[29], i0[29], i1[11]);
  and and_a29_b12 (and_12[29], i0[29], i1[12]);
  and and_a29_b13 (and_13[29], i0[29], i1[13]);
  and and_a29_b14 (and_14[29], i0[29], i1[14]);
  and and_a29_b15 (and_15[29], i0[29], i1[15]);
  and and_a29_b16 (and_16[29], i0[29], i1[16]);
  and and_a29_b17 (and_17[29], i0[29], i1[17]);
  and and_a29_b18 (and_18[29], i0[29], i1[18]);
  and and_a29_b19 (and_19[29], i0[29], i1[19]);
  and and_a29_b2 (and_2[29], i0[29], i1[2]);
  and and_a29_b20 (and_20[29], i0[29], i1[20]);
  and and_a29_b21 (and_21[29], i0[29], i1[21]);
  and and_a29_b22 (and_22[29], i0[29], i1[22]);
  and and_a29_b23 (and_23[29], i0[29], i1[23]);
  and and_a29_b24 (and_24[29], i0[29], i1[24]);
  and and_a29_b25 (and_25[29], i0[29], i1[25]);
  and and_a29_b26 (and_26[29], i0[29], i1[26]);
  and and_a29_b27 (and_27[29], i0[29], i1[27]);
  and and_a29_b28 (and_28[29], i0[29], i1[28]);
  and and_a29_b29 (and_29[29], i0[29], i1[29]);
  and and_a29_b3 (and_3[29], i0[29], i1[3]);
  and and_a29_b30 (and_30[29], i0[29], i1[30]);
  and and_a29_b31 (nand_31[29], i0[29], i1[31]);
  and and_a29_b4 (and_4[29], i0[29], i1[4]);
  and and_a29_b5 (and_5[29], i0[29], i1[5]);
  and and_a29_b6 (and_6[29], i0[29], i1[6]);
  and and_a29_b7 (and_7[29], i0[29], i1[7]);
  and and_a29_b8 (and_8[29], i0[29], i1[8]);
  and and_a29_b9 (and_9[29], i0[29], i1[9]);
  and and_a2_b0 (and_0[2], i0[2], i1[0]);
  and and_a2_b1 (and_1[2], i0[2], i1[1]);
  and and_a2_b10 (and_10[2], i0[2], i1[10]);
  and and_a2_b11 (and_11[2], i0[2], i1[11]);
  and and_a2_b12 (and_12[2], i0[2], i1[12]);
  and and_a2_b13 (and_13[2], i0[2], i1[13]);
  and and_a2_b14 (and_14[2], i0[2], i1[14]);
  and and_a2_b15 (and_15[2], i0[2], i1[15]);
  and and_a2_b16 (and_16[2], i0[2], i1[16]);
  and and_a2_b17 (and_17[2], i0[2], i1[17]);
  and and_a2_b18 (and_18[2], i0[2], i1[18]);
  and and_a2_b19 (and_19[2], i0[2], i1[19]);
  and and_a2_b2 (and_2[2], i0[2], i1[2]);
  and and_a2_b20 (and_20[2], i0[2], i1[20]);
  and and_a2_b21 (and_21[2], i0[2], i1[21]);
  and and_a2_b22 (and_22[2], i0[2], i1[22]);
  and and_a2_b23 (and_23[2], i0[2], i1[23]);
  and and_a2_b24 (and_24[2], i0[2], i1[24]);
  and and_a2_b25 (and_25[2], i0[2], i1[25]);
  and and_a2_b26 (and_26[2], i0[2], i1[26]);
  and and_a2_b27 (and_27[2], i0[2], i1[27]);
  and and_a2_b28 (and_28[2], i0[2], i1[28]);
  and and_a2_b29 (and_29[2], i0[2], i1[29]);
  and and_a2_b3 (and_3[2], i0[2], i1[3]);
  and and_a2_b30 (and_30[2], i0[2], i1[30]);
  and and_a2_b31 (nand_31[2], i0[2], i1[31]);
  and and_a2_b4 (and_4[2], i0[2], i1[4]);
  and and_a2_b5 (and_5[2], i0[2], i1[5]);
  and and_a2_b6 (and_6[2], i0[2], i1[6]);
  and and_a2_b7 (and_7[2], i0[2], i1[7]);
  and and_a2_b8 (and_8[2], i0[2], i1[8]);
  and and_a2_b9 (and_9[2], i0[2], i1[9]);
  and and_a30_b0 (and_0[30], i0[30], i1[0]);
  and and_a30_b1 (and_1[30], i0[30], i1[1]);
  and and_a30_b10 (and_10[30], i0[30], i1[10]);
  and and_a30_b11 (and_11[30], i0[30], i1[11]);
  and and_a30_b12 (and_12[30], i0[30], i1[12]);
  and and_a30_b13 (and_13[30], i0[30], i1[13]);
  and and_a30_b14 (and_14[30], i0[30], i1[14]);
  and and_a30_b15 (and_15[30], i0[30], i1[15]);
  and and_a30_b16 (and_16[30], i0[30], i1[16]);
  and and_a30_b17 (and_17[30], i0[30], i1[17]);
  and and_a30_b18 (and_18[30], i0[30], i1[18]);
  and and_a30_b19 (and_19[30], i0[30], i1[19]);
  and and_a30_b2 (and_2[30], i0[30], i1[2]);
  and and_a30_b20 (and_20[30], i0[30], i1[20]);
  and and_a30_b21 (and_21[30], i0[30], i1[21]);
  and and_a30_b22 (and_22[30], i0[30], i1[22]);
  and and_a30_b23 (and_23[30], i0[30], i1[23]);
  and and_a30_b24 (and_24[30], i0[30], i1[24]);
  and and_a30_b25 (and_25[30], i0[30], i1[25]);
  and and_a30_b26 (and_26[30], i0[30], i1[26]);
  and and_a30_b27 (and_27[30], i0[30], i1[27]);
  and and_a30_b28 (and_28[30], i0[30], i1[28]);
  and and_a30_b29 (and_29[30], i0[30], i1[29]);
  and and_a30_b3 (and_3[30], i0[30], i1[3]);
  and and_a30_b30 (and_30[30], i0[30], i1[30]);
  and and_a30_b31 (nand_31[30], i0[30], i1[31]);
  and and_a30_b4 (and_4[30], i0[30], i1[4]);
  and and_a30_b5 (and_5[30], i0[30], i1[5]);
  and and_a30_b6 (and_6[30], i0[30], i1[6]);
  and and_a30_b7 (and_7[30], i0[30], i1[7]);
  and and_a30_b8 (and_8[30], i0[30], i1[8]);
  and and_a30_b9 (and_9[30], i0[30], i1[9]);
  and and_a31_b0 (nand_0[31], i0[31], i1[0]);
  and and_a31_b1 (nand_1[31], i0[31], i1[1]);
  and and_a31_b10 (nand_10[31], i0[31], i1[10]);
  and and_a31_b11 (nand_11[31], i0[31], i1[11]);
  and and_a31_b12 (nand_12[31], i0[31], i1[12]);
  and and_a31_b13 (nand_13[31], i0[31], i1[13]);
  and and_a31_b14 (nand_14[31], i0[31], i1[14]);
  and and_a31_b15 (nand_15[31], i0[31], i1[15]);
  and and_a31_b16 (nand_16[31], i0[31], i1[16]);
  and and_a31_b17 (nand_17[31], i0[31], i1[17]);
  and and_a31_b18 (nand_18[31], i0[31], i1[18]);
  and and_a31_b19 (nand_19[31], i0[31], i1[19]);
  and and_a31_b2 (nand_2[31], i0[31], i1[2]);
  and and_a31_b20 (nand_20[31], i0[31], i1[20]);
  and and_a31_b21 (nand_21[31], i0[31], i1[21]);
  and and_a31_b22 (nand_22[31], i0[31], i1[22]);
  and and_a31_b23 (nand_23[31], i0[31], i1[23]);
  and and_a31_b24 (nand_24[31], i0[31], i1[24]);
  and and_a31_b25 (nand_25[31], i0[31], i1[25]);
  and and_a31_b26 (nand_26[31], i0[31], i1[26]);
  and and_a31_b27 (nand_27[31], i0[31], i1[27]);
  and and_a31_b28 (nand_28[31], i0[31], i1[28]);
  and and_a31_b29 (nand_29[31], i0[31], i1[29]);
  and and_a31_b3 (nand_3[31], i0[31], i1[3]);
  and and_a31_b30 (nand_30[31], i0[31], i1[30]);
  and and_a31_b31 (and_31[31], i0[31], i1[31]);
  and and_a31_b4 (nand_4[31], i0[31], i1[4]);
  and and_a31_b5 (nand_5[31], i0[31], i1[5]);
  and and_a31_b6 (nand_6[31], i0[31], i1[6]);
  and and_a31_b7 (nand_7[31], i0[31], i1[7]);
  and and_a31_b8 (nand_8[31], i0[31], i1[8]);
  and and_a31_b9 (nand_9[31], i0[31], i1[9]);
  and and_a3_b0 (and_0[3], i0[3], i1[0]);
  and and_a3_b1 (and_1[3], i0[3], i1[1]);
  and and_a3_b10 (and_10[3], i0[3], i1[10]);
  and and_a3_b11 (and_11[3], i0[3], i1[11]);
  and and_a3_b12 (and_12[3], i0[3], i1[12]);
  and and_a3_b13 (and_13[3], i0[3], i1[13]);
  and and_a3_b14 (and_14[3], i0[3], i1[14]);
  and and_a3_b15 (and_15[3], i0[3], i1[15]);
  and and_a3_b16 (and_16[3], i0[3], i1[16]);
  and and_a3_b17 (and_17[3], i0[3], i1[17]);
  and and_a3_b18 (and_18[3], i0[3], i1[18]);
  and and_a3_b19 (and_19[3], i0[3], i1[19]);
  and and_a3_b2 (and_2[3], i0[3], i1[2]);
  and and_a3_b20 (and_20[3], i0[3], i1[20]);
  and and_a3_b21 (and_21[3], i0[3], i1[21]);
  and and_a3_b22 (and_22[3], i0[3], i1[22]);
  and and_a3_b23 (and_23[3], i0[3], i1[23]);
  and and_a3_b24 (and_24[3], i0[3], i1[24]);
  and and_a3_b25 (and_25[3], i0[3], i1[25]);
  and and_a3_b26 (and_26[3], i0[3], i1[26]);
  and and_a3_b27 (and_27[3], i0[3], i1[27]);
  and and_a3_b28 (and_28[3], i0[3], i1[28]);
  and and_a3_b29 (and_29[3], i0[3], i1[29]);
  and and_a3_b3 (and_3[3], i0[3], i1[3]);
  and and_a3_b30 (and_30[3], i0[3], i1[30]);
  and and_a3_b31 (nand_31[3], i0[3], i1[31]);
  and and_a3_b4 (and_4[3], i0[3], i1[4]);
  and and_a3_b5 (and_5[3], i0[3], i1[5]);
  and and_a3_b6 (and_6[3], i0[3], i1[6]);
  and and_a3_b7 (and_7[3], i0[3], i1[7]);
  and and_a3_b8 (and_8[3], i0[3], i1[8]);
  and and_a3_b9 (and_9[3], i0[3], i1[9]);
  and and_a4_b0 (and_0[4], i0[4], i1[0]);
  and and_a4_b1 (and_1[4], i0[4], i1[1]);
  and and_a4_b10 (and_10[4], i0[4], i1[10]);
  and and_a4_b11 (and_11[4], i0[4], i1[11]);
  and and_a4_b12 (and_12[4], i0[4], i1[12]);
  and and_a4_b13 (and_13[4], i0[4], i1[13]);
  and and_a4_b14 (and_14[4], i0[4], i1[14]);
  and and_a4_b15 (and_15[4], i0[4], i1[15]);
  and and_a4_b16 (and_16[4], i0[4], i1[16]);
  and and_a4_b17 (and_17[4], i0[4], i1[17]);
  and and_a4_b18 (and_18[4], i0[4], i1[18]);
  and and_a4_b19 (and_19[4], i0[4], i1[19]);
  and and_a4_b2 (and_2[4], i0[4], i1[2]);
  and and_a4_b20 (and_20[4], i0[4], i1[20]);
  and and_a4_b21 (and_21[4], i0[4], i1[21]);
  and and_a4_b22 (and_22[4], i0[4], i1[22]);
  and and_a4_b23 (and_23[4], i0[4], i1[23]);
  and and_a4_b24 (and_24[4], i0[4], i1[24]);
  and and_a4_b25 (and_25[4], i0[4], i1[25]);
  and and_a4_b26 (and_26[4], i0[4], i1[26]);
  and and_a4_b27 (and_27[4], i0[4], i1[27]);
  and and_a4_b28 (and_28[4], i0[4], i1[28]);
  and and_a4_b29 (and_29[4], i0[4], i1[29]);
  and and_a4_b3 (and_3[4], i0[4], i1[3]);
  and and_a4_b30 (and_30[4], i0[4], i1[30]);
  and and_a4_b31 (nand_31[4], i0[4], i1[31]);
  and and_a4_b4 (and_4[4], i0[4], i1[4]);
  and and_a4_b5 (and_5[4], i0[4], i1[5]);
  and and_a4_b6 (and_6[4], i0[4], i1[6]);
  and and_a4_b7 (and_7[4], i0[4], i1[7]);
  and and_a4_b8 (and_8[4], i0[4], i1[8]);
  and and_a4_b9 (and_9[4], i0[4], i1[9]);
  and and_a5_b0 (and_0[5], i0[5], i1[0]);
  and and_a5_b1 (and_1[5], i0[5], i1[1]);
  and and_a5_b10 (and_10[5], i0[5], i1[10]);
  and and_a5_b11 (and_11[5], i0[5], i1[11]);
  and and_a5_b12 (and_12[5], i0[5], i1[12]);
  and and_a5_b13 (and_13[5], i0[5], i1[13]);
  and and_a5_b14 (and_14[5], i0[5], i1[14]);
  and and_a5_b15 (and_15[5], i0[5], i1[15]);
  and and_a5_b16 (and_16[5], i0[5], i1[16]);
  and and_a5_b17 (and_17[5], i0[5], i1[17]);
  and and_a5_b18 (and_18[5], i0[5], i1[18]);
  and and_a5_b19 (and_19[5], i0[5], i1[19]);
  and and_a5_b2 (and_2[5], i0[5], i1[2]);
  and and_a5_b20 (and_20[5], i0[5], i1[20]);
  and and_a5_b21 (and_21[5], i0[5], i1[21]);
  and and_a5_b22 (and_22[5], i0[5], i1[22]);
  and and_a5_b23 (and_23[5], i0[5], i1[23]);
  and and_a5_b24 (and_24[5], i0[5], i1[24]);
  and and_a5_b25 (and_25[5], i0[5], i1[25]);
  and and_a5_b26 (and_26[5], i0[5], i1[26]);
  and and_a5_b27 (and_27[5], i0[5], i1[27]);
  and and_a5_b28 (and_28[5], i0[5], i1[28]);
  and and_a5_b29 (and_29[5], i0[5], i1[29]);
  and and_a5_b3 (and_3[5], i0[5], i1[3]);
  and and_a5_b30 (and_30[5], i0[5], i1[30]);
  and and_a5_b31 (nand_31[5], i0[5], i1[31]);
  and and_a5_b4 (and_4[5], i0[5], i1[4]);
  and and_a5_b5 (and_5[5], i0[5], i1[5]);
  and and_a5_b6 (and_6[5], i0[5], i1[6]);
  and and_a5_b7 (and_7[5], i0[5], i1[7]);
  and and_a5_b8 (and_8[5], i0[5], i1[8]);
  and and_a5_b9 (and_9[5], i0[5], i1[9]);
  and and_a6_b0 (and_0[6], i0[6], i1[0]);
  and and_a6_b1 (and_1[6], i0[6], i1[1]);
  and and_a6_b10 (and_10[6], i0[6], i1[10]);
  and and_a6_b11 (and_11[6], i0[6], i1[11]);
  and and_a6_b12 (and_12[6], i0[6], i1[12]);
  and and_a6_b13 (and_13[6], i0[6], i1[13]);
  and and_a6_b14 (and_14[6], i0[6], i1[14]);
  and and_a6_b15 (and_15[6], i0[6], i1[15]);
  and and_a6_b16 (and_16[6], i0[6], i1[16]);
  and and_a6_b17 (and_17[6], i0[6], i1[17]);
  and and_a6_b18 (and_18[6], i0[6], i1[18]);
  and and_a6_b19 (and_19[6], i0[6], i1[19]);
  and and_a6_b2 (and_2[6], i0[6], i1[2]);
  and and_a6_b20 (and_20[6], i0[6], i1[20]);
  and and_a6_b21 (and_21[6], i0[6], i1[21]);
  and and_a6_b22 (and_22[6], i0[6], i1[22]);
  and and_a6_b23 (and_23[6], i0[6], i1[23]);
  and and_a6_b24 (and_24[6], i0[6], i1[24]);
  and and_a6_b25 (and_25[6], i0[6], i1[25]);
  and and_a6_b26 (and_26[6], i0[6], i1[26]);
  and and_a6_b27 (and_27[6], i0[6], i1[27]);
  and and_a6_b28 (and_28[6], i0[6], i1[28]);
  and and_a6_b29 (and_29[6], i0[6], i1[29]);
  and and_a6_b3 (and_3[6], i0[6], i1[3]);
  and and_a6_b30 (and_30[6], i0[6], i1[30]);
  and and_a6_b31 (nand_31[6], i0[6], i1[31]);
  and and_a6_b4 (and_4[6], i0[6], i1[4]);
  and and_a6_b5 (and_5[6], i0[6], i1[5]);
  and and_a6_b6 (and_6[6], i0[6], i1[6]);
  and and_a6_b7 (and_7[6], i0[6], i1[7]);
  and and_a6_b8 (and_8[6], i0[6], i1[8]);
  and and_a6_b9 (and_9[6], i0[6], i1[9]);
  and and_a7_b0 (and_0[7], i0[7], i1[0]);
  and and_a7_b1 (and_1[7], i0[7], i1[1]);
  and and_a7_b10 (and_10[7], i0[7], i1[10]);
  and and_a7_b11 (and_11[7], i0[7], i1[11]);
  and and_a7_b12 (and_12[7], i0[7], i1[12]);
  and and_a7_b13 (and_13[7], i0[7], i1[13]);
  and and_a7_b14 (and_14[7], i0[7], i1[14]);
  and and_a7_b15 (and_15[7], i0[7], i1[15]);
  and and_a7_b16 (and_16[7], i0[7], i1[16]);
  and and_a7_b17 (and_17[7], i0[7], i1[17]);
  and and_a7_b18 (and_18[7], i0[7], i1[18]);
  and and_a7_b19 (and_19[7], i0[7], i1[19]);
  and and_a7_b2 (and_2[7], i0[7], i1[2]);
  and and_a7_b20 (and_20[7], i0[7], i1[20]);
  and and_a7_b21 (and_21[7], i0[7], i1[21]);
  and and_a7_b22 (and_22[7], i0[7], i1[22]);
  and and_a7_b23 (and_23[7], i0[7], i1[23]);
  and and_a7_b24 (and_24[7], i0[7], i1[24]);
  and and_a7_b25 (and_25[7], i0[7], i1[25]);
  and and_a7_b26 (and_26[7], i0[7], i1[26]);
  and and_a7_b27 (and_27[7], i0[7], i1[27]);
  and and_a7_b28 (and_28[7], i0[7], i1[28]);
  and and_a7_b29 (and_29[7], i0[7], i1[29]);
  and and_a7_b3 (and_3[7], i0[7], i1[3]);
  and and_a7_b30 (and_30[7], i0[7], i1[30]);
  and and_a7_b31 (nand_31[7], i0[7], i1[31]);
  and and_a7_b4 (and_4[7], i0[7], i1[4]);
  and and_a7_b5 (and_5[7], i0[7], i1[5]);
  and and_a7_b6 (and_6[7], i0[7], i1[6]);
  and and_a7_b7 (and_7[7], i0[7], i1[7]);
  and and_a7_b8 (and_8[7], i0[7], i1[8]);
  and and_a7_b9 (and_9[7], i0[7], i1[9]);
  and and_a8_b0 (and_0[8], i0[8], i1[0]);
  and and_a8_b1 (and_1[8], i0[8], i1[1]);
  and and_a8_b10 (and_10[8], i0[8], i1[10]);
  and and_a8_b11 (and_11[8], i0[8], i1[11]);
  and and_a8_b12 (and_12[8], i0[8], i1[12]);
  and and_a8_b13 (and_13[8], i0[8], i1[13]);
  and and_a8_b14 (and_14[8], i0[8], i1[14]);
  and and_a8_b15 (and_15[8], i0[8], i1[15]);
  and and_a8_b16 (and_16[8], i0[8], i1[16]);
  and and_a8_b17 (and_17[8], i0[8], i1[17]);
  and and_a8_b18 (and_18[8], i0[8], i1[18]);
  and and_a8_b19 (and_19[8], i0[8], i1[19]);
  and and_a8_b2 (and_2[8], i0[8], i1[2]);
  and and_a8_b20 (and_20[8], i0[8], i1[20]);
  and and_a8_b21 (and_21[8], i0[8], i1[21]);
  and and_a8_b22 (and_22[8], i0[8], i1[22]);
  and and_a8_b23 (and_23[8], i0[8], i1[23]);
  and and_a8_b24 (and_24[8], i0[8], i1[24]);
  and and_a8_b25 (and_25[8], i0[8], i1[25]);
  and and_a8_b26 (and_26[8], i0[8], i1[26]);
  and and_a8_b27 (and_27[8], i0[8], i1[27]);
  and and_a8_b28 (and_28[8], i0[8], i1[28]);
  and and_a8_b29 (and_29[8], i0[8], i1[29]);
  and and_a8_b3 (and_3[8], i0[8], i1[3]);
  and and_a8_b30 (and_30[8], i0[8], i1[30]);
  and and_a8_b31 (nand_31[8], i0[8], i1[31]);
  and and_a8_b4 (and_4[8], i0[8], i1[4]);
  and and_a8_b5 (and_5[8], i0[8], i1[5]);
  and and_a8_b6 (and_6[8], i0[8], i1[6]);
  and and_a8_b7 (and_7[8], i0[8], i1[7]);
  and and_a8_b8 (and_8[8], i0[8], i1[8]);
  and and_a8_b9 (and_9[8], i0[8], i1[9]);
  and and_a9_b0 (and_0[9], i0[9], i1[0]);
  and and_a9_b1 (and_1[9], i0[9], i1[1]);
  and and_a9_b10 (and_10[9], i0[9], i1[10]);
  and and_a9_b11 (and_11[9], i0[9], i1[11]);
  and and_a9_b12 (and_12[9], i0[9], i1[12]);
  and and_a9_b13 (and_13[9], i0[9], i1[13]);
  and and_a9_b14 (and_14[9], i0[9], i1[14]);
  and and_a9_b15 (and_15[9], i0[9], i1[15]);
  and and_a9_b16 (and_16[9], i0[9], i1[16]);
  and and_a9_b17 (and_17[9], i0[9], i1[17]);
  and and_a9_b18 (and_18[9], i0[9], i1[18]);
  and and_a9_b19 (and_19[9], i0[9], i1[19]);
  and and_a9_b2 (and_2[9], i0[9], i1[2]);
  and and_a9_b20 (and_20[9], i0[9], i1[20]);
  and and_a9_b21 (and_21[9], i0[9], i1[21]);
  and and_a9_b22 (and_22[9], i0[9], i1[22]);
  and and_a9_b23 (and_23[9], i0[9], i1[23]);
  and and_a9_b24 (and_24[9], i0[9], i1[24]);
  and and_a9_b25 (and_25[9], i0[9], i1[25]);
  and and_a9_b26 (and_26[9], i0[9], i1[26]);
  and and_a9_b27 (and_27[9], i0[9], i1[27]);
  and and_a9_b28 (and_28[9], i0[9], i1[28]);
  and and_a9_b29 (and_29[9], i0[9], i1[29]);
  and and_a9_b3 (and_3[9], i0[9], i1[3]);
  and and_a9_b30 (and_30[9], i0[9], i1[30]);
  and and_a9_b31 (nand_31[9], i0[9], i1[31]);
  and and_a9_b4 (and_4[9], i0[9], i1[4]);
  and and_a9_b5 (and_5[9], i0[9], i1[5]);
  and and_a9_b6 (and_6[9], i0[9], i1[6]);
  and and_a9_b7 (and_7[9], i0[9], i1[7]);
  and and_a9_b8 (and_8[9], i0[9], i1[8]);
  and and_a9_b9 (and_9[9], i0[9], i1[9]);
  add_pu63_pu60_pu59_pu58_pu57_pu56_pu55_pu54_pu53_pu52_pu51_pu50_pu49_pu48_pu47_pu46_pu45_pu44_pu43_pu42_pu41_pu40_pu39_pu38_pu37_pu36_pu35_pu34_pu33_pu32_pu31_mu62_mu62_o64 sum (
    .i0({and_31[31],1'b0,and_30[30],and_29[30],and_28[30],and_27[30],and_26[30],and_25[30],and_24[30],and_23[30],and_22[30],and_21[30],and_20[30],and_19[30],and_18[30],and_17[30],and_16[30],and_15[30],and_14[30],and_13[30],and_12[30],and_11[30],and_10[30],and_9[30],and_8[30],and_7[30],and_6[30],and_5[30],and_4[30],and_3[30],and_2[30],and_1[30],and_0[30:0]}),
    .i1({and_30[29],and_29[29],and_28[29],and_27[29],and_26[29],and_25[29],and_24[29],and_23[29],and_22[29],and_21[29],and_20[29],and_19[29],and_18[29],and_17[29],and_16[29],and_15[29],and_14[29],and_13[29],and_12[29],and_11[29],and_10[29],and_9[29],and_8[29],and_7[29],and_6[29],and_5[29],and_4[29],and_3[29],and_2[29],and_1[29:0],1'b0}),
    .i10({and_30[20],and_29[20],and_28[20],and_27[20],and_26[20],and_25[20],and_24[20],and_23[20],and_22[20],and_21[20],and_20[20],and_19[20],and_18[20],and_17[20],and_16[20],and_15[20],and_14[20],and_13[20],and_12[20],and_11[20],and_10[20:0],10'b0000000000}),
    .i11({and_30[19],and_29[19],and_28[19],and_27[19],and_26[19],and_25[19],and_24[19],and_23[19],and_22[19],and_21[19],and_20[19],and_19[19],and_18[19],and_17[19],and_16[19],and_15[19],and_14[19],and_13[19],and_12[19],and_11[19:0],11'b00000000000}),
    .i12({and_30[18],and_29[18],and_28[18],and_27[18],and_26[18],and_25[18],and_24[18],and_23[18],and_22[18],and_21[18],and_20[18],and_19[18],and_18[18],and_17[18],and_16[18],and_15[18],and_14[18],and_13[18],and_12[18:0],12'b000000000000}),
    .i13({and_30[17],and_29[17],and_28[17],and_27[17],and_26[17],and_25[17],and_24[17],and_23[17],and_22[17],and_21[17],and_20[17],and_19[17],and_18[17],and_17[17],and_16[17],and_15[17],and_14[17],and_13[17:0],13'b0000000000000}),
    .i14({and_30[16],and_29[16],and_28[16],and_27[16],and_26[16],and_25[16],and_24[16],and_23[16],and_22[16],and_21[16],and_20[16],and_19[16],and_18[16],and_17[16],and_16[16],and_15[16],and_14[16:0],14'b00000000000000}),
    .i15({and_30[15],and_29[15],and_28[15],and_27[15],and_26[15],and_25[15],and_24[15],and_23[15],and_22[15],and_21[15],and_20[15],and_19[15],and_18[15],and_17[15],and_16[15],and_15[15:0],15'b000000000000000}),
    .i16({and_30[14],and_29[14],and_28[14],and_27[14],and_26[14],and_25[14],and_24[14],and_23[14],and_22[14],and_21[14],and_20[14],and_19[14],and_18[14],and_17[14],and_16[14:0],16'b0000000000000000}),
    .i17({and_30[13],and_29[13],and_28[13],and_27[13],and_26[13],and_25[13],and_24[13],and_23[13],and_22[13],and_21[13],and_20[13],and_19[13],and_18[13],and_17[13:0],17'b00000000000000000}),
    .i18({and_30[12],and_29[12],and_28[12],and_27[12],and_26[12],and_25[12],and_24[12],and_23[12],and_22[12],and_21[12],and_20[12],and_19[12],and_18[12:0],18'b000000000000000000}),
    .i19({and_30[11],and_29[11],and_28[11],and_27[11],and_26[11],and_25[11],and_24[11],and_23[11],and_22[11],and_21[11],and_20[11],and_19[11:0],19'b0000000000000000000}),
    .i2({and_30[28],and_29[28],and_28[28],and_27[28],and_26[28],and_25[28],and_24[28],and_23[28],and_22[28],and_21[28],and_20[28],and_19[28],and_18[28],and_17[28],and_16[28],and_15[28],and_14[28],and_13[28],and_12[28],and_11[28],and_10[28],and_9[28],and_8[28],and_7[28],and_6[28],and_5[28],and_4[28],and_3[28],and_2[28:0],2'b00}),
    .i20({and_30[10],and_29[10],and_28[10],and_27[10],and_26[10],and_25[10],and_24[10],and_23[10],and_22[10],and_21[10],and_20[10:0],20'b00000000000000000000}),
    .i21({and_30[9],and_29[9],and_28[9],and_27[9],and_26[9],and_25[9],and_24[9],and_23[9],and_22[9],and_21[9:0],21'b000000000000000000000}),
    .i22({and_30[8],and_29[8],and_28[8],and_27[8],and_26[8],and_25[8],and_24[8],and_23[8],and_22[8:0],22'b0000000000000000000000}),
    .i23({and_30[7],and_29[7],and_28[7],and_27[7],and_26[7],and_25[7],and_24[7],and_23[7:0],23'b00000000000000000000000}),
    .i24({and_30[6],and_29[6],and_28[6],and_27[6],and_26[6],and_25[6],and_24[6:0],24'b000000000000000000000000}),
    .i25({and_30[5],and_29[5],and_28[5],and_27[5],and_26[5],and_25[5:0],25'b0000000000000000000000000}),
    .i26({and_30[4],and_29[4],and_28[4],and_27[4],and_26[4:0],26'b00000000000000000000000000}),
    .i27({and_30[3],and_29[3],and_28[3],and_27[3:0],27'b000000000000000000000000000}),
    .i28({and_30[2],and_29[2],and_28[2:0],28'b0000000000000000000000000000}),
    .i29({and_30[1],and_29[1:0],29'b00000000000000000000000000000}),
    .i3({and_30[27],and_29[27],and_28[27],and_27[27],and_26[27],and_25[27],and_24[27],and_23[27],and_22[27],and_21[27],and_20[27],and_19[27],and_18[27],and_17[27],and_16[27],and_15[27],and_14[27],and_13[27],and_12[27],and_11[27],and_10[27],and_9[27],and_8[27],and_7[27],and_6[27],and_5[27],and_4[27],and_3[27:0],3'b000}),
    .i30({and_30[0],30'b000000000000000000000000000000}),
    .i31({nand_30[31],nand_29[31],nand_28[31],nand_27[31],nand_26[31],nand_25[31],nand_24[31],nand_23[31],nand_22[31],nand_21[31],nand_20[31],nand_19[31],nand_18[31],nand_17[31],nand_16[31],nand_15[31],nand_14[31],nand_13[31],nand_12[31],nand_11[31],nand_10[31],nand_9[31],nand_8[31],nand_7[31],nand_6[31],nand_5[31],nand_4[31],nand_3[31],nand_2[31],nand_1[31],nand_0[31],31'b0000000000000000000000000000000}),
    .i32({nand_31[30:0],31'b0000000000000000000000000000000}),
    .i4({and_30[26],and_29[26],and_28[26],and_27[26],and_26[26],and_25[26],and_24[26],and_23[26],and_22[26],and_21[26],and_20[26],and_19[26],and_18[26],and_17[26],and_16[26],and_15[26],and_14[26],and_13[26],and_12[26],and_11[26],and_10[26],and_9[26],and_8[26],and_7[26],and_6[26],and_5[26],and_4[26:0],4'b0000}),
    .i5({and_30[25],and_29[25],and_28[25],and_27[25],and_26[25],and_25[25],and_24[25],and_23[25],and_22[25],and_21[25],and_20[25],and_19[25],and_18[25],and_17[25],and_16[25],and_15[25],and_14[25],and_13[25],and_12[25],and_11[25],and_10[25],and_9[25],and_8[25],and_7[25],and_6[25],and_5[25:0],5'b00000}),
    .i6({and_30[24],and_29[24],and_28[24],and_27[24],and_26[24],and_25[24],and_24[24],and_23[24],and_22[24],and_21[24],and_20[24],and_19[24],and_18[24],and_17[24],and_16[24],and_15[24],and_14[24],and_13[24],and_12[24],and_11[24],and_10[24],and_9[24],and_8[24],and_7[24],and_6[24:0],6'b000000}),
    .i7({and_30[23],and_29[23],and_28[23],and_27[23],and_26[23],and_25[23],and_24[23],and_23[23],and_22[23],and_21[23],and_20[23],and_19[23],and_18[23],and_17[23],and_16[23],and_15[23],and_14[23],and_13[23],and_12[23],and_11[23],and_10[23],and_9[23],and_8[23],and_7[23:0],7'b0000000}),
    .i8({and_30[22],and_29[22],and_28[22],and_27[22],and_26[22],and_25[22],and_24[22],and_23[22],and_22[22],and_21[22],and_20[22],and_19[22],and_18[22],and_17[22],and_16[22],and_15[22],and_14[22],and_13[22],and_12[22],and_11[22],and_10[22],and_9[22],and_8[22:0],8'b00000000}),
    .i9({and_30[21],and_29[21],and_28[21],and_27[21],and_26[21],and_25[21],and_24[21],and_23[21],and_22[21],and_21[21],and_20[21],and_19[21],and_18[21],and_17[21],and_16[21],and_15[21],and_14[21],and_13[21],and_12[21],and_11[21],and_10[21],and_9[21:0],9'b000000000}),
    .o(o));

endmodule 

module mult_u32_u32_o64
  (
  i0,
  i1,
  o
  );

  input [31:0] i0;
  input [31:0] i1;
  output [63:0] o;

  wire [31:0] and_0;
  wire [31:0] and_1;
  wire [31:0] and_10;
  wire [31:0] and_11;
  wire [31:0] and_12;
  wire [31:0] and_13;
  wire [31:0] and_14;
  wire [31:0] and_15;
  wire [31:0] and_16;
  wire [31:0] and_17;
  wire [31:0] and_18;
  wire [31:0] and_19;
  wire [31:0] and_2;
  wire [31:0] and_20;
  wire [31:0] and_21;
  wire [31:0] and_22;
  wire [31:0] and_23;
  wire [31:0] and_24;
  wire [31:0] and_25;
  wire [31:0] and_26;
  wire [31:0] and_27;
  wire [31:0] and_28;
  wire [31:0] and_29;
  wire [31:0] and_3;
  wire [31:0] and_30;
  wire [31:0] and_31;
  wire [31:0] and_4;
  wire [31:0] and_5;
  wire [31:0] and_6;
  wire [31:0] and_7;
  wire [31:0] and_8;
  wire [31:0] and_9;
  wire [31:0] nand_0;
  wire [31:0] nand_1;
  wire [31:0] nand_10;
  wire [31:0] nand_11;
  wire [31:0] nand_12;
  wire [31:0] nand_13;
  wire [31:0] nand_14;
  wire [31:0] nand_15;
  wire [31:0] nand_16;
  wire [31:0] nand_17;
  wire [31:0] nand_18;
  wire [31:0] nand_19;
  wire [31:0] nand_2;
  wire [31:0] nand_20;
  wire [31:0] nand_21;
  wire [31:0] nand_22;
  wire [31:0] nand_23;
  wire [31:0] nand_24;
  wire [31:0] nand_25;
  wire [31:0] nand_26;
  wire [31:0] nand_27;
  wire [31:0] nand_28;
  wire [31:0] nand_29;
  wire [31:0] nand_3;
  wire [31:0] nand_30;
  wire [31:0] nand_31;
  wire [31:0] nand_4;
  wire [31:0] nand_5;
  wire [31:0] nand_6;
  wire [31:0] nand_7;
  wire [31:0] nand_8;
  wire [31:0] nand_9;

  and and_a0_b0 (and_0[0], i0[0], i1[0]);
  and and_a0_b1 (and_1[0], i0[0], i1[1]);
  and and_a0_b10 (and_10[0], i0[0], i1[10]);
  and and_a0_b11 (and_11[0], i0[0], i1[11]);
  and and_a0_b12 (and_12[0], i0[0], i1[12]);
  and and_a0_b13 (and_13[0], i0[0], i1[13]);
  and and_a0_b14 (and_14[0], i0[0], i1[14]);
  and and_a0_b15 (and_15[0], i0[0], i1[15]);
  and and_a0_b16 (and_16[0], i0[0], i1[16]);
  and and_a0_b17 (and_17[0], i0[0], i1[17]);
  and and_a0_b18 (and_18[0], i0[0], i1[18]);
  and and_a0_b19 (and_19[0], i0[0], i1[19]);
  and and_a0_b2 (and_2[0], i0[0], i1[2]);
  and and_a0_b20 (and_20[0], i0[0], i1[20]);
  and and_a0_b21 (and_21[0], i0[0], i1[21]);
  and and_a0_b22 (and_22[0], i0[0], i1[22]);
  and and_a0_b23 (and_23[0], i0[0], i1[23]);
  and and_a0_b24 (and_24[0], i0[0], i1[24]);
  and and_a0_b25 (and_25[0], i0[0], i1[25]);
  and and_a0_b26 (and_26[0], i0[0], i1[26]);
  and and_a0_b27 (and_27[0], i0[0], i1[27]);
  and and_a0_b28 (and_28[0], i0[0], i1[28]);
  and and_a0_b29 (and_29[0], i0[0], i1[29]);
  and and_a0_b3 (and_3[0], i0[0], i1[3]);
  and and_a0_b30 (and_30[0], i0[0], i1[30]);
  and and_a0_b31 (and_31[0], i0[0], i1[31]);
  and and_a0_b4 (and_4[0], i0[0], i1[4]);
  and and_a0_b5 (and_5[0], i0[0], i1[5]);
  and and_a0_b6 (and_6[0], i0[0], i1[6]);
  and and_a0_b7 (and_7[0], i0[0], i1[7]);
  and and_a0_b8 (and_8[0], i0[0], i1[8]);
  and and_a0_b9 (and_9[0], i0[0], i1[9]);
  and and_a10_b0 (and_0[10], i0[10], i1[0]);
  and and_a10_b1 (and_1[10], i0[10], i1[1]);
  and and_a10_b10 (and_10[10], i0[10], i1[10]);
  and and_a10_b11 (and_11[10], i0[10], i1[11]);
  and and_a10_b12 (and_12[10], i0[10], i1[12]);
  and and_a10_b13 (and_13[10], i0[10], i1[13]);
  and and_a10_b14 (and_14[10], i0[10], i1[14]);
  and and_a10_b15 (and_15[10], i0[10], i1[15]);
  and and_a10_b16 (and_16[10], i0[10], i1[16]);
  and and_a10_b17 (and_17[10], i0[10], i1[17]);
  and and_a10_b18 (and_18[10], i0[10], i1[18]);
  and and_a10_b19 (and_19[10], i0[10], i1[19]);
  and and_a10_b2 (and_2[10], i0[10], i1[2]);
  and and_a10_b20 (and_20[10], i0[10], i1[20]);
  and and_a10_b21 (and_21[10], i0[10], i1[21]);
  and and_a10_b22 (and_22[10], i0[10], i1[22]);
  and and_a10_b23 (and_23[10], i0[10], i1[23]);
  and and_a10_b24 (and_24[10], i0[10], i1[24]);
  and and_a10_b25 (and_25[10], i0[10], i1[25]);
  and and_a10_b26 (and_26[10], i0[10], i1[26]);
  and and_a10_b27 (and_27[10], i0[10], i1[27]);
  and and_a10_b28 (and_28[10], i0[10], i1[28]);
  and and_a10_b29 (and_29[10], i0[10], i1[29]);
  and and_a10_b3 (and_3[10], i0[10], i1[3]);
  and and_a10_b30 (and_30[10], i0[10], i1[30]);
  and and_a10_b31 (and_31[10], i0[10], i1[31]);
  and and_a10_b4 (and_4[10], i0[10], i1[4]);
  and and_a10_b5 (and_5[10], i0[10], i1[5]);
  and and_a10_b6 (and_6[10], i0[10], i1[6]);
  and and_a10_b7 (and_7[10], i0[10], i1[7]);
  and and_a10_b8 (and_8[10], i0[10], i1[8]);
  and and_a10_b9 (and_9[10], i0[10], i1[9]);
  and and_a11_b0 (and_0[11], i0[11], i1[0]);
  and and_a11_b1 (and_1[11], i0[11], i1[1]);
  and and_a11_b10 (and_10[11], i0[11], i1[10]);
  and and_a11_b11 (and_11[11], i0[11], i1[11]);
  and and_a11_b12 (and_12[11], i0[11], i1[12]);
  and and_a11_b13 (and_13[11], i0[11], i1[13]);
  and and_a11_b14 (and_14[11], i0[11], i1[14]);
  and and_a11_b15 (and_15[11], i0[11], i1[15]);
  and and_a11_b16 (and_16[11], i0[11], i1[16]);
  and and_a11_b17 (and_17[11], i0[11], i1[17]);
  and and_a11_b18 (and_18[11], i0[11], i1[18]);
  and and_a11_b19 (and_19[11], i0[11], i1[19]);
  and and_a11_b2 (and_2[11], i0[11], i1[2]);
  and and_a11_b20 (and_20[11], i0[11], i1[20]);
  and and_a11_b21 (and_21[11], i0[11], i1[21]);
  and and_a11_b22 (and_22[11], i0[11], i1[22]);
  and and_a11_b23 (and_23[11], i0[11], i1[23]);
  and and_a11_b24 (and_24[11], i0[11], i1[24]);
  and and_a11_b25 (and_25[11], i0[11], i1[25]);
  and and_a11_b26 (and_26[11], i0[11], i1[26]);
  and and_a11_b27 (and_27[11], i0[11], i1[27]);
  and and_a11_b28 (and_28[11], i0[11], i1[28]);
  and and_a11_b29 (and_29[11], i0[11], i1[29]);
  and and_a11_b3 (and_3[11], i0[11], i1[3]);
  and and_a11_b30 (and_30[11], i0[11], i1[30]);
  and and_a11_b31 (and_31[11], i0[11], i1[31]);
  and and_a11_b4 (and_4[11], i0[11], i1[4]);
  and and_a11_b5 (and_5[11], i0[11], i1[5]);
  and and_a11_b6 (and_6[11], i0[11], i1[6]);
  and and_a11_b7 (and_7[11], i0[11], i1[7]);
  and and_a11_b8 (and_8[11], i0[11], i1[8]);
  and and_a11_b9 (and_9[11], i0[11], i1[9]);
  and and_a12_b0 (and_0[12], i0[12], i1[0]);
  and and_a12_b1 (and_1[12], i0[12], i1[1]);
  and and_a12_b10 (and_10[12], i0[12], i1[10]);
  and and_a12_b11 (and_11[12], i0[12], i1[11]);
  and and_a12_b12 (and_12[12], i0[12], i1[12]);
  and and_a12_b13 (and_13[12], i0[12], i1[13]);
  and and_a12_b14 (and_14[12], i0[12], i1[14]);
  and and_a12_b15 (and_15[12], i0[12], i1[15]);
  and and_a12_b16 (and_16[12], i0[12], i1[16]);
  and and_a12_b17 (and_17[12], i0[12], i1[17]);
  and and_a12_b18 (and_18[12], i0[12], i1[18]);
  and and_a12_b19 (and_19[12], i0[12], i1[19]);
  and and_a12_b2 (and_2[12], i0[12], i1[2]);
  and and_a12_b20 (and_20[12], i0[12], i1[20]);
  and and_a12_b21 (and_21[12], i0[12], i1[21]);
  and and_a12_b22 (and_22[12], i0[12], i1[22]);
  and and_a12_b23 (and_23[12], i0[12], i1[23]);
  and and_a12_b24 (and_24[12], i0[12], i1[24]);
  and and_a12_b25 (and_25[12], i0[12], i1[25]);
  and and_a12_b26 (and_26[12], i0[12], i1[26]);
  and and_a12_b27 (and_27[12], i0[12], i1[27]);
  and and_a12_b28 (and_28[12], i0[12], i1[28]);
  and and_a12_b29 (and_29[12], i0[12], i1[29]);
  and and_a12_b3 (and_3[12], i0[12], i1[3]);
  and and_a12_b30 (and_30[12], i0[12], i1[30]);
  and and_a12_b31 (and_31[12], i0[12], i1[31]);
  and and_a12_b4 (and_4[12], i0[12], i1[4]);
  and and_a12_b5 (and_5[12], i0[12], i1[5]);
  and and_a12_b6 (and_6[12], i0[12], i1[6]);
  and and_a12_b7 (and_7[12], i0[12], i1[7]);
  and and_a12_b8 (and_8[12], i0[12], i1[8]);
  and and_a12_b9 (and_9[12], i0[12], i1[9]);
  and and_a13_b0 (and_0[13], i0[13], i1[0]);
  and and_a13_b1 (and_1[13], i0[13], i1[1]);
  and and_a13_b10 (and_10[13], i0[13], i1[10]);
  and and_a13_b11 (and_11[13], i0[13], i1[11]);
  and and_a13_b12 (and_12[13], i0[13], i1[12]);
  and and_a13_b13 (and_13[13], i0[13], i1[13]);
  and and_a13_b14 (and_14[13], i0[13], i1[14]);
  and and_a13_b15 (and_15[13], i0[13], i1[15]);
  and and_a13_b16 (and_16[13], i0[13], i1[16]);
  and and_a13_b17 (and_17[13], i0[13], i1[17]);
  and and_a13_b18 (and_18[13], i0[13], i1[18]);
  and and_a13_b19 (and_19[13], i0[13], i1[19]);
  and and_a13_b2 (and_2[13], i0[13], i1[2]);
  and and_a13_b20 (and_20[13], i0[13], i1[20]);
  and and_a13_b21 (and_21[13], i0[13], i1[21]);
  and and_a13_b22 (and_22[13], i0[13], i1[22]);
  and and_a13_b23 (and_23[13], i0[13], i1[23]);
  and and_a13_b24 (and_24[13], i0[13], i1[24]);
  and and_a13_b25 (and_25[13], i0[13], i1[25]);
  and and_a13_b26 (and_26[13], i0[13], i1[26]);
  and and_a13_b27 (and_27[13], i0[13], i1[27]);
  and and_a13_b28 (and_28[13], i0[13], i1[28]);
  and and_a13_b29 (and_29[13], i0[13], i1[29]);
  and and_a13_b3 (and_3[13], i0[13], i1[3]);
  and and_a13_b30 (and_30[13], i0[13], i1[30]);
  and and_a13_b31 (and_31[13], i0[13], i1[31]);
  and and_a13_b4 (and_4[13], i0[13], i1[4]);
  and and_a13_b5 (and_5[13], i0[13], i1[5]);
  and and_a13_b6 (and_6[13], i0[13], i1[6]);
  and and_a13_b7 (and_7[13], i0[13], i1[7]);
  and and_a13_b8 (and_8[13], i0[13], i1[8]);
  and and_a13_b9 (and_9[13], i0[13], i1[9]);
  and and_a14_b0 (and_0[14], i0[14], i1[0]);
  and and_a14_b1 (and_1[14], i0[14], i1[1]);
  and and_a14_b10 (and_10[14], i0[14], i1[10]);
  and and_a14_b11 (and_11[14], i0[14], i1[11]);
  and and_a14_b12 (and_12[14], i0[14], i1[12]);
  and and_a14_b13 (and_13[14], i0[14], i1[13]);
  and and_a14_b14 (and_14[14], i0[14], i1[14]);
  and and_a14_b15 (and_15[14], i0[14], i1[15]);
  and and_a14_b16 (and_16[14], i0[14], i1[16]);
  and and_a14_b17 (and_17[14], i0[14], i1[17]);
  and and_a14_b18 (and_18[14], i0[14], i1[18]);
  and and_a14_b19 (and_19[14], i0[14], i1[19]);
  and and_a14_b2 (and_2[14], i0[14], i1[2]);
  and and_a14_b20 (and_20[14], i0[14], i1[20]);
  and and_a14_b21 (and_21[14], i0[14], i1[21]);
  and and_a14_b22 (and_22[14], i0[14], i1[22]);
  and and_a14_b23 (and_23[14], i0[14], i1[23]);
  and and_a14_b24 (and_24[14], i0[14], i1[24]);
  and and_a14_b25 (and_25[14], i0[14], i1[25]);
  and and_a14_b26 (and_26[14], i0[14], i1[26]);
  and and_a14_b27 (and_27[14], i0[14], i1[27]);
  and and_a14_b28 (and_28[14], i0[14], i1[28]);
  and and_a14_b29 (and_29[14], i0[14], i1[29]);
  and and_a14_b3 (and_3[14], i0[14], i1[3]);
  and and_a14_b30 (and_30[14], i0[14], i1[30]);
  and and_a14_b31 (and_31[14], i0[14], i1[31]);
  and and_a14_b4 (and_4[14], i0[14], i1[4]);
  and and_a14_b5 (and_5[14], i0[14], i1[5]);
  and and_a14_b6 (and_6[14], i0[14], i1[6]);
  and and_a14_b7 (and_7[14], i0[14], i1[7]);
  and and_a14_b8 (and_8[14], i0[14], i1[8]);
  and and_a14_b9 (and_9[14], i0[14], i1[9]);
  and and_a15_b0 (and_0[15], i0[15], i1[0]);
  and and_a15_b1 (and_1[15], i0[15], i1[1]);
  and and_a15_b10 (and_10[15], i0[15], i1[10]);
  and and_a15_b11 (and_11[15], i0[15], i1[11]);
  and and_a15_b12 (and_12[15], i0[15], i1[12]);
  and and_a15_b13 (and_13[15], i0[15], i1[13]);
  and and_a15_b14 (and_14[15], i0[15], i1[14]);
  and and_a15_b15 (and_15[15], i0[15], i1[15]);
  and and_a15_b16 (and_16[15], i0[15], i1[16]);
  and and_a15_b17 (and_17[15], i0[15], i1[17]);
  and and_a15_b18 (and_18[15], i0[15], i1[18]);
  and and_a15_b19 (and_19[15], i0[15], i1[19]);
  and and_a15_b2 (and_2[15], i0[15], i1[2]);
  and and_a15_b20 (and_20[15], i0[15], i1[20]);
  and and_a15_b21 (and_21[15], i0[15], i1[21]);
  and and_a15_b22 (and_22[15], i0[15], i1[22]);
  and and_a15_b23 (and_23[15], i0[15], i1[23]);
  and and_a15_b24 (and_24[15], i0[15], i1[24]);
  and and_a15_b25 (and_25[15], i0[15], i1[25]);
  and and_a15_b26 (and_26[15], i0[15], i1[26]);
  and and_a15_b27 (and_27[15], i0[15], i1[27]);
  and and_a15_b28 (and_28[15], i0[15], i1[28]);
  and and_a15_b29 (and_29[15], i0[15], i1[29]);
  and and_a15_b3 (and_3[15], i0[15], i1[3]);
  and and_a15_b30 (and_30[15], i0[15], i1[30]);
  and and_a15_b31 (and_31[15], i0[15], i1[31]);
  and and_a15_b4 (and_4[15], i0[15], i1[4]);
  and and_a15_b5 (and_5[15], i0[15], i1[5]);
  and and_a15_b6 (and_6[15], i0[15], i1[6]);
  and and_a15_b7 (and_7[15], i0[15], i1[7]);
  and and_a15_b8 (and_8[15], i0[15], i1[8]);
  and and_a15_b9 (and_9[15], i0[15], i1[9]);
  and and_a16_b0 (and_0[16], i0[16], i1[0]);
  and and_a16_b1 (and_1[16], i0[16], i1[1]);
  and and_a16_b10 (and_10[16], i0[16], i1[10]);
  and and_a16_b11 (and_11[16], i0[16], i1[11]);
  and and_a16_b12 (and_12[16], i0[16], i1[12]);
  and and_a16_b13 (and_13[16], i0[16], i1[13]);
  and and_a16_b14 (and_14[16], i0[16], i1[14]);
  and and_a16_b15 (and_15[16], i0[16], i1[15]);
  and and_a16_b16 (and_16[16], i0[16], i1[16]);
  and and_a16_b17 (and_17[16], i0[16], i1[17]);
  and and_a16_b18 (and_18[16], i0[16], i1[18]);
  and and_a16_b19 (and_19[16], i0[16], i1[19]);
  and and_a16_b2 (and_2[16], i0[16], i1[2]);
  and and_a16_b20 (and_20[16], i0[16], i1[20]);
  and and_a16_b21 (and_21[16], i0[16], i1[21]);
  and and_a16_b22 (and_22[16], i0[16], i1[22]);
  and and_a16_b23 (and_23[16], i0[16], i1[23]);
  and and_a16_b24 (and_24[16], i0[16], i1[24]);
  and and_a16_b25 (and_25[16], i0[16], i1[25]);
  and and_a16_b26 (and_26[16], i0[16], i1[26]);
  and and_a16_b27 (and_27[16], i0[16], i1[27]);
  and and_a16_b28 (and_28[16], i0[16], i1[28]);
  and and_a16_b29 (and_29[16], i0[16], i1[29]);
  and and_a16_b3 (and_3[16], i0[16], i1[3]);
  and and_a16_b30 (and_30[16], i0[16], i1[30]);
  and and_a16_b31 (and_31[16], i0[16], i1[31]);
  and and_a16_b4 (and_4[16], i0[16], i1[4]);
  and and_a16_b5 (and_5[16], i0[16], i1[5]);
  and and_a16_b6 (and_6[16], i0[16], i1[6]);
  and and_a16_b7 (and_7[16], i0[16], i1[7]);
  and and_a16_b8 (and_8[16], i0[16], i1[8]);
  and and_a16_b9 (and_9[16], i0[16], i1[9]);
  and and_a17_b0 (and_0[17], i0[17], i1[0]);
  and and_a17_b1 (and_1[17], i0[17], i1[1]);
  and and_a17_b10 (and_10[17], i0[17], i1[10]);
  and and_a17_b11 (and_11[17], i0[17], i1[11]);
  and and_a17_b12 (and_12[17], i0[17], i1[12]);
  and and_a17_b13 (and_13[17], i0[17], i1[13]);
  and and_a17_b14 (and_14[17], i0[17], i1[14]);
  and and_a17_b15 (and_15[17], i0[17], i1[15]);
  and and_a17_b16 (and_16[17], i0[17], i1[16]);
  and and_a17_b17 (and_17[17], i0[17], i1[17]);
  and and_a17_b18 (and_18[17], i0[17], i1[18]);
  and and_a17_b19 (and_19[17], i0[17], i1[19]);
  and and_a17_b2 (and_2[17], i0[17], i1[2]);
  and and_a17_b20 (and_20[17], i0[17], i1[20]);
  and and_a17_b21 (and_21[17], i0[17], i1[21]);
  and and_a17_b22 (and_22[17], i0[17], i1[22]);
  and and_a17_b23 (and_23[17], i0[17], i1[23]);
  and and_a17_b24 (and_24[17], i0[17], i1[24]);
  and and_a17_b25 (and_25[17], i0[17], i1[25]);
  and and_a17_b26 (and_26[17], i0[17], i1[26]);
  and and_a17_b27 (and_27[17], i0[17], i1[27]);
  and and_a17_b28 (and_28[17], i0[17], i1[28]);
  and and_a17_b29 (and_29[17], i0[17], i1[29]);
  and and_a17_b3 (and_3[17], i0[17], i1[3]);
  and and_a17_b30 (and_30[17], i0[17], i1[30]);
  and and_a17_b31 (and_31[17], i0[17], i1[31]);
  and and_a17_b4 (and_4[17], i0[17], i1[4]);
  and and_a17_b5 (and_5[17], i0[17], i1[5]);
  and and_a17_b6 (and_6[17], i0[17], i1[6]);
  and and_a17_b7 (and_7[17], i0[17], i1[7]);
  and and_a17_b8 (and_8[17], i0[17], i1[8]);
  and and_a17_b9 (and_9[17], i0[17], i1[9]);
  and and_a18_b0 (and_0[18], i0[18], i1[0]);
  and and_a18_b1 (and_1[18], i0[18], i1[1]);
  and and_a18_b10 (and_10[18], i0[18], i1[10]);
  and and_a18_b11 (and_11[18], i0[18], i1[11]);
  and and_a18_b12 (and_12[18], i0[18], i1[12]);
  and and_a18_b13 (and_13[18], i0[18], i1[13]);
  and and_a18_b14 (and_14[18], i0[18], i1[14]);
  and and_a18_b15 (and_15[18], i0[18], i1[15]);
  and and_a18_b16 (and_16[18], i0[18], i1[16]);
  and and_a18_b17 (and_17[18], i0[18], i1[17]);
  and and_a18_b18 (and_18[18], i0[18], i1[18]);
  and and_a18_b19 (and_19[18], i0[18], i1[19]);
  and and_a18_b2 (and_2[18], i0[18], i1[2]);
  and and_a18_b20 (and_20[18], i0[18], i1[20]);
  and and_a18_b21 (and_21[18], i0[18], i1[21]);
  and and_a18_b22 (and_22[18], i0[18], i1[22]);
  and and_a18_b23 (and_23[18], i0[18], i1[23]);
  and and_a18_b24 (and_24[18], i0[18], i1[24]);
  and and_a18_b25 (and_25[18], i0[18], i1[25]);
  and and_a18_b26 (and_26[18], i0[18], i1[26]);
  and and_a18_b27 (and_27[18], i0[18], i1[27]);
  and and_a18_b28 (and_28[18], i0[18], i1[28]);
  and and_a18_b29 (and_29[18], i0[18], i1[29]);
  and and_a18_b3 (and_3[18], i0[18], i1[3]);
  and and_a18_b30 (and_30[18], i0[18], i1[30]);
  and and_a18_b31 (and_31[18], i0[18], i1[31]);
  and and_a18_b4 (and_4[18], i0[18], i1[4]);
  and and_a18_b5 (and_5[18], i0[18], i1[5]);
  and and_a18_b6 (and_6[18], i0[18], i1[6]);
  and and_a18_b7 (and_7[18], i0[18], i1[7]);
  and and_a18_b8 (and_8[18], i0[18], i1[8]);
  and and_a18_b9 (and_9[18], i0[18], i1[9]);
  and and_a19_b0 (and_0[19], i0[19], i1[0]);
  and and_a19_b1 (and_1[19], i0[19], i1[1]);
  and and_a19_b10 (and_10[19], i0[19], i1[10]);
  and and_a19_b11 (and_11[19], i0[19], i1[11]);
  and and_a19_b12 (and_12[19], i0[19], i1[12]);
  and and_a19_b13 (and_13[19], i0[19], i1[13]);
  and and_a19_b14 (and_14[19], i0[19], i1[14]);
  and and_a19_b15 (and_15[19], i0[19], i1[15]);
  and and_a19_b16 (and_16[19], i0[19], i1[16]);
  and and_a19_b17 (and_17[19], i0[19], i1[17]);
  and and_a19_b18 (and_18[19], i0[19], i1[18]);
  and and_a19_b19 (and_19[19], i0[19], i1[19]);
  and and_a19_b2 (and_2[19], i0[19], i1[2]);
  and and_a19_b20 (and_20[19], i0[19], i1[20]);
  and and_a19_b21 (and_21[19], i0[19], i1[21]);
  and and_a19_b22 (and_22[19], i0[19], i1[22]);
  and and_a19_b23 (and_23[19], i0[19], i1[23]);
  and and_a19_b24 (and_24[19], i0[19], i1[24]);
  and and_a19_b25 (and_25[19], i0[19], i1[25]);
  and and_a19_b26 (and_26[19], i0[19], i1[26]);
  and and_a19_b27 (and_27[19], i0[19], i1[27]);
  and and_a19_b28 (and_28[19], i0[19], i1[28]);
  and and_a19_b29 (and_29[19], i0[19], i1[29]);
  and and_a19_b3 (and_3[19], i0[19], i1[3]);
  and and_a19_b30 (and_30[19], i0[19], i1[30]);
  and and_a19_b31 (and_31[19], i0[19], i1[31]);
  and and_a19_b4 (and_4[19], i0[19], i1[4]);
  and and_a19_b5 (and_5[19], i0[19], i1[5]);
  and and_a19_b6 (and_6[19], i0[19], i1[6]);
  and and_a19_b7 (and_7[19], i0[19], i1[7]);
  and and_a19_b8 (and_8[19], i0[19], i1[8]);
  and and_a19_b9 (and_9[19], i0[19], i1[9]);
  and and_a1_b0 (and_0[1], i0[1], i1[0]);
  and and_a1_b1 (and_1[1], i0[1], i1[1]);
  and and_a1_b10 (and_10[1], i0[1], i1[10]);
  and and_a1_b11 (and_11[1], i0[1], i1[11]);
  and and_a1_b12 (and_12[1], i0[1], i1[12]);
  and and_a1_b13 (and_13[1], i0[1], i1[13]);
  and and_a1_b14 (and_14[1], i0[1], i1[14]);
  and and_a1_b15 (and_15[1], i0[1], i1[15]);
  and and_a1_b16 (and_16[1], i0[1], i1[16]);
  and and_a1_b17 (and_17[1], i0[1], i1[17]);
  and and_a1_b18 (and_18[1], i0[1], i1[18]);
  and and_a1_b19 (and_19[1], i0[1], i1[19]);
  and and_a1_b2 (and_2[1], i0[1], i1[2]);
  and and_a1_b20 (and_20[1], i0[1], i1[20]);
  and and_a1_b21 (and_21[1], i0[1], i1[21]);
  and and_a1_b22 (and_22[1], i0[1], i1[22]);
  and and_a1_b23 (and_23[1], i0[1], i1[23]);
  and and_a1_b24 (and_24[1], i0[1], i1[24]);
  and and_a1_b25 (and_25[1], i0[1], i1[25]);
  and and_a1_b26 (and_26[1], i0[1], i1[26]);
  and and_a1_b27 (and_27[1], i0[1], i1[27]);
  and and_a1_b28 (and_28[1], i0[1], i1[28]);
  and and_a1_b29 (and_29[1], i0[1], i1[29]);
  and and_a1_b3 (and_3[1], i0[1], i1[3]);
  and and_a1_b30 (and_30[1], i0[1], i1[30]);
  and and_a1_b31 (and_31[1], i0[1], i1[31]);
  and and_a1_b4 (and_4[1], i0[1], i1[4]);
  and and_a1_b5 (and_5[1], i0[1], i1[5]);
  and and_a1_b6 (and_6[1], i0[1], i1[6]);
  and and_a1_b7 (and_7[1], i0[1], i1[7]);
  and and_a1_b8 (and_8[1], i0[1], i1[8]);
  and and_a1_b9 (and_9[1], i0[1], i1[9]);
  and and_a20_b0 (and_0[20], i0[20], i1[0]);
  and and_a20_b1 (and_1[20], i0[20], i1[1]);
  and and_a20_b10 (and_10[20], i0[20], i1[10]);
  and and_a20_b11 (and_11[20], i0[20], i1[11]);
  and and_a20_b12 (and_12[20], i0[20], i1[12]);
  and and_a20_b13 (and_13[20], i0[20], i1[13]);
  and and_a20_b14 (and_14[20], i0[20], i1[14]);
  and and_a20_b15 (and_15[20], i0[20], i1[15]);
  and and_a20_b16 (and_16[20], i0[20], i1[16]);
  and and_a20_b17 (and_17[20], i0[20], i1[17]);
  and and_a20_b18 (and_18[20], i0[20], i1[18]);
  and and_a20_b19 (and_19[20], i0[20], i1[19]);
  and and_a20_b2 (and_2[20], i0[20], i1[2]);
  and and_a20_b20 (and_20[20], i0[20], i1[20]);
  and and_a20_b21 (and_21[20], i0[20], i1[21]);
  and and_a20_b22 (and_22[20], i0[20], i1[22]);
  and and_a20_b23 (and_23[20], i0[20], i1[23]);
  and and_a20_b24 (and_24[20], i0[20], i1[24]);
  and and_a20_b25 (and_25[20], i0[20], i1[25]);
  and and_a20_b26 (and_26[20], i0[20], i1[26]);
  and and_a20_b27 (and_27[20], i0[20], i1[27]);
  and and_a20_b28 (and_28[20], i0[20], i1[28]);
  and and_a20_b29 (and_29[20], i0[20], i1[29]);
  and and_a20_b3 (and_3[20], i0[20], i1[3]);
  and and_a20_b30 (and_30[20], i0[20], i1[30]);
  and and_a20_b31 (and_31[20], i0[20], i1[31]);
  and and_a20_b4 (and_4[20], i0[20], i1[4]);
  and and_a20_b5 (and_5[20], i0[20], i1[5]);
  and and_a20_b6 (and_6[20], i0[20], i1[6]);
  and and_a20_b7 (and_7[20], i0[20], i1[7]);
  and and_a20_b8 (and_8[20], i0[20], i1[8]);
  and and_a20_b9 (and_9[20], i0[20], i1[9]);
  and and_a21_b0 (and_0[21], i0[21], i1[0]);
  and and_a21_b1 (and_1[21], i0[21], i1[1]);
  and and_a21_b10 (and_10[21], i0[21], i1[10]);
  and and_a21_b11 (and_11[21], i0[21], i1[11]);
  and and_a21_b12 (and_12[21], i0[21], i1[12]);
  and and_a21_b13 (and_13[21], i0[21], i1[13]);
  and and_a21_b14 (and_14[21], i0[21], i1[14]);
  and and_a21_b15 (and_15[21], i0[21], i1[15]);
  and and_a21_b16 (and_16[21], i0[21], i1[16]);
  and and_a21_b17 (and_17[21], i0[21], i1[17]);
  and and_a21_b18 (and_18[21], i0[21], i1[18]);
  and and_a21_b19 (and_19[21], i0[21], i1[19]);
  and and_a21_b2 (and_2[21], i0[21], i1[2]);
  and and_a21_b20 (and_20[21], i0[21], i1[20]);
  and and_a21_b21 (and_21[21], i0[21], i1[21]);
  and and_a21_b22 (and_22[21], i0[21], i1[22]);
  and and_a21_b23 (and_23[21], i0[21], i1[23]);
  and and_a21_b24 (and_24[21], i0[21], i1[24]);
  and and_a21_b25 (and_25[21], i0[21], i1[25]);
  and and_a21_b26 (and_26[21], i0[21], i1[26]);
  and and_a21_b27 (and_27[21], i0[21], i1[27]);
  and and_a21_b28 (and_28[21], i0[21], i1[28]);
  and and_a21_b29 (and_29[21], i0[21], i1[29]);
  and and_a21_b3 (and_3[21], i0[21], i1[3]);
  and and_a21_b30 (and_30[21], i0[21], i1[30]);
  and and_a21_b31 (and_31[21], i0[21], i1[31]);
  and and_a21_b4 (and_4[21], i0[21], i1[4]);
  and and_a21_b5 (and_5[21], i0[21], i1[5]);
  and and_a21_b6 (and_6[21], i0[21], i1[6]);
  and and_a21_b7 (and_7[21], i0[21], i1[7]);
  and and_a21_b8 (and_8[21], i0[21], i1[8]);
  and and_a21_b9 (and_9[21], i0[21], i1[9]);
  and and_a22_b0 (and_0[22], i0[22], i1[0]);
  and and_a22_b1 (and_1[22], i0[22], i1[1]);
  and and_a22_b10 (and_10[22], i0[22], i1[10]);
  and and_a22_b11 (and_11[22], i0[22], i1[11]);
  and and_a22_b12 (and_12[22], i0[22], i1[12]);
  and and_a22_b13 (and_13[22], i0[22], i1[13]);
  and and_a22_b14 (and_14[22], i0[22], i1[14]);
  and and_a22_b15 (and_15[22], i0[22], i1[15]);
  and and_a22_b16 (and_16[22], i0[22], i1[16]);
  and and_a22_b17 (and_17[22], i0[22], i1[17]);
  and and_a22_b18 (and_18[22], i0[22], i1[18]);
  and and_a22_b19 (and_19[22], i0[22], i1[19]);
  and and_a22_b2 (and_2[22], i0[22], i1[2]);
  and and_a22_b20 (and_20[22], i0[22], i1[20]);
  and and_a22_b21 (and_21[22], i0[22], i1[21]);
  and and_a22_b22 (and_22[22], i0[22], i1[22]);
  and and_a22_b23 (and_23[22], i0[22], i1[23]);
  and and_a22_b24 (and_24[22], i0[22], i1[24]);
  and and_a22_b25 (and_25[22], i0[22], i1[25]);
  and and_a22_b26 (and_26[22], i0[22], i1[26]);
  and and_a22_b27 (and_27[22], i0[22], i1[27]);
  and and_a22_b28 (and_28[22], i0[22], i1[28]);
  and and_a22_b29 (and_29[22], i0[22], i1[29]);
  and and_a22_b3 (and_3[22], i0[22], i1[3]);
  and and_a22_b30 (and_30[22], i0[22], i1[30]);
  and and_a22_b31 (and_31[22], i0[22], i1[31]);
  and and_a22_b4 (and_4[22], i0[22], i1[4]);
  and and_a22_b5 (and_5[22], i0[22], i1[5]);
  and and_a22_b6 (and_6[22], i0[22], i1[6]);
  and and_a22_b7 (and_7[22], i0[22], i1[7]);
  and and_a22_b8 (and_8[22], i0[22], i1[8]);
  and and_a22_b9 (and_9[22], i0[22], i1[9]);
  and and_a23_b0 (and_0[23], i0[23], i1[0]);
  and and_a23_b1 (and_1[23], i0[23], i1[1]);
  and and_a23_b10 (and_10[23], i0[23], i1[10]);
  and and_a23_b11 (and_11[23], i0[23], i1[11]);
  and and_a23_b12 (and_12[23], i0[23], i1[12]);
  and and_a23_b13 (and_13[23], i0[23], i1[13]);
  and and_a23_b14 (and_14[23], i0[23], i1[14]);
  and and_a23_b15 (and_15[23], i0[23], i1[15]);
  and and_a23_b16 (and_16[23], i0[23], i1[16]);
  and and_a23_b17 (and_17[23], i0[23], i1[17]);
  and and_a23_b18 (and_18[23], i0[23], i1[18]);
  and and_a23_b19 (and_19[23], i0[23], i1[19]);
  and and_a23_b2 (and_2[23], i0[23], i1[2]);
  and and_a23_b20 (and_20[23], i0[23], i1[20]);
  and and_a23_b21 (and_21[23], i0[23], i1[21]);
  and and_a23_b22 (and_22[23], i0[23], i1[22]);
  and and_a23_b23 (and_23[23], i0[23], i1[23]);
  and and_a23_b24 (and_24[23], i0[23], i1[24]);
  and and_a23_b25 (and_25[23], i0[23], i1[25]);
  and and_a23_b26 (and_26[23], i0[23], i1[26]);
  and and_a23_b27 (and_27[23], i0[23], i1[27]);
  and and_a23_b28 (and_28[23], i0[23], i1[28]);
  and and_a23_b29 (and_29[23], i0[23], i1[29]);
  and and_a23_b3 (and_3[23], i0[23], i1[3]);
  and and_a23_b30 (and_30[23], i0[23], i1[30]);
  and and_a23_b31 (and_31[23], i0[23], i1[31]);
  and and_a23_b4 (and_4[23], i0[23], i1[4]);
  and and_a23_b5 (and_5[23], i0[23], i1[5]);
  and and_a23_b6 (and_6[23], i0[23], i1[6]);
  and and_a23_b7 (and_7[23], i0[23], i1[7]);
  and and_a23_b8 (and_8[23], i0[23], i1[8]);
  and and_a23_b9 (and_9[23], i0[23], i1[9]);
  and and_a24_b0 (and_0[24], i0[24], i1[0]);
  and and_a24_b1 (and_1[24], i0[24], i1[1]);
  and and_a24_b10 (and_10[24], i0[24], i1[10]);
  and and_a24_b11 (and_11[24], i0[24], i1[11]);
  and and_a24_b12 (and_12[24], i0[24], i1[12]);
  and and_a24_b13 (and_13[24], i0[24], i1[13]);
  and and_a24_b14 (and_14[24], i0[24], i1[14]);
  and and_a24_b15 (and_15[24], i0[24], i1[15]);
  and and_a24_b16 (and_16[24], i0[24], i1[16]);
  and and_a24_b17 (and_17[24], i0[24], i1[17]);
  and and_a24_b18 (and_18[24], i0[24], i1[18]);
  and and_a24_b19 (and_19[24], i0[24], i1[19]);
  and and_a24_b2 (and_2[24], i0[24], i1[2]);
  and and_a24_b20 (and_20[24], i0[24], i1[20]);
  and and_a24_b21 (and_21[24], i0[24], i1[21]);
  and and_a24_b22 (and_22[24], i0[24], i1[22]);
  and and_a24_b23 (and_23[24], i0[24], i1[23]);
  and and_a24_b24 (and_24[24], i0[24], i1[24]);
  and and_a24_b25 (and_25[24], i0[24], i1[25]);
  and and_a24_b26 (and_26[24], i0[24], i1[26]);
  and and_a24_b27 (and_27[24], i0[24], i1[27]);
  and and_a24_b28 (and_28[24], i0[24], i1[28]);
  and and_a24_b29 (and_29[24], i0[24], i1[29]);
  and and_a24_b3 (and_3[24], i0[24], i1[3]);
  and and_a24_b30 (and_30[24], i0[24], i1[30]);
  and and_a24_b31 (and_31[24], i0[24], i1[31]);
  and and_a24_b4 (and_4[24], i0[24], i1[4]);
  and and_a24_b5 (and_5[24], i0[24], i1[5]);
  and and_a24_b6 (and_6[24], i0[24], i1[6]);
  and and_a24_b7 (and_7[24], i0[24], i1[7]);
  and and_a24_b8 (and_8[24], i0[24], i1[8]);
  and and_a24_b9 (and_9[24], i0[24], i1[9]);
  and and_a25_b0 (and_0[25], i0[25], i1[0]);
  and and_a25_b1 (and_1[25], i0[25], i1[1]);
  and and_a25_b10 (and_10[25], i0[25], i1[10]);
  and and_a25_b11 (and_11[25], i0[25], i1[11]);
  and and_a25_b12 (and_12[25], i0[25], i1[12]);
  and and_a25_b13 (and_13[25], i0[25], i1[13]);
  and and_a25_b14 (and_14[25], i0[25], i1[14]);
  and and_a25_b15 (and_15[25], i0[25], i1[15]);
  and and_a25_b16 (and_16[25], i0[25], i1[16]);
  and and_a25_b17 (and_17[25], i0[25], i1[17]);
  and and_a25_b18 (and_18[25], i0[25], i1[18]);
  and and_a25_b19 (and_19[25], i0[25], i1[19]);
  and and_a25_b2 (and_2[25], i0[25], i1[2]);
  and and_a25_b20 (and_20[25], i0[25], i1[20]);
  and and_a25_b21 (and_21[25], i0[25], i1[21]);
  and and_a25_b22 (and_22[25], i0[25], i1[22]);
  and and_a25_b23 (and_23[25], i0[25], i1[23]);
  and and_a25_b24 (and_24[25], i0[25], i1[24]);
  and and_a25_b25 (and_25[25], i0[25], i1[25]);
  and and_a25_b26 (and_26[25], i0[25], i1[26]);
  and and_a25_b27 (and_27[25], i0[25], i1[27]);
  and and_a25_b28 (and_28[25], i0[25], i1[28]);
  and and_a25_b29 (and_29[25], i0[25], i1[29]);
  and and_a25_b3 (and_3[25], i0[25], i1[3]);
  and and_a25_b30 (and_30[25], i0[25], i1[30]);
  and and_a25_b31 (and_31[25], i0[25], i1[31]);
  and and_a25_b4 (and_4[25], i0[25], i1[4]);
  and and_a25_b5 (and_5[25], i0[25], i1[5]);
  and and_a25_b6 (and_6[25], i0[25], i1[6]);
  and and_a25_b7 (and_7[25], i0[25], i1[7]);
  and and_a25_b8 (and_8[25], i0[25], i1[8]);
  and and_a25_b9 (and_9[25], i0[25], i1[9]);
  and and_a26_b0 (and_0[26], i0[26], i1[0]);
  and and_a26_b1 (and_1[26], i0[26], i1[1]);
  and and_a26_b10 (and_10[26], i0[26], i1[10]);
  and and_a26_b11 (and_11[26], i0[26], i1[11]);
  and and_a26_b12 (and_12[26], i0[26], i1[12]);
  and and_a26_b13 (and_13[26], i0[26], i1[13]);
  and and_a26_b14 (and_14[26], i0[26], i1[14]);
  and and_a26_b15 (and_15[26], i0[26], i1[15]);
  and and_a26_b16 (and_16[26], i0[26], i1[16]);
  and and_a26_b17 (and_17[26], i0[26], i1[17]);
  and and_a26_b18 (and_18[26], i0[26], i1[18]);
  and and_a26_b19 (and_19[26], i0[26], i1[19]);
  and and_a26_b2 (and_2[26], i0[26], i1[2]);
  and and_a26_b20 (and_20[26], i0[26], i1[20]);
  and and_a26_b21 (and_21[26], i0[26], i1[21]);
  and and_a26_b22 (and_22[26], i0[26], i1[22]);
  and and_a26_b23 (and_23[26], i0[26], i1[23]);
  and and_a26_b24 (and_24[26], i0[26], i1[24]);
  and and_a26_b25 (and_25[26], i0[26], i1[25]);
  and and_a26_b26 (and_26[26], i0[26], i1[26]);
  and and_a26_b27 (and_27[26], i0[26], i1[27]);
  and and_a26_b28 (and_28[26], i0[26], i1[28]);
  and and_a26_b29 (and_29[26], i0[26], i1[29]);
  and and_a26_b3 (and_3[26], i0[26], i1[3]);
  and and_a26_b30 (and_30[26], i0[26], i1[30]);
  and and_a26_b31 (and_31[26], i0[26], i1[31]);
  and and_a26_b4 (and_4[26], i0[26], i1[4]);
  and and_a26_b5 (and_5[26], i0[26], i1[5]);
  and and_a26_b6 (and_6[26], i0[26], i1[6]);
  and and_a26_b7 (and_7[26], i0[26], i1[7]);
  and and_a26_b8 (and_8[26], i0[26], i1[8]);
  and and_a26_b9 (and_9[26], i0[26], i1[9]);
  and and_a27_b0 (and_0[27], i0[27], i1[0]);
  and and_a27_b1 (and_1[27], i0[27], i1[1]);
  and and_a27_b10 (and_10[27], i0[27], i1[10]);
  and and_a27_b11 (and_11[27], i0[27], i1[11]);
  and and_a27_b12 (and_12[27], i0[27], i1[12]);
  and and_a27_b13 (and_13[27], i0[27], i1[13]);
  and and_a27_b14 (and_14[27], i0[27], i1[14]);
  and and_a27_b15 (and_15[27], i0[27], i1[15]);
  and and_a27_b16 (and_16[27], i0[27], i1[16]);
  and and_a27_b17 (and_17[27], i0[27], i1[17]);
  and and_a27_b18 (and_18[27], i0[27], i1[18]);
  and and_a27_b19 (and_19[27], i0[27], i1[19]);
  and and_a27_b2 (and_2[27], i0[27], i1[2]);
  and and_a27_b20 (and_20[27], i0[27], i1[20]);
  and and_a27_b21 (and_21[27], i0[27], i1[21]);
  and and_a27_b22 (and_22[27], i0[27], i1[22]);
  and and_a27_b23 (and_23[27], i0[27], i1[23]);
  and and_a27_b24 (and_24[27], i0[27], i1[24]);
  and and_a27_b25 (and_25[27], i0[27], i1[25]);
  and and_a27_b26 (and_26[27], i0[27], i1[26]);
  and and_a27_b27 (and_27[27], i0[27], i1[27]);
  and and_a27_b28 (and_28[27], i0[27], i1[28]);
  and and_a27_b29 (and_29[27], i0[27], i1[29]);
  and and_a27_b3 (and_3[27], i0[27], i1[3]);
  and and_a27_b30 (and_30[27], i0[27], i1[30]);
  and and_a27_b31 (and_31[27], i0[27], i1[31]);
  and and_a27_b4 (and_4[27], i0[27], i1[4]);
  and and_a27_b5 (and_5[27], i0[27], i1[5]);
  and and_a27_b6 (and_6[27], i0[27], i1[6]);
  and and_a27_b7 (and_7[27], i0[27], i1[7]);
  and and_a27_b8 (and_8[27], i0[27], i1[8]);
  and and_a27_b9 (and_9[27], i0[27], i1[9]);
  and and_a28_b0 (and_0[28], i0[28], i1[0]);
  and and_a28_b1 (and_1[28], i0[28], i1[1]);
  and and_a28_b10 (and_10[28], i0[28], i1[10]);
  and and_a28_b11 (and_11[28], i0[28], i1[11]);
  and and_a28_b12 (and_12[28], i0[28], i1[12]);
  and and_a28_b13 (and_13[28], i0[28], i1[13]);
  and and_a28_b14 (and_14[28], i0[28], i1[14]);
  and and_a28_b15 (and_15[28], i0[28], i1[15]);
  and and_a28_b16 (and_16[28], i0[28], i1[16]);
  and and_a28_b17 (and_17[28], i0[28], i1[17]);
  and and_a28_b18 (and_18[28], i0[28], i1[18]);
  and and_a28_b19 (and_19[28], i0[28], i1[19]);
  and and_a28_b2 (and_2[28], i0[28], i1[2]);
  and and_a28_b20 (and_20[28], i0[28], i1[20]);
  and and_a28_b21 (and_21[28], i0[28], i1[21]);
  and and_a28_b22 (and_22[28], i0[28], i1[22]);
  and and_a28_b23 (and_23[28], i0[28], i1[23]);
  and and_a28_b24 (and_24[28], i0[28], i1[24]);
  and and_a28_b25 (and_25[28], i0[28], i1[25]);
  and and_a28_b26 (and_26[28], i0[28], i1[26]);
  and and_a28_b27 (and_27[28], i0[28], i1[27]);
  and and_a28_b28 (and_28[28], i0[28], i1[28]);
  and and_a28_b29 (and_29[28], i0[28], i1[29]);
  and and_a28_b3 (and_3[28], i0[28], i1[3]);
  and and_a28_b30 (and_30[28], i0[28], i1[30]);
  and and_a28_b31 (and_31[28], i0[28], i1[31]);
  and and_a28_b4 (and_4[28], i0[28], i1[4]);
  and and_a28_b5 (and_5[28], i0[28], i1[5]);
  and and_a28_b6 (and_6[28], i0[28], i1[6]);
  and and_a28_b7 (and_7[28], i0[28], i1[7]);
  and and_a28_b8 (and_8[28], i0[28], i1[8]);
  and and_a28_b9 (and_9[28], i0[28], i1[9]);
  and and_a29_b0 (and_0[29], i0[29], i1[0]);
  and and_a29_b1 (and_1[29], i0[29], i1[1]);
  and and_a29_b10 (and_10[29], i0[29], i1[10]);
  and and_a29_b11 (and_11[29], i0[29], i1[11]);
  and and_a29_b12 (and_12[29], i0[29], i1[12]);
  and and_a29_b13 (and_13[29], i0[29], i1[13]);
  and and_a29_b14 (and_14[29], i0[29], i1[14]);
  and and_a29_b15 (and_15[29], i0[29], i1[15]);
  and and_a29_b16 (and_16[29], i0[29], i1[16]);
  and and_a29_b17 (and_17[29], i0[29], i1[17]);
  and and_a29_b18 (and_18[29], i0[29], i1[18]);
  and and_a29_b19 (and_19[29], i0[29], i1[19]);
  and and_a29_b2 (and_2[29], i0[29], i1[2]);
  and and_a29_b20 (and_20[29], i0[29], i1[20]);
  and and_a29_b21 (and_21[29], i0[29], i1[21]);
  and and_a29_b22 (and_22[29], i0[29], i1[22]);
  and and_a29_b23 (and_23[29], i0[29], i1[23]);
  and and_a29_b24 (and_24[29], i0[29], i1[24]);
  and and_a29_b25 (and_25[29], i0[29], i1[25]);
  and and_a29_b26 (and_26[29], i0[29], i1[26]);
  and and_a29_b27 (and_27[29], i0[29], i1[27]);
  and and_a29_b28 (and_28[29], i0[29], i1[28]);
  and and_a29_b29 (and_29[29], i0[29], i1[29]);
  and and_a29_b3 (and_3[29], i0[29], i1[3]);
  and and_a29_b30 (and_30[29], i0[29], i1[30]);
  and and_a29_b31 (and_31[29], i0[29], i1[31]);
  and and_a29_b4 (and_4[29], i0[29], i1[4]);
  and and_a29_b5 (and_5[29], i0[29], i1[5]);
  and and_a29_b6 (and_6[29], i0[29], i1[6]);
  and and_a29_b7 (and_7[29], i0[29], i1[7]);
  and and_a29_b8 (and_8[29], i0[29], i1[8]);
  and and_a29_b9 (and_9[29], i0[29], i1[9]);
  and and_a2_b0 (and_0[2], i0[2], i1[0]);
  and and_a2_b1 (and_1[2], i0[2], i1[1]);
  and and_a2_b10 (and_10[2], i0[2], i1[10]);
  and and_a2_b11 (and_11[2], i0[2], i1[11]);
  and and_a2_b12 (and_12[2], i0[2], i1[12]);
  and and_a2_b13 (and_13[2], i0[2], i1[13]);
  and and_a2_b14 (and_14[2], i0[2], i1[14]);
  and and_a2_b15 (and_15[2], i0[2], i1[15]);
  and and_a2_b16 (and_16[2], i0[2], i1[16]);
  and and_a2_b17 (and_17[2], i0[2], i1[17]);
  and and_a2_b18 (and_18[2], i0[2], i1[18]);
  and and_a2_b19 (and_19[2], i0[2], i1[19]);
  and and_a2_b2 (and_2[2], i0[2], i1[2]);
  and and_a2_b20 (and_20[2], i0[2], i1[20]);
  and and_a2_b21 (and_21[2], i0[2], i1[21]);
  and and_a2_b22 (and_22[2], i0[2], i1[22]);
  and and_a2_b23 (and_23[2], i0[2], i1[23]);
  and and_a2_b24 (and_24[2], i0[2], i1[24]);
  and and_a2_b25 (and_25[2], i0[2], i1[25]);
  and and_a2_b26 (and_26[2], i0[2], i1[26]);
  and and_a2_b27 (and_27[2], i0[2], i1[27]);
  and and_a2_b28 (and_28[2], i0[2], i1[28]);
  and and_a2_b29 (and_29[2], i0[2], i1[29]);
  and and_a2_b3 (and_3[2], i0[2], i1[3]);
  and and_a2_b30 (and_30[2], i0[2], i1[30]);
  and and_a2_b31 (and_31[2], i0[2], i1[31]);
  and and_a2_b4 (and_4[2], i0[2], i1[4]);
  and and_a2_b5 (and_5[2], i0[2], i1[5]);
  and and_a2_b6 (and_6[2], i0[2], i1[6]);
  and and_a2_b7 (and_7[2], i0[2], i1[7]);
  and and_a2_b8 (and_8[2], i0[2], i1[8]);
  and and_a2_b9 (and_9[2], i0[2], i1[9]);
  and and_a30_b0 (and_0[30], i0[30], i1[0]);
  and and_a30_b1 (and_1[30], i0[30], i1[1]);
  and and_a30_b10 (and_10[30], i0[30], i1[10]);
  and and_a30_b11 (and_11[30], i0[30], i1[11]);
  and and_a30_b12 (and_12[30], i0[30], i1[12]);
  and and_a30_b13 (and_13[30], i0[30], i1[13]);
  and and_a30_b14 (and_14[30], i0[30], i1[14]);
  and and_a30_b15 (and_15[30], i0[30], i1[15]);
  and and_a30_b16 (and_16[30], i0[30], i1[16]);
  and and_a30_b17 (and_17[30], i0[30], i1[17]);
  and and_a30_b18 (and_18[30], i0[30], i1[18]);
  and and_a30_b19 (and_19[30], i0[30], i1[19]);
  and and_a30_b2 (and_2[30], i0[30], i1[2]);
  and and_a30_b20 (and_20[30], i0[30], i1[20]);
  and and_a30_b21 (and_21[30], i0[30], i1[21]);
  and and_a30_b22 (and_22[30], i0[30], i1[22]);
  and and_a30_b23 (and_23[30], i0[30], i1[23]);
  and and_a30_b24 (and_24[30], i0[30], i1[24]);
  and and_a30_b25 (and_25[30], i0[30], i1[25]);
  and and_a30_b26 (and_26[30], i0[30], i1[26]);
  and and_a30_b27 (and_27[30], i0[30], i1[27]);
  and and_a30_b28 (and_28[30], i0[30], i1[28]);
  and and_a30_b29 (and_29[30], i0[30], i1[29]);
  and and_a30_b3 (and_3[30], i0[30], i1[3]);
  and and_a30_b30 (and_30[30], i0[30], i1[30]);
  and and_a30_b31 (and_31[30], i0[30], i1[31]);
  and and_a30_b4 (and_4[30], i0[30], i1[4]);
  and and_a30_b5 (and_5[30], i0[30], i1[5]);
  and and_a30_b6 (and_6[30], i0[30], i1[6]);
  and and_a30_b7 (and_7[30], i0[30], i1[7]);
  and and_a30_b8 (and_8[30], i0[30], i1[8]);
  and and_a30_b9 (and_9[30], i0[30], i1[9]);
  and and_a31_b0 (and_0[31], i0[31], i1[0]);
  and and_a31_b1 (and_1[31], i0[31], i1[1]);
  and and_a31_b10 (and_10[31], i0[31], i1[10]);
  and and_a31_b11 (and_11[31], i0[31], i1[11]);
  and and_a31_b12 (and_12[31], i0[31], i1[12]);
  and and_a31_b13 (and_13[31], i0[31], i1[13]);
  and and_a31_b14 (and_14[31], i0[31], i1[14]);
  and and_a31_b15 (and_15[31], i0[31], i1[15]);
  and and_a31_b16 (and_16[31], i0[31], i1[16]);
  and and_a31_b17 (and_17[31], i0[31], i1[17]);
  and and_a31_b18 (and_18[31], i0[31], i1[18]);
  and and_a31_b19 (and_19[31], i0[31], i1[19]);
  and and_a31_b2 (and_2[31], i0[31], i1[2]);
  and and_a31_b20 (and_20[31], i0[31], i1[20]);
  and and_a31_b21 (and_21[31], i0[31], i1[21]);
  and and_a31_b22 (and_22[31], i0[31], i1[22]);
  and and_a31_b23 (and_23[31], i0[31], i1[23]);
  and and_a31_b24 (and_24[31], i0[31], i1[24]);
  and and_a31_b25 (and_25[31], i0[31], i1[25]);
  and and_a31_b26 (and_26[31], i0[31], i1[26]);
  and and_a31_b27 (and_27[31], i0[31], i1[27]);
  and and_a31_b28 (and_28[31], i0[31], i1[28]);
  and and_a31_b29 (and_29[31], i0[31], i1[29]);
  and and_a31_b3 (and_3[31], i0[31], i1[3]);
  and and_a31_b30 (and_30[31], i0[31], i1[30]);
  and and_a31_b31 (and_31[31], i0[31], i1[31]);
  and and_a31_b4 (and_4[31], i0[31], i1[4]);
  and and_a31_b5 (and_5[31], i0[31], i1[5]);
  and and_a31_b6 (and_6[31], i0[31], i1[6]);
  and and_a31_b7 (and_7[31], i0[31], i1[7]);
  and and_a31_b8 (and_8[31], i0[31], i1[8]);
  and and_a31_b9 (and_9[31], i0[31], i1[9]);
  and and_a3_b0 (and_0[3], i0[3], i1[0]);
  and and_a3_b1 (and_1[3], i0[3], i1[1]);
  and and_a3_b10 (and_10[3], i0[3], i1[10]);
  and and_a3_b11 (and_11[3], i0[3], i1[11]);
  and and_a3_b12 (and_12[3], i0[3], i1[12]);
  and and_a3_b13 (and_13[3], i0[3], i1[13]);
  and and_a3_b14 (and_14[3], i0[3], i1[14]);
  and and_a3_b15 (and_15[3], i0[3], i1[15]);
  and and_a3_b16 (and_16[3], i0[3], i1[16]);
  and and_a3_b17 (and_17[3], i0[3], i1[17]);
  and and_a3_b18 (and_18[3], i0[3], i1[18]);
  and and_a3_b19 (and_19[3], i0[3], i1[19]);
  and and_a3_b2 (and_2[3], i0[3], i1[2]);
  and and_a3_b20 (and_20[3], i0[3], i1[20]);
  and and_a3_b21 (and_21[3], i0[3], i1[21]);
  and and_a3_b22 (and_22[3], i0[3], i1[22]);
  and and_a3_b23 (and_23[3], i0[3], i1[23]);
  and and_a3_b24 (and_24[3], i0[3], i1[24]);
  and and_a3_b25 (and_25[3], i0[3], i1[25]);
  and and_a3_b26 (and_26[3], i0[3], i1[26]);
  and and_a3_b27 (and_27[3], i0[3], i1[27]);
  and and_a3_b28 (and_28[3], i0[3], i1[28]);
  and and_a3_b29 (and_29[3], i0[3], i1[29]);
  and and_a3_b3 (and_3[3], i0[3], i1[3]);
  and and_a3_b30 (and_30[3], i0[3], i1[30]);
  and and_a3_b31 (and_31[3], i0[3], i1[31]);
  and and_a3_b4 (and_4[3], i0[3], i1[4]);
  and and_a3_b5 (and_5[3], i0[3], i1[5]);
  and and_a3_b6 (and_6[3], i0[3], i1[6]);
  and and_a3_b7 (and_7[3], i0[3], i1[7]);
  and and_a3_b8 (and_8[3], i0[3], i1[8]);
  and and_a3_b9 (and_9[3], i0[3], i1[9]);
  and and_a4_b0 (and_0[4], i0[4], i1[0]);
  and and_a4_b1 (and_1[4], i0[4], i1[1]);
  and and_a4_b10 (and_10[4], i0[4], i1[10]);
  and and_a4_b11 (and_11[4], i0[4], i1[11]);
  and and_a4_b12 (and_12[4], i0[4], i1[12]);
  and and_a4_b13 (and_13[4], i0[4], i1[13]);
  and and_a4_b14 (and_14[4], i0[4], i1[14]);
  and and_a4_b15 (and_15[4], i0[4], i1[15]);
  and and_a4_b16 (and_16[4], i0[4], i1[16]);
  and and_a4_b17 (and_17[4], i0[4], i1[17]);
  and and_a4_b18 (and_18[4], i0[4], i1[18]);
  and and_a4_b19 (and_19[4], i0[4], i1[19]);
  and and_a4_b2 (and_2[4], i0[4], i1[2]);
  and and_a4_b20 (and_20[4], i0[4], i1[20]);
  and and_a4_b21 (and_21[4], i0[4], i1[21]);
  and and_a4_b22 (and_22[4], i0[4], i1[22]);
  and and_a4_b23 (and_23[4], i0[4], i1[23]);
  and and_a4_b24 (and_24[4], i0[4], i1[24]);
  and and_a4_b25 (and_25[4], i0[4], i1[25]);
  and and_a4_b26 (and_26[4], i0[4], i1[26]);
  and and_a4_b27 (and_27[4], i0[4], i1[27]);
  and and_a4_b28 (and_28[4], i0[4], i1[28]);
  and and_a4_b29 (and_29[4], i0[4], i1[29]);
  and and_a4_b3 (and_3[4], i0[4], i1[3]);
  and and_a4_b30 (and_30[4], i0[4], i1[30]);
  and and_a4_b31 (and_31[4], i0[4], i1[31]);
  and and_a4_b4 (and_4[4], i0[4], i1[4]);
  and and_a4_b5 (and_5[4], i0[4], i1[5]);
  and and_a4_b6 (and_6[4], i0[4], i1[6]);
  and and_a4_b7 (and_7[4], i0[4], i1[7]);
  and and_a4_b8 (and_8[4], i0[4], i1[8]);
  and and_a4_b9 (and_9[4], i0[4], i1[9]);
  and and_a5_b0 (and_0[5], i0[5], i1[0]);
  and and_a5_b1 (and_1[5], i0[5], i1[1]);
  and and_a5_b10 (and_10[5], i0[5], i1[10]);
  and and_a5_b11 (and_11[5], i0[5], i1[11]);
  and and_a5_b12 (and_12[5], i0[5], i1[12]);
  and and_a5_b13 (and_13[5], i0[5], i1[13]);
  and and_a5_b14 (and_14[5], i0[5], i1[14]);
  and and_a5_b15 (and_15[5], i0[5], i1[15]);
  and and_a5_b16 (and_16[5], i0[5], i1[16]);
  and and_a5_b17 (and_17[5], i0[5], i1[17]);
  and and_a5_b18 (and_18[5], i0[5], i1[18]);
  and and_a5_b19 (and_19[5], i0[5], i1[19]);
  and and_a5_b2 (and_2[5], i0[5], i1[2]);
  and and_a5_b20 (and_20[5], i0[5], i1[20]);
  and and_a5_b21 (and_21[5], i0[5], i1[21]);
  and and_a5_b22 (and_22[5], i0[5], i1[22]);
  and and_a5_b23 (and_23[5], i0[5], i1[23]);
  and and_a5_b24 (and_24[5], i0[5], i1[24]);
  and and_a5_b25 (and_25[5], i0[5], i1[25]);
  and and_a5_b26 (and_26[5], i0[5], i1[26]);
  and and_a5_b27 (and_27[5], i0[5], i1[27]);
  and and_a5_b28 (and_28[5], i0[5], i1[28]);
  and and_a5_b29 (and_29[5], i0[5], i1[29]);
  and and_a5_b3 (and_3[5], i0[5], i1[3]);
  and and_a5_b30 (and_30[5], i0[5], i1[30]);
  and and_a5_b31 (and_31[5], i0[5], i1[31]);
  and and_a5_b4 (and_4[5], i0[5], i1[4]);
  and and_a5_b5 (and_5[5], i0[5], i1[5]);
  and and_a5_b6 (and_6[5], i0[5], i1[6]);
  and and_a5_b7 (and_7[5], i0[5], i1[7]);
  and and_a5_b8 (and_8[5], i0[5], i1[8]);
  and and_a5_b9 (and_9[5], i0[5], i1[9]);
  and and_a6_b0 (and_0[6], i0[6], i1[0]);
  and and_a6_b1 (and_1[6], i0[6], i1[1]);
  and and_a6_b10 (and_10[6], i0[6], i1[10]);
  and and_a6_b11 (and_11[6], i0[6], i1[11]);
  and and_a6_b12 (and_12[6], i0[6], i1[12]);
  and and_a6_b13 (and_13[6], i0[6], i1[13]);
  and and_a6_b14 (and_14[6], i0[6], i1[14]);
  and and_a6_b15 (and_15[6], i0[6], i1[15]);
  and and_a6_b16 (and_16[6], i0[6], i1[16]);
  and and_a6_b17 (and_17[6], i0[6], i1[17]);
  and and_a6_b18 (and_18[6], i0[6], i1[18]);
  and and_a6_b19 (and_19[6], i0[6], i1[19]);
  and and_a6_b2 (and_2[6], i0[6], i1[2]);
  and and_a6_b20 (and_20[6], i0[6], i1[20]);
  and and_a6_b21 (and_21[6], i0[6], i1[21]);
  and and_a6_b22 (and_22[6], i0[6], i1[22]);
  and and_a6_b23 (and_23[6], i0[6], i1[23]);
  and and_a6_b24 (and_24[6], i0[6], i1[24]);
  and and_a6_b25 (and_25[6], i0[6], i1[25]);
  and and_a6_b26 (and_26[6], i0[6], i1[26]);
  and and_a6_b27 (and_27[6], i0[6], i1[27]);
  and and_a6_b28 (and_28[6], i0[6], i1[28]);
  and and_a6_b29 (and_29[6], i0[6], i1[29]);
  and and_a6_b3 (and_3[6], i0[6], i1[3]);
  and and_a6_b30 (and_30[6], i0[6], i1[30]);
  and and_a6_b31 (and_31[6], i0[6], i1[31]);
  and and_a6_b4 (and_4[6], i0[6], i1[4]);
  and and_a6_b5 (and_5[6], i0[6], i1[5]);
  and and_a6_b6 (and_6[6], i0[6], i1[6]);
  and and_a6_b7 (and_7[6], i0[6], i1[7]);
  and and_a6_b8 (and_8[6], i0[6], i1[8]);
  and and_a6_b9 (and_9[6], i0[6], i1[9]);
  and and_a7_b0 (and_0[7], i0[7], i1[0]);
  and and_a7_b1 (and_1[7], i0[7], i1[1]);
  and and_a7_b10 (and_10[7], i0[7], i1[10]);
  and and_a7_b11 (and_11[7], i0[7], i1[11]);
  and and_a7_b12 (and_12[7], i0[7], i1[12]);
  and and_a7_b13 (and_13[7], i0[7], i1[13]);
  and and_a7_b14 (and_14[7], i0[7], i1[14]);
  and and_a7_b15 (and_15[7], i0[7], i1[15]);
  and and_a7_b16 (and_16[7], i0[7], i1[16]);
  and and_a7_b17 (and_17[7], i0[7], i1[17]);
  and and_a7_b18 (and_18[7], i0[7], i1[18]);
  and and_a7_b19 (and_19[7], i0[7], i1[19]);
  and and_a7_b2 (and_2[7], i0[7], i1[2]);
  and and_a7_b20 (and_20[7], i0[7], i1[20]);
  and and_a7_b21 (and_21[7], i0[7], i1[21]);
  and and_a7_b22 (and_22[7], i0[7], i1[22]);
  and and_a7_b23 (and_23[7], i0[7], i1[23]);
  and and_a7_b24 (and_24[7], i0[7], i1[24]);
  and and_a7_b25 (and_25[7], i0[7], i1[25]);
  and and_a7_b26 (and_26[7], i0[7], i1[26]);
  and and_a7_b27 (and_27[7], i0[7], i1[27]);
  and and_a7_b28 (and_28[7], i0[7], i1[28]);
  and and_a7_b29 (and_29[7], i0[7], i1[29]);
  and and_a7_b3 (and_3[7], i0[7], i1[3]);
  and and_a7_b30 (and_30[7], i0[7], i1[30]);
  and and_a7_b31 (and_31[7], i0[7], i1[31]);
  and and_a7_b4 (and_4[7], i0[7], i1[4]);
  and and_a7_b5 (and_5[7], i0[7], i1[5]);
  and and_a7_b6 (and_6[7], i0[7], i1[6]);
  and and_a7_b7 (and_7[7], i0[7], i1[7]);
  and and_a7_b8 (and_8[7], i0[7], i1[8]);
  and and_a7_b9 (and_9[7], i0[7], i1[9]);
  and and_a8_b0 (and_0[8], i0[8], i1[0]);
  and and_a8_b1 (and_1[8], i0[8], i1[1]);
  and and_a8_b10 (and_10[8], i0[8], i1[10]);
  and and_a8_b11 (and_11[8], i0[8], i1[11]);
  and and_a8_b12 (and_12[8], i0[8], i1[12]);
  and and_a8_b13 (and_13[8], i0[8], i1[13]);
  and and_a8_b14 (and_14[8], i0[8], i1[14]);
  and and_a8_b15 (and_15[8], i0[8], i1[15]);
  and and_a8_b16 (and_16[8], i0[8], i1[16]);
  and and_a8_b17 (and_17[8], i0[8], i1[17]);
  and and_a8_b18 (and_18[8], i0[8], i1[18]);
  and and_a8_b19 (and_19[8], i0[8], i1[19]);
  and and_a8_b2 (and_2[8], i0[8], i1[2]);
  and and_a8_b20 (and_20[8], i0[8], i1[20]);
  and and_a8_b21 (and_21[8], i0[8], i1[21]);
  and and_a8_b22 (and_22[8], i0[8], i1[22]);
  and and_a8_b23 (and_23[8], i0[8], i1[23]);
  and and_a8_b24 (and_24[8], i0[8], i1[24]);
  and and_a8_b25 (and_25[8], i0[8], i1[25]);
  and and_a8_b26 (and_26[8], i0[8], i1[26]);
  and and_a8_b27 (and_27[8], i0[8], i1[27]);
  and and_a8_b28 (and_28[8], i0[8], i1[28]);
  and and_a8_b29 (and_29[8], i0[8], i1[29]);
  and and_a8_b3 (and_3[8], i0[8], i1[3]);
  and and_a8_b30 (and_30[8], i0[8], i1[30]);
  and and_a8_b31 (and_31[8], i0[8], i1[31]);
  and and_a8_b4 (and_4[8], i0[8], i1[4]);
  and and_a8_b5 (and_5[8], i0[8], i1[5]);
  and and_a8_b6 (and_6[8], i0[8], i1[6]);
  and and_a8_b7 (and_7[8], i0[8], i1[7]);
  and and_a8_b8 (and_8[8], i0[8], i1[8]);
  and and_a8_b9 (and_9[8], i0[8], i1[9]);
  and and_a9_b0 (and_0[9], i0[9], i1[0]);
  and and_a9_b1 (and_1[9], i0[9], i1[1]);
  and and_a9_b10 (and_10[9], i0[9], i1[10]);
  and and_a9_b11 (and_11[9], i0[9], i1[11]);
  and and_a9_b12 (and_12[9], i0[9], i1[12]);
  and and_a9_b13 (and_13[9], i0[9], i1[13]);
  and and_a9_b14 (and_14[9], i0[9], i1[14]);
  and and_a9_b15 (and_15[9], i0[9], i1[15]);
  and and_a9_b16 (and_16[9], i0[9], i1[16]);
  and and_a9_b17 (and_17[9], i0[9], i1[17]);
  and and_a9_b18 (and_18[9], i0[9], i1[18]);
  and and_a9_b19 (and_19[9], i0[9], i1[19]);
  and and_a9_b2 (and_2[9], i0[9], i1[2]);
  and and_a9_b20 (and_20[9], i0[9], i1[20]);
  and and_a9_b21 (and_21[9], i0[9], i1[21]);
  and and_a9_b22 (and_22[9], i0[9], i1[22]);
  and and_a9_b23 (and_23[9], i0[9], i1[23]);
  and and_a9_b24 (and_24[9], i0[9], i1[24]);
  and and_a9_b25 (and_25[9], i0[9], i1[25]);
  and and_a9_b26 (and_26[9], i0[9], i1[26]);
  and and_a9_b27 (and_27[9], i0[9], i1[27]);
  and and_a9_b28 (and_28[9], i0[9], i1[28]);
  and and_a9_b29 (and_29[9], i0[9], i1[29]);
  and and_a9_b3 (and_3[9], i0[9], i1[3]);
  and and_a9_b30 (and_30[9], i0[9], i1[30]);
  and and_a9_b31 (and_31[9], i0[9], i1[31]);
  and and_a9_b4 (and_4[9], i0[9], i1[4]);
  and and_a9_b5 (and_5[9], i0[9], i1[5]);
  and and_a9_b6 (and_6[9], i0[9], i1[6]);
  and and_a9_b7 (and_7[9], i0[9], i1[7]);
  and and_a9_b8 (and_8[9], i0[9], i1[8]);
  and and_a9_b9 (and_9[9], i0[9], i1[9]);
  add_pu63_pu62_pu61_pu60_pu59_pu58_pu57_pu56_pu55_pu54_pu53_pu52_pu51_pu50_pu49_pu48_pu47_pu46_pu45_pu44_pu43_pu42_pu41_pu40_pu39_pu38_pu37_pu36_pu35_pu34_pu33_pu32_o64 sum (
    .i0({and_31[31],and_30[31],and_29[31],and_28[31],and_27[31],and_26[31],and_25[31],and_24[31],and_23[31],and_22[31],and_21[31],and_20[31],and_19[31],and_18[31],and_17[31],and_16[31],and_15[31],and_14[31],and_13[31],and_12[31],and_11[31],and_10[31],and_9[31],and_8[31],and_7[31],and_6[31],and_5[31],and_4[31],and_3[31],and_2[31],and_1[31],and_0}),
    .i1({and_31[30],and_30[30],and_29[30],and_28[30],and_27[30],and_26[30],and_25[30],and_24[30],and_23[30],and_22[30],and_21[30],and_20[30],and_19[30],and_18[30],and_17[30],and_16[30],and_15[30],and_14[30],and_13[30],and_12[30],and_11[30],and_10[30],and_9[30],and_8[30],and_7[30],and_6[30],and_5[30],and_4[30],and_3[30],and_2[30],and_1[30:0],1'b0}),
    .i10({and_31[21],and_30[21],and_29[21],and_28[21],and_27[21],and_26[21],and_25[21],and_24[21],and_23[21],and_22[21],and_21[21],and_20[21],and_19[21],and_18[21],and_17[21],and_16[21],and_15[21],and_14[21],and_13[21],and_12[21],and_11[21],and_10[21:0],10'b0000000000}),
    .i11({and_31[20],and_30[20],and_29[20],and_28[20],and_27[20],and_26[20],and_25[20],and_24[20],and_23[20],and_22[20],and_21[20],and_20[20],and_19[20],and_18[20],and_17[20],and_16[20],and_15[20],and_14[20],and_13[20],and_12[20],and_11[20:0],11'b00000000000}),
    .i12({and_31[19],and_30[19],and_29[19],and_28[19],and_27[19],and_26[19],and_25[19],and_24[19],and_23[19],and_22[19],and_21[19],and_20[19],and_19[19],and_18[19],and_17[19],and_16[19],and_15[19],and_14[19],and_13[19],and_12[19:0],12'b000000000000}),
    .i13({and_31[18],and_30[18],and_29[18],and_28[18],and_27[18],and_26[18],and_25[18],and_24[18],and_23[18],and_22[18],and_21[18],and_20[18],and_19[18],and_18[18],and_17[18],and_16[18],and_15[18],and_14[18],and_13[18:0],13'b0000000000000}),
    .i14({and_31[17],and_30[17],and_29[17],and_28[17],and_27[17],and_26[17],and_25[17],and_24[17],and_23[17],and_22[17],and_21[17],and_20[17],and_19[17],and_18[17],and_17[17],and_16[17],and_15[17],and_14[17:0],14'b00000000000000}),
    .i15({and_31[16],and_30[16],and_29[16],and_28[16],and_27[16],and_26[16],and_25[16],and_24[16],and_23[16],and_22[16],and_21[16],and_20[16],and_19[16],and_18[16],and_17[16],and_16[16],and_15[16:0],15'b000000000000000}),
    .i16({and_31[15],and_30[15],and_29[15],and_28[15],and_27[15],and_26[15],and_25[15],and_24[15],and_23[15],and_22[15],and_21[15],and_20[15],and_19[15],and_18[15],and_17[15],and_16[15:0],16'b0000000000000000}),
    .i17({and_31[14],and_30[14],and_29[14],and_28[14],and_27[14],and_26[14],and_25[14],and_24[14],and_23[14],and_22[14],and_21[14],and_20[14],and_19[14],and_18[14],and_17[14:0],17'b00000000000000000}),
    .i18({and_31[13],and_30[13],and_29[13],and_28[13],and_27[13],and_26[13],and_25[13],and_24[13],and_23[13],and_22[13],and_21[13],and_20[13],and_19[13],and_18[13:0],18'b000000000000000000}),
    .i19({and_31[12],and_30[12],and_29[12],and_28[12],and_27[12],and_26[12],and_25[12],and_24[12],and_23[12],and_22[12],and_21[12],and_20[12],and_19[12:0],19'b0000000000000000000}),
    .i2({and_31[29],and_30[29],and_29[29],and_28[29],and_27[29],and_26[29],and_25[29],and_24[29],and_23[29],and_22[29],and_21[29],and_20[29],and_19[29],and_18[29],and_17[29],and_16[29],and_15[29],and_14[29],and_13[29],and_12[29],and_11[29],and_10[29],and_9[29],and_8[29],and_7[29],and_6[29],and_5[29],and_4[29],and_3[29],and_2[29:0],2'b00}),
    .i20({and_31[11],and_30[11],and_29[11],and_28[11],and_27[11],and_26[11],and_25[11],and_24[11],and_23[11],and_22[11],and_21[11],and_20[11:0],20'b00000000000000000000}),
    .i21({and_31[10],and_30[10],and_29[10],and_28[10],and_27[10],and_26[10],and_25[10],and_24[10],and_23[10],and_22[10],and_21[10:0],21'b000000000000000000000}),
    .i22({and_31[9],and_30[9],and_29[9],and_28[9],and_27[9],and_26[9],and_25[9],and_24[9],and_23[9],and_22[9:0],22'b0000000000000000000000}),
    .i23({and_31[8],and_30[8],and_29[8],and_28[8],and_27[8],and_26[8],and_25[8],and_24[8],and_23[8:0],23'b00000000000000000000000}),
    .i24({and_31[7],and_30[7],and_29[7],and_28[7],and_27[7],and_26[7],and_25[7],and_24[7:0],24'b000000000000000000000000}),
    .i25({and_31[6],and_30[6],and_29[6],and_28[6],and_27[6],and_26[6],and_25[6:0],25'b0000000000000000000000000}),
    .i26({and_31[5],and_30[5],and_29[5],and_28[5],and_27[5],and_26[5:0],26'b00000000000000000000000000}),
    .i27({and_31[4],and_30[4],and_29[4],and_28[4],and_27[4:0],27'b000000000000000000000000000}),
    .i28({and_31[3],and_30[3],and_29[3],and_28[3:0],28'b0000000000000000000000000000}),
    .i29({and_31[2],and_30[2],and_29[2:0],29'b00000000000000000000000000000}),
    .i3({and_31[28],and_30[28],and_29[28],and_28[28],and_27[28],and_26[28],and_25[28],and_24[28],and_23[28],and_22[28],and_21[28],and_20[28],and_19[28],and_18[28],and_17[28],and_16[28],and_15[28],and_14[28],and_13[28],and_12[28],and_11[28],and_10[28],and_9[28],and_8[28],and_7[28],and_6[28],and_5[28],and_4[28],and_3[28:0],3'b000}),
    .i30({and_31[1],and_30[1:0],30'b000000000000000000000000000000}),
    .i31({and_31[0],31'b0000000000000000000000000000000}),
    .i4({and_31[27],and_30[27],and_29[27],and_28[27],and_27[27],and_26[27],and_25[27],and_24[27],and_23[27],and_22[27],and_21[27],and_20[27],and_19[27],and_18[27],and_17[27],and_16[27],and_15[27],and_14[27],and_13[27],and_12[27],and_11[27],and_10[27],and_9[27],and_8[27],and_7[27],and_6[27],and_5[27],and_4[27:0],4'b0000}),
    .i5({and_31[26],and_30[26],and_29[26],and_28[26],and_27[26],and_26[26],and_25[26],and_24[26],and_23[26],and_22[26],and_21[26],and_20[26],and_19[26],and_18[26],and_17[26],and_16[26],and_15[26],and_14[26],and_13[26],and_12[26],and_11[26],and_10[26],and_9[26],and_8[26],and_7[26],and_6[26],and_5[26:0],5'b00000}),
    .i6({and_31[25],and_30[25],and_29[25],and_28[25],and_27[25],and_26[25],and_25[25],and_24[25],and_23[25],and_22[25],and_21[25],and_20[25],and_19[25],and_18[25],and_17[25],and_16[25],and_15[25],and_14[25],and_13[25],and_12[25],and_11[25],and_10[25],and_9[25],and_8[25],and_7[25],and_6[25:0],6'b000000}),
    .i7({and_31[24],and_30[24],and_29[24],and_28[24],and_27[24],and_26[24],and_25[24],and_24[24],and_23[24],and_22[24],and_21[24],and_20[24],and_19[24],and_18[24],and_17[24],and_16[24],and_15[24],and_14[24],and_13[24],and_12[24],and_11[24],and_10[24],and_9[24],and_8[24],and_7[24:0],7'b0000000}),
    .i8({and_31[23],and_30[23],and_29[23],and_28[23],and_27[23],and_26[23],and_25[23],and_24[23],and_23[23],and_22[23],and_21[23],and_20[23],and_19[23],and_18[23],and_17[23],and_16[23],and_15[23],and_14[23],and_13[23],and_12[23],and_11[23],and_10[23],and_9[23],and_8[23:0],8'b00000000}),
    .i9({and_31[22],and_30[22],and_29[22],and_28[22],and_27[22],and_26[22],and_25[22],and_24[22],and_23[22],and_22[22],and_21[22],and_20[22],and_19[22],and_18[22],and_17[22],and_16[22],and_15[22],and_14[22],and_13[22],and_12[22],and_11[22],and_10[22],and_9[22:0],9'b000000000}),
    .o(o));

endmodule 

module mult_s32_s33_o64
  (
  i0,
  i1,
  o
  );

  input signed [31:0] i0;
  input signed [32:0] i1;
  output [63:0] o;

  wire [31:0] and_0;
  wire [31:0] and_1;
  wire [31:0] and_10;
  wire [31:0] and_11;
  wire [31:0] and_12;
  wire [31:0] and_13;
  wire [31:0] and_14;
  wire [31:0] and_15;
  wire [31:0] and_16;
  wire [31:0] and_17;
  wire [31:0] and_18;
  wire [31:0] and_19;
  wire [31:0] and_2;
  wire [31:0] and_20;
  wire [31:0] and_21;
  wire [31:0] and_22;
  wire [31:0] and_23;
  wire [31:0] and_24;
  wire [31:0] and_25;
  wire [31:0] and_26;
  wire [31:0] and_27;
  wire [31:0] and_28;
  wire [31:0] and_29;
  wire [31:0] and_3;
  wire [31:0] and_30;
  wire [31:0] and_31;
  wire [31:0] and_32;
  wire [31:0] and_4;
  wire [31:0] and_5;
  wire [31:0] and_6;
  wire [31:0] and_7;
  wire [31:0] and_8;
  wire [31:0] and_9;
  wire [31:0] nand_0;
  wire [31:0] nand_1;
  wire [31:0] nand_10;
  wire [31:0] nand_11;
  wire [31:0] nand_12;
  wire [31:0] nand_13;
  wire [31:0] nand_14;
  wire [31:0] nand_15;
  wire [31:0] nand_16;
  wire [31:0] nand_17;
  wire [31:0] nand_18;
  wire [31:0] nand_19;
  wire [31:0] nand_2;
  wire [31:0] nand_20;
  wire [31:0] nand_21;
  wire [31:0] nand_22;
  wire [31:0] nand_23;
  wire [31:0] nand_24;
  wire [31:0] nand_25;
  wire [31:0] nand_26;
  wire [31:0] nand_27;
  wire [31:0] nand_28;
  wire [31:0] nand_29;
  wire [31:0] nand_3;
  wire [31:0] nand_30;
  wire [31:0] nand_31;
  wire [31:0] nand_32;
  wire [31:0] nand_4;
  wire [31:0] nand_5;
  wire [31:0] nand_6;
  wire [31:0] nand_7;
  wire [31:0] nand_8;
  wire [31:0] nand_9;

  and and_a0_b0 (and_0[0], i0[0], i1[0]);
  and and_a0_b1 (and_1[0], i0[0], i1[1]);
  and and_a0_b10 (and_10[0], i0[0], i1[10]);
  and and_a0_b11 (and_11[0], i0[0], i1[11]);
  and and_a0_b12 (and_12[0], i0[0], i1[12]);
  and and_a0_b13 (and_13[0], i0[0], i1[13]);
  and and_a0_b14 (and_14[0], i0[0], i1[14]);
  and and_a0_b15 (and_15[0], i0[0], i1[15]);
  and and_a0_b16 (and_16[0], i0[0], i1[16]);
  and and_a0_b17 (and_17[0], i0[0], i1[17]);
  and and_a0_b18 (and_18[0], i0[0], i1[18]);
  and and_a0_b19 (and_19[0], i0[0], i1[19]);
  and and_a0_b2 (and_2[0], i0[0], i1[2]);
  and and_a0_b20 (and_20[0], i0[0], i1[20]);
  and and_a0_b21 (and_21[0], i0[0], i1[21]);
  and and_a0_b22 (and_22[0], i0[0], i1[22]);
  and and_a0_b23 (and_23[0], i0[0], i1[23]);
  and and_a0_b24 (and_24[0], i0[0], i1[24]);
  and and_a0_b25 (and_25[0], i0[0], i1[25]);
  and and_a0_b26 (and_26[0], i0[0], i1[26]);
  and and_a0_b27 (and_27[0], i0[0], i1[27]);
  and and_a0_b28 (and_28[0], i0[0], i1[28]);
  and and_a0_b29 (and_29[0], i0[0], i1[29]);
  and and_a0_b3 (and_3[0], i0[0], i1[3]);
  and and_a0_b30 (and_30[0], i0[0], i1[30]);
  and and_a0_b31 (and_31[0], i0[0], i1[31]);
  and and_a0_b32 (nand_32[0], i0[0], i1[32]);
  and and_a0_b4 (and_4[0], i0[0], i1[4]);
  and and_a0_b5 (and_5[0], i0[0], i1[5]);
  and and_a0_b6 (and_6[0], i0[0], i1[6]);
  and and_a0_b7 (and_7[0], i0[0], i1[7]);
  and and_a0_b8 (and_8[0], i0[0], i1[8]);
  and and_a0_b9 (and_9[0], i0[0], i1[9]);
  and and_a10_b0 (and_0[10], i0[10], i1[0]);
  and and_a10_b1 (and_1[10], i0[10], i1[1]);
  and and_a10_b10 (and_10[10], i0[10], i1[10]);
  and and_a10_b11 (and_11[10], i0[10], i1[11]);
  and and_a10_b12 (and_12[10], i0[10], i1[12]);
  and and_a10_b13 (and_13[10], i0[10], i1[13]);
  and and_a10_b14 (and_14[10], i0[10], i1[14]);
  and and_a10_b15 (and_15[10], i0[10], i1[15]);
  and and_a10_b16 (and_16[10], i0[10], i1[16]);
  and and_a10_b17 (and_17[10], i0[10], i1[17]);
  and and_a10_b18 (and_18[10], i0[10], i1[18]);
  and and_a10_b19 (and_19[10], i0[10], i1[19]);
  and and_a10_b2 (and_2[10], i0[10], i1[2]);
  and and_a10_b20 (and_20[10], i0[10], i1[20]);
  and and_a10_b21 (and_21[10], i0[10], i1[21]);
  and and_a10_b22 (and_22[10], i0[10], i1[22]);
  and and_a10_b23 (and_23[10], i0[10], i1[23]);
  and and_a10_b24 (and_24[10], i0[10], i1[24]);
  and and_a10_b25 (and_25[10], i0[10], i1[25]);
  and and_a10_b26 (and_26[10], i0[10], i1[26]);
  and and_a10_b27 (and_27[10], i0[10], i1[27]);
  and and_a10_b28 (and_28[10], i0[10], i1[28]);
  and and_a10_b29 (and_29[10], i0[10], i1[29]);
  and and_a10_b3 (and_3[10], i0[10], i1[3]);
  and and_a10_b30 (and_30[10], i0[10], i1[30]);
  and and_a10_b31 (and_31[10], i0[10], i1[31]);
  and and_a10_b32 (nand_32[10], i0[10], i1[32]);
  and and_a10_b4 (and_4[10], i0[10], i1[4]);
  and and_a10_b5 (and_5[10], i0[10], i1[5]);
  and and_a10_b6 (and_6[10], i0[10], i1[6]);
  and and_a10_b7 (and_7[10], i0[10], i1[7]);
  and and_a10_b8 (and_8[10], i0[10], i1[8]);
  and and_a10_b9 (and_9[10], i0[10], i1[9]);
  and and_a11_b0 (and_0[11], i0[11], i1[0]);
  and and_a11_b1 (and_1[11], i0[11], i1[1]);
  and and_a11_b10 (and_10[11], i0[11], i1[10]);
  and and_a11_b11 (and_11[11], i0[11], i1[11]);
  and and_a11_b12 (and_12[11], i0[11], i1[12]);
  and and_a11_b13 (and_13[11], i0[11], i1[13]);
  and and_a11_b14 (and_14[11], i0[11], i1[14]);
  and and_a11_b15 (and_15[11], i0[11], i1[15]);
  and and_a11_b16 (and_16[11], i0[11], i1[16]);
  and and_a11_b17 (and_17[11], i0[11], i1[17]);
  and and_a11_b18 (and_18[11], i0[11], i1[18]);
  and and_a11_b19 (and_19[11], i0[11], i1[19]);
  and and_a11_b2 (and_2[11], i0[11], i1[2]);
  and and_a11_b20 (and_20[11], i0[11], i1[20]);
  and and_a11_b21 (and_21[11], i0[11], i1[21]);
  and and_a11_b22 (and_22[11], i0[11], i1[22]);
  and and_a11_b23 (and_23[11], i0[11], i1[23]);
  and and_a11_b24 (and_24[11], i0[11], i1[24]);
  and and_a11_b25 (and_25[11], i0[11], i1[25]);
  and and_a11_b26 (and_26[11], i0[11], i1[26]);
  and and_a11_b27 (and_27[11], i0[11], i1[27]);
  and and_a11_b28 (and_28[11], i0[11], i1[28]);
  and and_a11_b29 (and_29[11], i0[11], i1[29]);
  and and_a11_b3 (and_3[11], i0[11], i1[3]);
  and and_a11_b30 (and_30[11], i0[11], i1[30]);
  and and_a11_b31 (and_31[11], i0[11], i1[31]);
  and and_a11_b32 (nand_32[11], i0[11], i1[32]);
  and and_a11_b4 (and_4[11], i0[11], i1[4]);
  and and_a11_b5 (and_5[11], i0[11], i1[5]);
  and and_a11_b6 (and_6[11], i0[11], i1[6]);
  and and_a11_b7 (and_7[11], i0[11], i1[7]);
  and and_a11_b8 (and_8[11], i0[11], i1[8]);
  and and_a11_b9 (and_9[11], i0[11], i1[9]);
  and and_a12_b0 (and_0[12], i0[12], i1[0]);
  and and_a12_b1 (and_1[12], i0[12], i1[1]);
  and and_a12_b10 (and_10[12], i0[12], i1[10]);
  and and_a12_b11 (and_11[12], i0[12], i1[11]);
  and and_a12_b12 (and_12[12], i0[12], i1[12]);
  and and_a12_b13 (and_13[12], i0[12], i1[13]);
  and and_a12_b14 (and_14[12], i0[12], i1[14]);
  and and_a12_b15 (and_15[12], i0[12], i1[15]);
  and and_a12_b16 (and_16[12], i0[12], i1[16]);
  and and_a12_b17 (and_17[12], i0[12], i1[17]);
  and and_a12_b18 (and_18[12], i0[12], i1[18]);
  and and_a12_b19 (and_19[12], i0[12], i1[19]);
  and and_a12_b2 (and_2[12], i0[12], i1[2]);
  and and_a12_b20 (and_20[12], i0[12], i1[20]);
  and and_a12_b21 (and_21[12], i0[12], i1[21]);
  and and_a12_b22 (and_22[12], i0[12], i1[22]);
  and and_a12_b23 (and_23[12], i0[12], i1[23]);
  and and_a12_b24 (and_24[12], i0[12], i1[24]);
  and and_a12_b25 (and_25[12], i0[12], i1[25]);
  and and_a12_b26 (and_26[12], i0[12], i1[26]);
  and and_a12_b27 (and_27[12], i0[12], i1[27]);
  and and_a12_b28 (and_28[12], i0[12], i1[28]);
  and and_a12_b29 (and_29[12], i0[12], i1[29]);
  and and_a12_b3 (and_3[12], i0[12], i1[3]);
  and and_a12_b30 (and_30[12], i0[12], i1[30]);
  and and_a12_b31 (and_31[12], i0[12], i1[31]);
  and and_a12_b32 (nand_32[12], i0[12], i1[32]);
  and and_a12_b4 (and_4[12], i0[12], i1[4]);
  and and_a12_b5 (and_5[12], i0[12], i1[5]);
  and and_a12_b6 (and_6[12], i0[12], i1[6]);
  and and_a12_b7 (and_7[12], i0[12], i1[7]);
  and and_a12_b8 (and_8[12], i0[12], i1[8]);
  and and_a12_b9 (and_9[12], i0[12], i1[9]);
  and and_a13_b0 (and_0[13], i0[13], i1[0]);
  and and_a13_b1 (and_1[13], i0[13], i1[1]);
  and and_a13_b10 (and_10[13], i0[13], i1[10]);
  and and_a13_b11 (and_11[13], i0[13], i1[11]);
  and and_a13_b12 (and_12[13], i0[13], i1[12]);
  and and_a13_b13 (and_13[13], i0[13], i1[13]);
  and and_a13_b14 (and_14[13], i0[13], i1[14]);
  and and_a13_b15 (and_15[13], i0[13], i1[15]);
  and and_a13_b16 (and_16[13], i0[13], i1[16]);
  and and_a13_b17 (and_17[13], i0[13], i1[17]);
  and and_a13_b18 (and_18[13], i0[13], i1[18]);
  and and_a13_b19 (and_19[13], i0[13], i1[19]);
  and and_a13_b2 (and_2[13], i0[13], i1[2]);
  and and_a13_b20 (and_20[13], i0[13], i1[20]);
  and and_a13_b21 (and_21[13], i0[13], i1[21]);
  and and_a13_b22 (and_22[13], i0[13], i1[22]);
  and and_a13_b23 (and_23[13], i0[13], i1[23]);
  and and_a13_b24 (and_24[13], i0[13], i1[24]);
  and and_a13_b25 (and_25[13], i0[13], i1[25]);
  and and_a13_b26 (and_26[13], i0[13], i1[26]);
  and and_a13_b27 (and_27[13], i0[13], i1[27]);
  and and_a13_b28 (and_28[13], i0[13], i1[28]);
  and and_a13_b29 (and_29[13], i0[13], i1[29]);
  and and_a13_b3 (and_3[13], i0[13], i1[3]);
  and and_a13_b30 (and_30[13], i0[13], i1[30]);
  and and_a13_b31 (and_31[13], i0[13], i1[31]);
  and and_a13_b32 (nand_32[13], i0[13], i1[32]);
  and and_a13_b4 (and_4[13], i0[13], i1[4]);
  and and_a13_b5 (and_5[13], i0[13], i1[5]);
  and and_a13_b6 (and_6[13], i0[13], i1[6]);
  and and_a13_b7 (and_7[13], i0[13], i1[7]);
  and and_a13_b8 (and_8[13], i0[13], i1[8]);
  and and_a13_b9 (and_9[13], i0[13], i1[9]);
  and and_a14_b0 (and_0[14], i0[14], i1[0]);
  and and_a14_b1 (and_1[14], i0[14], i1[1]);
  and and_a14_b10 (and_10[14], i0[14], i1[10]);
  and and_a14_b11 (and_11[14], i0[14], i1[11]);
  and and_a14_b12 (and_12[14], i0[14], i1[12]);
  and and_a14_b13 (and_13[14], i0[14], i1[13]);
  and and_a14_b14 (and_14[14], i0[14], i1[14]);
  and and_a14_b15 (and_15[14], i0[14], i1[15]);
  and and_a14_b16 (and_16[14], i0[14], i1[16]);
  and and_a14_b17 (and_17[14], i0[14], i1[17]);
  and and_a14_b18 (and_18[14], i0[14], i1[18]);
  and and_a14_b19 (and_19[14], i0[14], i1[19]);
  and and_a14_b2 (and_2[14], i0[14], i1[2]);
  and and_a14_b20 (and_20[14], i0[14], i1[20]);
  and and_a14_b21 (and_21[14], i0[14], i1[21]);
  and and_a14_b22 (and_22[14], i0[14], i1[22]);
  and and_a14_b23 (and_23[14], i0[14], i1[23]);
  and and_a14_b24 (and_24[14], i0[14], i1[24]);
  and and_a14_b25 (and_25[14], i0[14], i1[25]);
  and and_a14_b26 (and_26[14], i0[14], i1[26]);
  and and_a14_b27 (and_27[14], i0[14], i1[27]);
  and and_a14_b28 (and_28[14], i0[14], i1[28]);
  and and_a14_b29 (and_29[14], i0[14], i1[29]);
  and and_a14_b3 (and_3[14], i0[14], i1[3]);
  and and_a14_b30 (and_30[14], i0[14], i1[30]);
  and and_a14_b31 (and_31[14], i0[14], i1[31]);
  and and_a14_b32 (nand_32[14], i0[14], i1[32]);
  and and_a14_b4 (and_4[14], i0[14], i1[4]);
  and and_a14_b5 (and_5[14], i0[14], i1[5]);
  and and_a14_b6 (and_6[14], i0[14], i1[6]);
  and and_a14_b7 (and_7[14], i0[14], i1[7]);
  and and_a14_b8 (and_8[14], i0[14], i1[8]);
  and and_a14_b9 (and_9[14], i0[14], i1[9]);
  and and_a15_b0 (and_0[15], i0[15], i1[0]);
  and and_a15_b1 (and_1[15], i0[15], i1[1]);
  and and_a15_b10 (and_10[15], i0[15], i1[10]);
  and and_a15_b11 (and_11[15], i0[15], i1[11]);
  and and_a15_b12 (and_12[15], i0[15], i1[12]);
  and and_a15_b13 (and_13[15], i0[15], i1[13]);
  and and_a15_b14 (and_14[15], i0[15], i1[14]);
  and and_a15_b15 (and_15[15], i0[15], i1[15]);
  and and_a15_b16 (and_16[15], i0[15], i1[16]);
  and and_a15_b17 (and_17[15], i0[15], i1[17]);
  and and_a15_b18 (and_18[15], i0[15], i1[18]);
  and and_a15_b19 (and_19[15], i0[15], i1[19]);
  and and_a15_b2 (and_2[15], i0[15], i1[2]);
  and and_a15_b20 (and_20[15], i0[15], i1[20]);
  and and_a15_b21 (and_21[15], i0[15], i1[21]);
  and and_a15_b22 (and_22[15], i0[15], i1[22]);
  and and_a15_b23 (and_23[15], i0[15], i1[23]);
  and and_a15_b24 (and_24[15], i0[15], i1[24]);
  and and_a15_b25 (and_25[15], i0[15], i1[25]);
  and and_a15_b26 (and_26[15], i0[15], i1[26]);
  and and_a15_b27 (and_27[15], i0[15], i1[27]);
  and and_a15_b28 (and_28[15], i0[15], i1[28]);
  and and_a15_b29 (and_29[15], i0[15], i1[29]);
  and and_a15_b3 (and_3[15], i0[15], i1[3]);
  and and_a15_b30 (and_30[15], i0[15], i1[30]);
  and and_a15_b31 (and_31[15], i0[15], i1[31]);
  and and_a15_b32 (nand_32[15], i0[15], i1[32]);
  and and_a15_b4 (and_4[15], i0[15], i1[4]);
  and and_a15_b5 (and_5[15], i0[15], i1[5]);
  and and_a15_b6 (and_6[15], i0[15], i1[6]);
  and and_a15_b7 (and_7[15], i0[15], i1[7]);
  and and_a15_b8 (and_8[15], i0[15], i1[8]);
  and and_a15_b9 (and_9[15], i0[15], i1[9]);
  and and_a16_b0 (and_0[16], i0[16], i1[0]);
  and and_a16_b1 (and_1[16], i0[16], i1[1]);
  and and_a16_b10 (and_10[16], i0[16], i1[10]);
  and and_a16_b11 (and_11[16], i0[16], i1[11]);
  and and_a16_b12 (and_12[16], i0[16], i1[12]);
  and and_a16_b13 (and_13[16], i0[16], i1[13]);
  and and_a16_b14 (and_14[16], i0[16], i1[14]);
  and and_a16_b15 (and_15[16], i0[16], i1[15]);
  and and_a16_b16 (and_16[16], i0[16], i1[16]);
  and and_a16_b17 (and_17[16], i0[16], i1[17]);
  and and_a16_b18 (and_18[16], i0[16], i1[18]);
  and and_a16_b19 (and_19[16], i0[16], i1[19]);
  and and_a16_b2 (and_2[16], i0[16], i1[2]);
  and and_a16_b20 (and_20[16], i0[16], i1[20]);
  and and_a16_b21 (and_21[16], i0[16], i1[21]);
  and and_a16_b22 (and_22[16], i0[16], i1[22]);
  and and_a16_b23 (and_23[16], i0[16], i1[23]);
  and and_a16_b24 (and_24[16], i0[16], i1[24]);
  and and_a16_b25 (and_25[16], i0[16], i1[25]);
  and and_a16_b26 (and_26[16], i0[16], i1[26]);
  and and_a16_b27 (and_27[16], i0[16], i1[27]);
  and and_a16_b28 (and_28[16], i0[16], i1[28]);
  and and_a16_b29 (and_29[16], i0[16], i1[29]);
  and and_a16_b3 (and_3[16], i0[16], i1[3]);
  and and_a16_b30 (and_30[16], i0[16], i1[30]);
  and and_a16_b31 (and_31[16], i0[16], i1[31]);
  and and_a16_b32 (nand_32[16], i0[16], i1[32]);
  and and_a16_b4 (and_4[16], i0[16], i1[4]);
  and and_a16_b5 (and_5[16], i0[16], i1[5]);
  and and_a16_b6 (and_6[16], i0[16], i1[6]);
  and and_a16_b7 (and_7[16], i0[16], i1[7]);
  and and_a16_b8 (and_8[16], i0[16], i1[8]);
  and and_a16_b9 (and_9[16], i0[16], i1[9]);
  and and_a17_b0 (and_0[17], i0[17], i1[0]);
  and and_a17_b1 (and_1[17], i0[17], i1[1]);
  and and_a17_b10 (and_10[17], i0[17], i1[10]);
  and and_a17_b11 (and_11[17], i0[17], i1[11]);
  and and_a17_b12 (and_12[17], i0[17], i1[12]);
  and and_a17_b13 (and_13[17], i0[17], i1[13]);
  and and_a17_b14 (and_14[17], i0[17], i1[14]);
  and and_a17_b15 (and_15[17], i0[17], i1[15]);
  and and_a17_b16 (and_16[17], i0[17], i1[16]);
  and and_a17_b17 (and_17[17], i0[17], i1[17]);
  and and_a17_b18 (and_18[17], i0[17], i1[18]);
  and and_a17_b19 (and_19[17], i0[17], i1[19]);
  and and_a17_b2 (and_2[17], i0[17], i1[2]);
  and and_a17_b20 (and_20[17], i0[17], i1[20]);
  and and_a17_b21 (and_21[17], i0[17], i1[21]);
  and and_a17_b22 (and_22[17], i0[17], i1[22]);
  and and_a17_b23 (and_23[17], i0[17], i1[23]);
  and and_a17_b24 (and_24[17], i0[17], i1[24]);
  and and_a17_b25 (and_25[17], i0[17], i1[25]);
  and and_a17_b26 (and_26[17], i0[17], i1[26]);
  and and_a17_b27 (and_27[17], i0[17], i1[27]);
  and and_a17_b28 (and_28[17], i0[17], i1[28]);
  and and_a17_b29 (and_29[17], i0[17], i1[29]);
  and and_a17_b3 (and_3[17], i0[17], i1[3]);
  and and_a17_b30 (and_30[17], i0[17], i1[30]);
  and and_a17_b31 (and_31[17], i0[17], i1[31]);
  and and_a17_b32 (nand_32[17], i0[17], i1[32]);
  and and_a17_b4 (and_4[17], i0[17], i1[4]);
  and and_a17_b5 (and_5[17], i0[17], i1[5]);
  and and_a17_b6 (and_6[17], i0[17], i1[6]);
  and and_a17_b7 (and_7[17], i0[17], i1[7]);
  and and_a17_b8 (and_8[17], i0[17], i1[8]);
  and and_a17_b9 (and_9[17], i0[17], i1[9]);
  and and_a18_b0 (and_0[18], i0[18], i1[0]);
  and and_a18_b1 (and_1[18], i0[18], i1[1]);
  and and_a18_b10 (and_10[18], i0[18], i1[10]);
  and and_a18_b11 (and_11[18], i0[18], i1[11]);
  and and_a18_b12 (and_12[18], i0[18], i1[12]);
  and and_a18_b13 (and_13[18], i0[18], i1[13]);
  and and_a18_b14 (and_14[18], i0[18], i1[14]);
  and and_a18_b15 (and_15[18], i0[18], i1[15]);
  and and_a18_b16 (and_16[18], i0[18], i1[16]);
  and and_a18_b17 (and_17[18], i0[18], i1[17]);
  and and_a18_b18 (and_18[18], i0[18], i1[18]);
  and and_a18_b19 (and_19[18], i0[18], i1[19]);
  and and_a18_b2 (and_2[18], i0[18], i1[2]);
  and and_a18_b20 (and_20[18], i0[18], i1[20]);
  and and_a18_b21 (and_21[18], i0[18], i1[21]);
  and and_a18_b22 (and_22[18], i0[18], i1[22]);
  and and_a18_b23 (and_23[18], i0[18], i1[23]);
  and and_a18_b24 (and_24[18], i0[18], i1[24]);
  and and_a18_b25 (and_25[18], i0[18], i1[25]);
  and and_a18_b26 (and_26[18], i0[18], i1[26]);
  and and_a18_b27 (and_27[18], i0[18], i1[27]);
  and and_a18_b28 (and_28[18], i0[18], i1[28]);
  and and_a18_b29 (and_29[18], i0[18], i1[29]);
  and and_a18_b3 (and_3[18], i0[18], i1[3]);
  and and_a18_b30 (and_30[18], i0[18], i1[30]);
  and and_a18_b31 (and_31[18], i0[18], i1[31]);
  and and_a18_b32 (nand_32[18], i0[18], i1[32]);
  and and_a18_b4 (and_4[18], i0[18], i1[4]);
  and and_a18_b5 (and_5[18], i0[18], i1[5]);
  and and_a18_b6 (and_6[18], i0[18], i1[6]);
  and and_a18_b7 (and_7[18], i0[18], i1[7]);
  and and_a18_b8 (and_8[18], i0[18], i1[8]);
  and and_a18_b9 (and_9[18], i0[18], i1[9]);
  and and_a19_b0 (and_0[19], i0[19], i1[0]);
  and and_a19_b1 (and_1[19], i0[19], i1[1]);
  and and_a19_b10 (and_10[19], i0[19], i1[10]);
  and and_a19_b11 (and_11[19], i0[19], i1[11]);
  and and_a19_b12 (and_12[19], i0[19], i1[12]);
  and and_a19_b13 (and_13[19], i0[19], i1[13]);
  and and_a19_b14 (and_14[19], i0[19], i1[14]);
  and and_a19_b15 (and_15[19], i0[19], i1[15]);
  and and_a19_b16 (and_16[19], i0[19], i1[16]);
  and and_a19_b17 (and_17[19], i0[19], i1[17]);
  and and_a19_b18 (and_18[19], i0[19], i1[18]);
  and and_a19_b19 (and_19[19], i0[19], i1[19]);
  and and_a19_b2 (and_2[19], i0[19], i1[2]);
  and and_a19_b20 (and_20[19], i0[19], i1[20]);
  and and_a19_b21 (and_21[19], i0[19], i1[21]);
  and and_a19_b22 (and_22[19], i0[19], i1[22]);
  and and_a19_b23 (and_23[19], i0[19], i1[23]);
  and and_a19_b24 (and_24[19], i0[19], i1[24]);
  and and_a19_b25 (and_25[19], i0[19], i1[25]);
  and and_a19_b26 (and_26[19], i0[19], i1[26]);
  and and_a19_b27 (and_27[19], i0[19], i1[27]);
  and and_a19_b28 (and_28[19], i0[19], i1[28]);
  and and_a19_b29 (and_29[19], i0[19], i1[29]);
  and and_a19_b3 (and_3[19], i0[19], i1[3]);
  and and_a19_b30 (and_30[19], i0[19], i1[30]);
  and and_a19_b31 (and_31[19], i0[19], i1[31]);
  and and_a19_b32 (nand_32[19], i0[19], i1[32]);
  and and_a19_b4 (and_4[19], i0[19], i1[4]);
  and and_a19_b5 (and_5[19], i0[19], i1[5]);
  and and_a19_b6 (and_6[19], i0[19], i1[6]);
  and and_a19_b7 (and_7[19], i0[19], i1[7]);
  and and_a19_b8 (and_8[19], i0[19], i1[8]);
  and and_a19_b9 (and_9[19], i0[19], i1[9]);
  and and_a1_b0 (and_0[1], i0[1], i1[0]);
  and and_a1_b1 (and_1[1], i0[1], i1[1]);
  and and_a1_b10 (and_10[1], i0[1], i1[10]);
  and and_a1_b11 (and_11[1], i0[1], i1[11]);
  and and_a1_b12 (and_12[1], i0[1], i1[12]);
  and and_a1_b13 (and_13[1], i0[1], i1[13]);
  and and_a1_b14 (and_14[1], i0[1], i1[14]);
  and and_a1_b15 (and_15[1], i0[1], i1[15]);
  and and_a1_b16 (and_16[1], i0[1], i1[16]);
  and and_a1_b17 (and_17[1], i0[1], i1[17]);
  and and_a1_b18 (and_18[1], i0[1], i1[18]);
  and and_a1_b19 (and_19[1], i0[1], i1[19]);
  and and_a1_b2 (and_2[1], i0[1], i1[2]);
  and and_a1_b20 (and_20[1], i0[1], i1[20]);
  and and_a1_b21 (and_21[1], i0[1], i1[21]);
  and and_a1_b22 (and_22[1], i0[1], i1[22]);
  and and_a1_b23 (and_23[1], i0[1], i1[23]);
  and and_a1_b24 (and_24[1], i0[1], i1[24]);
  and and_a1_b25 (and_25[1], i0[1], i1[25]);
  and and_a1_b26 (and_26[1], i0[1], i1[26]);
  and and_a1_b27 (and_27[1], i0[1], i1[27]);
  and and_a1_b28 (and_28[1], i0[1], i1[28]);
  and and_a1_b29 (and_29[1], i0[1], i1[29]);
  and and_a1_b3 (and_3[1], i0[1], i1[3]);
  and and_a1_b30 (and_30[1], i0[1], i1[30]);
  and and_a1_b31 (and_31[1], i0[1], i1[31]);
  and and_a1_b32 (nand_32[1], i0[1], i1[32]);
  and and_a1_b4 (and_4[1], i0[1], i1[4]);
  and and_a1_b5 (and_5[1], i0[1], i1[5]);
  and and_a1_b6 (and_6[1], i0[1], i1[6]);
  and and_a1_b7 (and_7[1], i0[1], i1[7]);
  and and_a1_b8 (and_8[1], i0[1], i1[8]);
  and and_a1_b9 (and_9[1], i0[1], i1[9]);
  and and_a20_b0 (and_0[20], i0[20], i1[0]);
  and and_a20_b1 (and_1[20], i0[20], i1[1]);
  and and_a20_b10 (and_10[20], i0[20], i1[10]);
  and and_a20_b11 (and_11[20], i0[20], i1[11]);
  and and_a20_b12 (and_12[20], i0[20], i1[12]);
  and and_a20_b13 (and_13[20], i0[20], i1[13]);
  and and_a20_b14 (and_14[20], i0[20], i1[14]);
  and and_a20_b15 (and_15[20], i0[20], i1[15]);
  and and_a20_b16 (and_16[20], i0[20], i1[16]);
  and and_a20_b17 (and_17[20], i0[20], i1[17]);
  and and_a20_b18 (and_18[20], i0[20], i1[18]);
  and and_a20_b19 (and_19[20], i0[20], i1[19]);
  and and_a20_b2 (and_2[20], i0[20], i1[2]);
  and and_a20_b20 (and_20[20], i0[20], i1[20]);
  and and_a20_b21 (and_21[20], i0[20], i1[21]);
  and and_a20_b22 (and_22[20], i0[20], i1[22]);
  and and_a20_b23 (and_23[20], i0[20], i1[23]);
  and and_a20_b24 (and_24[20], i0[20], i1[24]);
  and and_a20_b25 (and_25[20], i0[20], i1[25]);
  and and_a20_b26 (and_26[20], i0[20], i1[26]);
  and and_a20_b27 (and_27[20], i0[20], i1[27]);
  and and_a20_b28 (and_28[20], i0[20], i1[28]);
  and and_a20_b29 (and_29[20], i0[20], i1[29]);
  and and_a20_b3 (and_3[20], i0[20], i1[3]);
  and and_a20_b30 (and_30[20], i0[20], i1[30]);
  and and_a20_b31 (and_31[20], i0[20], i1[31]);
  and and_a20_b32 (nand_32[20], i0[20], i1[32]);
  and and_a20_b4 (and_4[20], i0[20], i1[4]);
  and and_a20_b5 (and_5[20], i0[20], i1[5]);
  and and_a20_b6 (and_6[20], i0[20], i1[6]);
  and and_a20_b7 (and_7[20], i0[20], i1[7]);
  and and_a20_b8 (and_8[20], i0[20], i1[8]);
  and and_a20_b9 (and_9[20], i0[20], i1[9]);
  and and_a21_b0 (and_0[21], i0[21], i1[0]);
  and and_a21_b1 (and_1[21], i0[21], i1[1]);
  and and_a21_b10 (and_10[21], i0[21], i1[10]);
  and and_a21_b11 (and_11[21], i0[21], i1[11]);
  and and_a21_b12 (and_12[21], i0[21], i1[12]);
  and and_a21_b13 (and_13[21], i0[21], i1[13]);
  and and_a21_b14 (and_14[21], i0[21], i1[14]);
  and and_a21_b15 (and_15[21], i0[21], i1[15]);
  and and_a21_b16 (and_16[21], i0[21], i1[16]);
  and and_a21_b17 (and_17[21], i0[21], i1[17]);
  and and_a21_b18 (and_18[21], i0[21], i1[18]);
  and and_a21_b19 (and_19[21], i0[21], i1[19]);
  and and_a21_b2 (and_2[21], i0[21], i1[2]);
  and and_a21_b20 (and_20[21], i0[21], i1[20]);
  and and_a21_b21 (and_21[21], i0[21], i1[21]);
  and and_a21_b22 (and_22[21], i0[21], i1[22]);
  and and_a21_b23 (and_23[21], i0[21], i1[23]);
  and and_a21_b24 (and_24[21], i0[21], i1[24]);
  and and_a21_b25 (and_25[21], i0[21], i1[25]);
  and and_a21_b26 (and_26[21], i0[21], i1[26]);
  and and_a21_b27 (and_27[21], i0[21], i1[27]);
  and and_a21_b28 (and_28[21], i0[21], i1[28]);
  and and_a21_b29 (and_29[21], i0[21], i1[29]);
  and and_a21_b3 (and_3[21], i0[21], i1[3]);
  and and_a21_b30 (and_30[21], i0[21], i1[30]);
  and and_a21_b31 (and_31[21], i0[21], i1[31]);
  and and_a21_b32 (nand_32[21], i0[21], i1[32]);
  and and_a21_b4 (and_4[21], i0[21], i1[4]);
  and and_a21_b5 (and_5[21], i0[21], i1[5]);
  and and_a21_b6 (and_6[21], i0[21], i1[6]);
  and and_a21_b7 (and_7[21], i0[21], i1[7]);
  and and_a21_b8 (and_8[21], i0[21], i1[8]);
  and and_a21_b9 (and_9[21], i0[21], i1[9]);
  and and_a22_b0 (and_0[22], i0[22], i1[0]);
  and and_a22_b1 (and_1[22], i0[22], i1[1]);
  and and_a22_b10 (and_10[22], i0[22], i1[10]);
  and and_a22_b11 (and_11[22], i0[22], i1[11]);
  and and_a22_b12 (and_12[22], i0[22], i1[12]);
  and and_a22_b13 (and_13[22], i0[22], i1[13]);
  and and_a22_b14 (and_14[22], i0[22], i1[14]);
  and and_a22_b15 (and_15[22], i0[22], i1[15]);
  and and_a22_b16 (and_16[22], i0[22], i1[16]);
  and and_a22_b17 (and_17[22], i0[22], i1[17]);
  and and_a22_b18 (and_18[22], i0[22], i1[18]);
  and and_a22_b19 (and_19[22], i0[22], i1[19]);
  and and_a22_b2 (and_2[22], i0[22], i1[2]);
  and and_a22_b20 (and_20[22], i0[22], i1[20]);
  and and_a22_b21 (and_21[22], i0[22], i1[21]);
  and and_a22_b22 (and_22[22], i0[22], i1[22]);
  and and_a22_b23 (and_23[22], i0[22], i1[23]);
  and and_a22_b24 (and_24[22], i0[22], i1[24]);
  and and_a22_b25 (and_25[22], i0[22], i1[25]);
  and and_a22_b26 (and_26[22], i0[22], i1[26]);
  and and_a22_b27 (and_27[22], i0[22], i1[27]);
  and and_a22_b28 (and_28[22], i0[22], i1[28]);
  and and_a22_b29 (and_29[22], i0[22], i1[29]);
  and and_a22_b3 (and_3[22], i0[22], i1[3]);
  and and_a22_b30 (and_30[22], i0[22], i1[30]);
  and and_a22_b31 (and_31[22], i0[22], i1[31]);
  and and_a22_b32 (nand_32[22], i0[22], i1[32]);
  and and_a22_b4 (and_4[22], i0[22], i1[4]);
  and and_a22_b5 (and_5[22], i0[22], i1[5]);
  and and_a22_b6 (and_6[22], i0[22], i1[6]);
  and and_a22_b7 (and_7[22], i0[22], i1[7]);
  and and_a22_b8 (and_8[22], i0[22], i1[8]);
  and and_a22_b9 (and_9[22], i0[22], i1[9]);
  and and_a23_b0 (and_0[23], i0[23], i1[0]);
  and and_a23_b1 (and_1[23], i0[23], i1[1]);
  and and_a23_b10 (and_10[23], i0[23], i1[10]);
  and and_a23_b11 (and_11[23], i0[23], i1[11]);
  and and_a23_b12 (and_12[23], i0[23], i1[12]);
  and and_a23_b13 (and_13[23], i0[23], i1[13]);
  and and_a23_b14 (and_14[23], i0[23], i1[14]);
  and and_a23_b15 (and_15[23], i0[23], i1[15]);
  and and_a23_b16 (and_16[23], i0[23], i1[16]);
  and and_a23_b17 (and_17[23], i0[23], i1[17]);
  and and_a23_b18 (and_18[23], i0[23], i1[18]);
  and and_a23_b19 (and_19[23], i0[23], i1[19]);
  and and_a23_b2 (and_2[23], i0[23], i1[2]);
  and and_a23_b20 (and_20[23], i0[23], i1[20]);
  and and_a23_b21 (and_21[23], i0[23], i1[21]);
  and and_a23_b22 (and_22[23], i0[23], i1[22]);
  and and_a23_b23 (and_23[23], i0[23], i1[23]);
  and and_a23_b24 (and_24[23], i0[23], i1[24]);
  and and_a23_b25 (and_25[23], i0[23], i1[25]);
  and and_a23_b26 (and_26[23], i0[23], i1[26]);
  and and_a23_b27 (and_27[23], i0[23], i1[27]);
  and and_a23_b28 (and_28[23], i0[23], i1[28]);
  and and_a23_b29 (and_29[23], i0[23], i1[29]);
  and and_a23_b3 (and_3[23], i0[23], i1[3]);
  and and_a23_b30 (and_30[23], i0[23], i1[30]);
  and and_a23_b31 (and_31[23], i0[23], i1[31]);
  and and_a23_b32 (nand_32[23], i0[23], i1[32]);
  and and_a23_b4 (and_4[23], i0[23], i1[4]);
  and and_a23_b5 (and_5[23], i0[23], i1[5]);
  and and_a23_b6 (and_6[23], i0[23], i1[6]);
  and and_a23_b7 (and_7[23], i0[23], i1[7]);
  and and_a23_b8 (and_8[23], i0[23], i1[8]);
  and and_a23_b9 (and_9[23], i0[23], i1[9]);
  and and_a24_b0 (and_0[24], i0[24], i1[0]);
  and and_a24_b1 (and_1[24], i0[24], i1[1]);
  and and_a24_b10 (and_10[24], i0[24], i1[10]);
  and and_a24_b11 (and_11[24], i0[24], i1[11]);
  and and_a24_b12 (and_12[24], i0[24], i1[12]);
  and and_a24_b13 (and_13[24], i0[24], i1[13]);
  and and_a24_b14 (and_14[24], i0[24], i1[14]);
  and and_a24_b15 (and_15[24], i0[24], i1[15]);
  and and_a24_b16 (and_16[24], i0[24], i1[16]);
  and and_a24_b17 (and_17[24], i0[24], i1[17]);
  and and_a24_b18 (and_18[24], i0[24], i1[18]);
  and and_a24_b19 (and_19[24], i0[24], i1[19]);
  and and_a24_b2 (and_2[24], i0[24], i1[2]);
  and and_a24_b20 (and_20[24], i0[24], i1[20]);
  and and_a24_b21 (and_21[24], i0[24], i1[21]);
  and and_a24_b22 (and_22[24], i0[24], i1[22]);
  and and_a24_b23 (and_23[24], i0[24], i1[23]);
  and and_a24_b24 (and_24[24], i0[24], i1[24]);
  and and_a24_b25 (and_25[24], i0[24], i1[25]);
  and and_a24_b26 (and_26[24], i0[24], i1[26]);
  and and_a24_b27 (and_27[24], i0[24], i1[27]);
  and and_a24_b28 (and_28[24], i0[24], i1[28]);
  and and_a24_b29 (and_29[24], i0[24], i1[29]);
  and and_a24_b3 (and_3[24], i0[24], i1[3]);
  and and_a24_b30 (and_30[24], i0[24], i1[30]);
  and and_a24_b31 (and_31[24], i0[24], i1[31]);
  and and_a24_b32 (nand_32[24], i0[24], i1[32]);
  and and_a24_b4 (and_4[24], i0[24], i1[4]);
  and and_a24_b5 (and_5[24], i0[24], i1[5]);
  and and_a24_b6 (and_6[24], i0[24], i1[6]);
  and and_a24_b7 (and_7[24], i0[24], i1[7]);
  and and_a24_b8 (and_8[24], i0[24], i1[8]);
  and and_a24_b9 (and_9[24], i0[24], i1[9]);
  and and_a25_b0 (and_0[25], i0[25], i1[0]);
  and and_a25_b1 (and_1[25], i0[25], i1[1]);
  and and_a25_b10 (and_10[25], i0[25], i1[10]);
  and and_a25_b11 (and_11[25], i0[25], i1[11]);
  and and_a25_b12 (and_12[25], i0[25], i1[12]);
  and and_a25_b13 (and_13[25], i0[25], i1[13]);
  and and_a25_b14 (and_14[25], i0[25], i1[14]);
  and and_a25_b15 (and_15[25], i0[25], i1[15]);
  and and_a25_b16 (and_16[25], i0[25], i1[16]);
  and and_a25_b17 (and_17[25], i0[25], i1[17]);
  and and_a25_b18 (and_18[25], i0[25], i1[18]);
  and and_a25_b19 (and_19[25], i0[25], i1[19]);
  and and_a25_b2 (and_2[25], i0[25], i1[2]);
  and and_a25_b20 (and_20[25], i0[25], i1[20]);
  and and_a25_b21 (and_21[25], i0[25], i1[21]);
  and and_a25_b22 (and_22[25], i0[25], i1[22]);
  and and_a25_b23 (and_23[25], i0[25], i1[23]);
  and and_a25_b24 (and_24[25], i0[25], i1[24]);
  and and_a25_b25 (and_25[25], i0[25], i1[25]);
  and and_a25_b26 (and_26[25], i0[25], i1[26]);
  and and_a25_b27 (and_27[25], i0[25], i1[27]);
  and and_a25_b28 (and_28[25], i0[25], i1[28]);
  and and_a25_b29 (and_29[25], i0[25], i1[29]);
  and and_a25_b3 (and_3[25], i0[25], i1[3]);
  and and_a25_b30 (and_30[25], i0[25], i1[30]);
  and and_a25_b31 (and_31[25], i0[25], i1[31]);
  and and_a25_b32 (nand_32[25], i0[25], i1[32]);
  and and_a25_b4 (and_4[25], i0[25], i1[4]);
  and and_a25_b5 (and_5[25], i0[25], i1[5]);
  and and_a25_b6 (and_6[25], i0[25], i1[6]);
  and and_a25_b7 (and_7[25], i0[25], i1[7]);
  and and_a25_b8 (and_8[25], i0[25], i1[8]);
  and and_a25_b9 (and_9[25], i0[25], i1[9]);
  and and_a26_b0 (and_0[26], i0[26], i1[0]);
  and and_a26_b1 (and_1[26], i0[26], i1[1]);
  and and_a26_b10 (and_10[26], i0[26], i1[10]);
  and and_a26_b11 (and_11[26], i0[26], i1[11]);
  and and_a26_b12 (and_12[26], i0[26], i1[12]);
  and and_a26_b13 (and_13[26], i0[26], i1[13]);
  and and_a26_b14 (and_14[26], i0[26], i1[14]);
  and and_a26_b15 (and_15[26], i0[26], i1[15]);
  and and_a26_b16 (and_16[26], i0[26], i1[16]);
  and and_a26_b17 (and_17[26], i0[26], i1[17]);
  and and_a26_b18 (and_18[26], i0[26], i1[18]);
  and and_a26_b19 (and_19[26], i0[26], i1[19]);
  and and_a26_b2 (and_2[26], i0[26], i1[2]);
  and and_a26_b20 (and_20[26], i0[26], i1[20]);
  and and_a26_b21 (and_21[26], i0[26], i1[21]);
  and and_a26_b22 (and_22[26], i0[26], i1[22]);
  and and_a26_b23 (and_23[26], i0[26], i1[23]);
  and and_a26_b24 (and_24[26], i0[26], i1[24]);
  and and_a26_b25 (and_25[26], i0[26], i1[25]);
  and and_a26_b26 (and_26[26], i0[26], i1[26]);
  and and_a26_b27 (and_27[26], i0[26], i1[27]);
  and and_a26_b28 (and_28[26], i0[26], i1[28]);
  and and_a26_b29 (and_29[26], i0[26], i1[29]);
  and and_a26_b3 (and_3[26], i0[26], i1[3]);
  and and_a26_b30 (and_30[26], i0[26], i1[30]);
  and and_a26_b31 (and_31[26], i0[26], i1[31]);
  and and_a26_b32 (nand_32[26], i0[26], i1[32]);
  and and_a26_b4 (and_4[26], i0[26], i1[4]);
  and and_a26_b5 (and_5[26], i0[26], i1[5]);
  and and_a26_b6 (and_6[26], i0[26], i1[6]);
  and and_a26_b7 (and_7[26], i0[26], i1[7]);
  and and_a26_b8 (and_8[26], i0[26], i1[8]);
  and and_a26_b9 (and_9[26], i0[26], i1[9]);
  and and_a27_b0 (and_0[27], i0[27], i1[0]);
  and and_a27_b1 (and_1[27], i0[27], i1[1]);
  and and_a27_b10 (and_10[27], i0[27], i1[10]);
  and and_a27_b11 (and_11[27], i0[27], i1[11]);
  and and_a27_b12 (and_12[27], i0[27], i1[12]);
  and and_a27_b13 (and_13[27], i0[27], i1[13]);
  and and_a27_b14 (and_14[27], i0[27], i1[14]);
  and and_a27_b15 (and_15[27], i0[27], i1[15]);
  and and_a27_b16 (and_16[27], i0[27], i1[16]);
  and and_a27_b17 (and_17[27], i0[27], i1[17]);
  and and_a27_b18 (and_18[27], i0[27], i1[18]);
  and and_a27_b19 (and_19[27], i0[27], i1[19]);
  and and_a27_b2 (and_2[27], i0[27], i1[2]);
  and and_a27_b20 (and_20[27], i0[27], i1[20]);
  and and_a27_b21 (and_21[27], i0[27], i1[21]);
  and and_a27_b22 (and_22[27], i0[27], i1[22]);
  and and_a27_b23 (and_23[27], i0[27], i1[23]);
  and and_a27_b24 (and_24[27], i0[27], i1[24]);
  and and_a27_b25 (and_25[27], i0[27], i1[25]);
  and and_a27_b26 (and_26[27], i0[27], i1[26]);
  and and_a27_b27 (and_27[27], i0[27], i1[27]);
  and and_a27_b28 (and_28[27], i0[27], i1[28]);
  and and_a27_b29 (and_29[27], i0[27], i1[29]);
  and and_a27_b3 (and_3[27], i0[27], i1[3]);
  and and_a27_b30 (and_30[27], i0[27], i1[30]);
  and and_a27_b31 (and_31[27], i0[27], i1[31]);
  and and_a27_b32 (nand_32[27], i0[27], i1[32]);
  and and_a27_b4 (and_4[27], i0[27], i1[4]);
  and and_a27_b5 (and_5[27], i0[27], i1[5]);
  and and_a27_b6 (and_6[27], i0[27], i1[6]);
  and and_a27_b7 (and_7[27], i0[27], i1[7]);
  and and_a27_b8 (and_8[27], i0[27], i1[8]);
  and and_a27_b9 (and_9[27], i0[27], i1[9]);
  and and_a28_b0 (and_0[28], i0[28], i1[0]);
  and and_a28_b1 (and_1[28], i0[28], i1[1]);
  and and_a28_b10 (and_10[28], i0[28], i1[10]);
  and and_a28_b11 (and_11[28], i0[28], i1[11]);
  and and_a28_b12 (and_12[28], i0[28], i1[12]);
  and and_a28_b13 (and_13[28], i0[28], i1[13]);
  and and_a28_b14 (and_14[28], i0[28], i1[14]);
  and and_a28_b15 (and_15[28], i0[28], i1[15]);
  and and_a28_b16 (and_16[28], i0[28], i1[16]);
  and and_a28_b17 (and_17[28], i0[28], i1[17]);
  and and_a28_b18 (and_18[28], i0[28], i1[18]);
  and and_a28_b19 (and_19[28], i0[28], i1[19]);
  and and_a28_b2 (and_2[28], i0[28], i1[2]);
  and and_a28_b20 (and_20[28], i0[28], i1[20]);
  and and_a28_b21 (and_21[28], i0[28], i1[21]);
  and and_a28_b22 (and_22[28], i0[28], i1[22]);
  and and_a28_b23 (and_23[28], i0[28], i1[23]);
  and and_a28_b24 (and_24[28], i0[28], i1[24]);
  and and_a28_b25 (and_25[28], i0[28], i1[25]);
  and and_a28_b26 (and_26[28], i0[28], i1[26]);
  and and_a28_b27 (and_27[28], i0[28], i1[27]);
  and and_a28_b28 (and_28[28], i0[28], i1[28]);
  and and_a28_b29 (and_29[28], i0[28], i1[29]);
  and and_a28_b3 (and_3[28], i0[28], i1[3]);
  and and_a28_b30 (and_30[28], i0[28], i1[30]);
  and and_a28_b31 (and_31[28], i0[28], i1[31]);
  and and_a28_b32 (nand_32[28], i0[28], i1[32]);
  and and_a28_b4 (and_4[28], i0[28], i1[4]);
  and and_a28_b5 (and_5[28], i0[28], i1[5]);
  and and_a28_b6 (and_6[28], i0[28], i1[6]);
  and and_a28_b7 (and_7[28], i0[28], i1[7]);
  and and_a28_b8 (and_8[28], i0[28], i1[8]);
  and and_a28_b9 (and_9[28], i0[28], i1[9]);
  and and_a29_b0 (and_0[29], i0[29], i1[0]);
  and and_a29_b1 (and_1[29], i0[29], i1[1]);
  and and_a29_b10 (and_10[29], i0[29], i1[10]);
  and and_a29_b11 (and_11[29], i0[29], i1[11]);
  and and_a29_b12 (and_12[29], i0[29], i1[12]);
  and and_a29_b13 (and_13[29], i0[29], i1[13]);
  and and_a29_b14 (and_14[29], i0[29], i1[14]);
  and and_a29_b15 (and_15[29], i0[29], i1[15]);
  and and_a29_b16 (and_16[29], i0[29], i1[16]);
  and and_a29_b17 (and_17[29], i0[29], i1[17]);
  and and_a29_b18 (and_18[29], i0[29], i1[18]);
  and and_a29_b19 (and_19[29], i0[29], i1[19]);
  and and_a29_b2 (and_2[29], i0[29], i1[2]);
  and and_a29_b20 (and_20[29], i0[29], i1[20]);
  and and_a29_b21 (and_21[29], i0[29], i1[21]);
  and and_a29_b22 (and_22[29], i0[29], i1[22]);
  and and_a29_b23 (and_23[29], i0[29], i1[23]);
  and and_a29_b24 (and_24[29], i0[29], i1[24]);
  and and_a29_b25 (and_25[29], i0[29], i1[25]);
  and and_a29_b26 (and_26[29], i0[29], i1[26]);
  and and_a29_b27 (and_27[29], i0[29], i1[27]);
  and and_a29_b28 (and_28[29], i0[29], i1[28]);
  and and_a29_b29 (and_29[29], i0[29], i1[29]);
  and and_a29_b3 (and_3[29], i0[29], i1[3]);
  and and_a29_b30 (and_30[29], i0[29], i1[30]);
  and and_a29_b31 (and_31[29], i0[29], i1[31]);
  and and_a29_b32 (nand_32[29], i0[29], i1[32]);
  and and_a29_b4 (and_4[29], i0[29], i1[4]);
  and and_a29_b5 (and_5[29], i0[29], i1[5]);
  and and_a29_b6 (and_6[29], i0[29], i1[6]);
  and and_a29_b7 (and_7[29], i0[29], i1[7]);
  and and_a29_b8 (and_8[29], i0[29], i1[8]);
  and and_a29_b9 (and_9[29], i0[29], i1[9]);
  and and_a2_b0 (and_0[2], i0[2], i1[0]);
  and and_a2_b1 (and_1[2], i0[2], i1[1]);
  and and_a2_b10 (and_10[2], i0[2], i1[10]);
  and and_a2_b11 (and_11[2], i0[2], i1[11]);
  and and_a2_b12 (and_12[2], i0[2], i1[12]);
  and and_a2_b13 (and_13[2], i0[2], i1[13]);
  and and_a2_b14 (and_14[2], i0[2], i1[14]);
  and and_a2_b15 (and_15[2], i0[2], i1[15]);
  and and_a2_b16 (and_16[2], i0[2], i1[16]);
  and and_a2_b17 (and_17[2], i0[2], i1[17]);
  and and_a2_b18 (and_18[2], i0[2], i1[18]);
  and and_a2_b19 (and_19[2], i0[2], i1[19]);
  and and_a2_b2 (and_2[2], i0[2], i1[2]);
  and and_a2_b20 (and_20[2], i0[2], i1[20]);
  and and_a2_b21 (and_21[2], i0[2], i1[21]);
  and and_a2_b22 (and_22[2], i0[2], i1[22]);
  and and_a2_b23 (and_23[2], i0[2], i1[23]);
  and and_a2_b24 (and_24[2], i0[2], i1[24]);
  and and_a2_b25 (and_25[2], i0[2], i1[25]);
  and and_a2_b26 (and_26[2], i0[2], i1[26]);
  and and_a2_b27 (and_27[2], i0[2], i1[27]);
  and and_a2_b28 (and_28[2], i0[2], i1[28]);
  and and_a2_b29 (and_29[2], i0[2], i1[29]);
  and and_a2_b3 (and_3[2], i0[2], i1[3]);
  and and_a2_b30 (and_30[2], i0[2], i1[30]);
  and and_a2_b31 (and_31[2], i0[2], i1[31]);
  and and_a2_b32 (nand_32[2], i0[2], i1[32]);
  and and_a2_b4 (and_4[2], i0[2], i1[4]);
  and and_a2_b5 (and_5[2], i0[2], i1[5]);
  and and_a2_b6 (and_6[2], i0[2], i1[6]);
  and and_a2_b7 (and_7[2], i0[2], i1[7]);
  and and_a2_b8 (and_8[2], i0[2], i1[8]);
  and and_a2_b9 (and_9[2], i0[2], i1[9]);
  and and_a30_b0 (and_0[30], i0[30], i1[0]);
  and and_a30_b1 (and_1[30], i0[30], i1[1]);
  and and_a30_b10 (and_10[30], i0[30], i1[10]);
  and and_a30_b11 (and_11[30], i0[30], i1[11]);
  and and_a30_b12 (and_12[30], i0[30], i1[12]);
  and and_a30_b13 (and_13[30], i0[30], i1[13]);
  and and_a30_b14 (and_14[30], i0[30], i1[14]);
  and and_a30_b15 (and_15[30], i0[30], i1[15]);
  and and_a30_b16 (and_16[30], i0[30], i1[16]);
  and and_a30_b17 (and_17[30], i0[30], i1[17]);
  and and_a30_b18 (and_18[30], i0[30], i1[18]);
  and and_a30_b19 (and_19[30], i0[30], i1[19]);
  and and_a30_b2 (and_2[30], i0[30], i1[2]);
  and and_a30_b20 (and_20[30], i0[30], i1[20]);
  and and_a30_b21 (and_21[30], i0[30], i1[21]);
  and and_a30_b22 (and_22[30], i0[30], i1[22]);
  and and_a30_b23 (and_23[30], i0[30], i1[23]);
  and and_a30_b24 (and_24[30], i0[30], i1[24]);
  and and_a30_b25 (and_25[30], i0[30], i1[25]);
  and and_a30_b26 (and_26[30], i0[30], i1[26]);
  and and_a30_b27 (and_27[30], i0[30], i1[27]);
  and and_a30_b28 (and_28[30], i0[30], i1[28]);
  and and_a30_b29 (and_29[30], i0[30], i1[29]);
  and and_a30_b3 (and_3[30], i0[30], i1[3]);
  and and_a30_b30 (and_30[30], i0[30], i1[30]);
  and and_a30_b31 (and_31[30], i0[30], i1[31]);
  and and_a30_b32 (nand_32[30], i0[30], i1[32]);
  and and_a30_b4 (and_4[30], i0[30], i1[4]);
  and and_a30_b5 (and_5[30], i0[30], i1[5]);
  and and_a30_b6 (and_6[30], i0[30], i1[6]);
  and and_a30_b7 (and_7[30], i0[30], i1[7]);
  and and_a30_b8 (and_8[30], i0[30], i1[8]);
  and and_a30_b9 (and_9[30], i0[30], i1[9]);
  and and_a31_b0 (nand_0[31], i0[31], i1[0]);
  and and_a31_b1 (nand_1[31], i0[31], i1[1]);
  and and_a31_b10 (nand_10[31], i0[31], i1[10]);
  and and_a31_b11 (nand_11[31], i0[31], i1[11]);
  and and_a31_b12 (nand_12[31], i0[31], i1[12]);
  and and_a31_b13 (nand_13[31], i0[31], i1[13]);
  and and_a31_b14 (nand_14[31], i0[31], i1[14]);
  and and_a31_b15 (nand_15[31], i0[31], i1[15]);
  and and_a31_b16 (nand_16[31], i0[31], i1[16]);
  and and_a31_b17 (nand_17[31], i0[31], i1[17]);
  and and_a31_b18 (nand_18[31], i0[31], i1[18]);
  and and_a31_b19 (nand_19[31], i0[31], i1[19]);
  and and_a31_b2 (nand_2[31], i0[31], i1[2]);
  and and_a31_b20 (nand_20[31], i0[31], i1[20]);
  and and_a31_b21 (nand_21[31], i0[31], i1[21]);
  and and_a31_b22 (nand_22[31], i0[31], i1[22]);
  and and_a31_b23 (nand_23[31], i0[31], i1[23]);
  and and_a31_b24 (nand_24[31], i0[31], i1[24]);
  and and_a31_b25 (nand_25[31], i0[31], i1[25]);
  and and_a31_b26 (nand_26[31], i0[31], i1[26]);
  and and_a31_b27 (nand_27[31], i0[31], i1[27]);
  and and_a31_b28 (nand_28[31], i0[31], i1[28]);
  and and_a31_b29 (nand_29[31], i0[31], i1[29]);
  and and_a31_b3 (nand_3[31], i0[31], i1[3]);
  and and_a31_b30 (nand_30[31], i0[31], i1[30]);
  and and_a31_b31 (nand_31[31], i0[31], i1[31]);
  and and_a31_b32 (and_32[31], i0[31], i1[32]);
  and and_a31_b4 (nand_4[31], i0[31], i1[4]);
  and and_a31_b5 (nand_5[31], i0[31], i1[5]);
  and and_a31_b6 (nand_6[31], i0[31], i1[6]);
  and and_a31_b7 (nand_7[31], i0[31], i1[7]);
  and and_a31_b8 (nand_8[31], i0[31], i1[8]);
  and and_a31_b9 (nand_9[31], i0[31], i1[9]);
  and and_a3_b0 (and_0[3], i0[3], i1[0]);
  and and_a3_b1 (and_1[3], i0[3], i1[1]);
  and and_a3_b10 (and_10[3], i0[3], i1[10]);
  and and_a3_b11 (and_11[3], i0[3], i1[11]);
  and and_a3_b12 (and_12[3], i0[3], i1[12]);
  and and_a3_b13 (and_13[3], i0[3], i1[13]);
  and and_a3_b14 (and_14[3], i0[3], i1[14]);
  and and_a3_b15 (and_15[3], i0[3], i1[15]);
  and and_a3_b16 (and_16[3], i0[3], i1[16]);
  and and_a3_b17 (and_17[3], i0[3], i1[17]);
  and and_a3_b18 (and_18[3], i0[3], i1[18]);
  and and_a3_b19 (and_19[3], i0[3], i1[19]);
  and and_a3_b2 (and_2[3], i0[3], i1[2]);
  and and_a3_b20 (and_20[3], i0[3], i1[20]);
  and and_a3_b21 (and_21[3], i0[3], i1[21]);
  and and_a3_b22 (and_22[3], i0[3], i1[22]);
  and and_a3_b23 (and_23[3], i0[3], i1[23]);
  and and_a3_b24 (and_24[3], i0[3], i1[24]);
  and and_a3_b25 (and_25[3], i0[3], i1[25]);
  and and_a3_b26 (and_26[3], i0[3], i1[26]);
  and and_a3_b27 (and_27[3], i0[3], i1[27]);
  and and_a3_b28 (and_28[3], i0[3], i1[28]);
  and and_a3_b29 (and_29[3], i0[3], i1[29]);
  and and_a3_b3 (and_3[3], i0[3], i1[3]);
  and and_a3_b30 (and_30[3], i0[3], i1[30]);
  and and_a3_b31 (and_31[3], i0[3], i1[31]);
  and and_a3_b32 (nand_32[3], i0[3], i1[32]);
  and and_a3_b4 (and_4[3], i0[3], i1[4]);
  and and_a3_b5 (and_5[3], i0[3], i1[5]);
  and and_a3_b6 (and_6[3], i0[3], i1[6]);
  and and_a3_b7 (and_7[3], i0[3], i1[7]);
  and and_a3_b8 (and_8[3], i0[3], i1[8]);
  and and_a3_b9 (and_9[3], i0[3], i1[9]);
  and and_a4_b0 (and_0[4], i0[4], i1[0]);
  and and_a4_b1 (and_1[4], i0[4], i1[1]);
  and and_a4_b10 (and_10[4], i0[4], i1[10]);
  and and_a4_b11 (and_11[4], i0[4], i1[11]);
  and and_a4_b12 (and_12[4], i0[4], i1[12]);
  and and_a4_b13 (and_13[4], i0[4], i1[13]);
  and and_a4_b14 (and_14[4], i0[4], i1[14]);
  and and_a4_b15 (and_15[4], i0[4], i1[15]);
  and and_a4_b16 (and_16[4], i0[4], i1[16]);
  and and_a4_b17 (and_17[4], i0[4], i1[17]);
  and and_a4_b18 (and_18[4], i0[4], i1[18]);
  and and_a4_b19 (and_19[4], i0[4], i1[19]);
  and and_a4_b2 (and_2[4], i0[4], i1[2]);
  and and_a4_b20 (and_20[4], i0[4], i1[20]);
  and and_a4_b21 (and_21[4], i0[4], i1[21]);
  and and_a4_b22 (and_22[4], i0[4], i1[22]);
  and and_a4_b23 (and_23[4], i0[4], i1[23]);
  and and_a4_b24 (and_24[4], i0[4], i1[24]);
  and and_a4_b25 (and_25[4], i0[4], i1[25]);
  and and_a4_b26 (and_26[4], i0[4], i1[26]);
  and and_a4_b27 (and_27[4], i0[4], i1[27]);
  and and_a4_b28 (and_28[4], i0[4], i1[28]);
  and and_a4_b29 (and_29[4], i0[4], i1[29]);
  and and_a4_b3 (and_3[4], i0[4], i1[3]);
  and and_a4_b30 (and_30[4], i0[4], i1[30]);
  and and_a4_b31 (and_31[4], i0[4], i1[31]);
  and and_a4_b32 (nand_32[4], i0[4], i1[32]);
  and and_a4_b4 (and_4[4], i0[4], i1[4]);
  and and_a4_b5 (and_5[4], i0[4], i1[5]);
  and and_a4_b6 (and_6[4], i0[4], i1[6]);
  and and_a4_b7 (and_7[4], i0[4], i1[7]);
  and and_a4_b8 (and_8[4], i0[4], i1[8]);
  and and_a4_b9 (and_9[4], i0[4], i1[9]);
  and and_a5_b0 (and_0[5], i0[5], i1[0]);
  and and_a5_b1 (and_1[5], i0[5], i1[1]);
  and and_a5_b10 (and_10[5], i0[5], i1[10]);
  and and_a5_b11 (and_11[5], i0[5], i1[11]);
  and and_a5_b12 (and_12[5], i0[5], i1[12]);
  and and_a5_b13 (and_13[5], i0[5], i1[13]);
  and and_a5_b14 (and_14[5], i0[5], i1[14]);
  and and_a5_b15 (and_15[5], i0[5], i1[15]);
  and and_a5_b16 (and_16[5], i0[5], i1[16]);
  and and_a5_b17 (and_17[5], i0[5], i1[17]);
  and and_a5_b18 (and_18[5], i0[5], i1[18]);
  and and_a5_b19 (and_19[5], i0[5], i1[19]);
  and and_a5_b2 (and_2[5], i0[5], i1[2]);
  and and_a5_b20 (and_20[5], i0[5], i1[20]);
  and and_a5_b21 (and_21[5], i0[5], i1[21]);
  and and_a5_b22 (and_22[5], i0[5], i1[22]);
  and and_a5_b23 (and_23[5], i0[5], i1[23]);
  and and_a5_b24 (and_24[5], i0[5], i1[24]);
  and and_a5_b25 (and_25[5], i0[5], i1[25]);
  and and_a5_b26 (and_26[5], i0[5], i1[26]);
  and and_a5_b27 (and_27[5], i0[5], i1[27]);
  and and_a5_b28 (and_28[5], i0[5], i1[28]);
  and and_a5_b29 (and_29[5], i0[5], i1[29]);
  and and_a5_b3 (and_3[5], i0[5], i1[3]);
  and and_a5_b30 (and_30[5], i0[5], i1[30]);
  and and_a5_b31 (and_31[5], i0[5], i1[31]);
  and and_a5_b32 (nand_32[5], i0[5], i1[32]);
  and and_a5_b4 (and_4[5], i0[5], i1[4]);
  and and_a5_b5 (and_5[5], i0[5], i1[5]);
  and and_a5_b6 (and_6[5], i0[5], i1[6]);
  and and_a5_b7 (and_7[5], i0[5], i1[7]);
  and and_a5_b8 (and_8[5], i0[5], i1[8]);
  and and_a5_b9 (and_9[5], i0[5], i1[9]);
  and and_a6_b0 (and_0[6], i0[6], i1[0]);
  and and_a6_b1 (and_1[6], i0[6], i1[1]);
  and and_a6_b10 (and_10[6], i0[6], i1[10]);
  and and_a6_b11 (and_11[6], i0[6], i1[11]);
  and and_a6_b12 (and_12[6], i0[6], i1[12]);
  and and_a6_b13 (and_13[6], i0[6], i1[13]);
  and and_a6_b14 (and_14[6], i0[6], i1[14]);
  and and_a6_b15 (and_15[6], i0[6], i1[15]);
  and and_a6_b16 (and_16[6], i0[6], i1[16]);
  and and_a6_b17 (and_17[6], i0[6], i1[17]);
  and and_a6_b18 (and_18[6], i0[6], i1[18]);
  and and_a6_b19 (and_19[6], i0[6], i1[19]);
  and and_a6_b2 (and_2[6], i0[6], i1[2]);
  and and_a6_b20 (and_20[6], i0[6], i1[20]);
  and and_a6_b21 (and_21[6], i0[6], i1[21]);
  and and_a6_b22 (and_22[6], i0[6], i1[22]);
  and and_a6_b23 (and_23[6], i0[6], i1[23]);
  and and_a6_b24 (and_24[6], i0[6], i1[24]);
  and and_a6_b25 (and_25[6], i0[6], i1[25]);
  and and_a6_b26 (and_26[6], i0[6], i1[26]);
  and and_a6_b27 (and_27[6], i0[6], i1[27]);
  and and_a6_b28 (and_28[6], i0[6], i1[28]);
  and and_a6_b29 (and_29[6], i0[6], i1[29]);
  and and_a6_b3 (and_3[6], i0[6], i1[3]);
  and and_a6_b30 (and_30[6], i0[6], i1[30]);
  and and_a6_b31 (and_31[6], i0[6], i1[31]);
  and and_a6_b32 (nand_32[6], i0[6], i1[32]);
  and and_a6_b4 (and_4[6], i0[6], i1[4]);
  and and_a6_b5 (and_5[6], i0[6], i1[5]);
  and and_a6_b6 (and_6[6], i0[6], i1[6]);
  and and_a6_b7 (and_7[6], i0[6], i1[7]);
  and and_a6_b8 (and_8[6], i0[6], i1[8]);
  and and_a6_b9 (and_9[6], i0[6], i1[9]);
  and and_a7_b0 (and_0[7], i0[7], i1[0]);
  and and_a7_b1 (and_1[7], i0[7], i1[1]);
  and and_a7_b10 (and_10[7], i0[7], i1[10]);
  and and_a7_b11 (and_11[7], i0[7], i1[11]);
  and and_a7_b12 (and_12[7], i0[7], i1[12]);
  and and_a7_b13 (and_13[7], i0[7], i1[13]);
  and and_a7_b14 (and_14[7], i0[7], i1[14]);
  and and_a7_b15 (and_15[7], i0[7], i1[15]);
  and and_a7_b16 (and_16[7], i0[7], i1[16]);
  and and_a7_b17 (and_17[7], i0[7], i1[17]);
  and and_a7_b18 (and_18[7], i0[7], i1[18]);
  and and_a7_b19 (and_19[7], i0[7], i1[19]);
  and and_a7_b2 (and_2[7], i0[7], i1[2]);
  and and_a7_b20 (and_20[7], i0[7], i1[20]);
  and and_a7_b21 (and_21[7], i0[7], i1[21]);
  and and_a7_b22 (and_22[7], i0[7], i1[22]);
  and and_a7_b23 (and_23[7], i0[7], i1[23]);
  and and_a7_b24 (and_24[7], i0[7], i1[24]);
  and and_a7_b25 (and_25[7], i0[7], i1[25]);
  and and_a7_b26 (and_26[7], i0[7], i1[26]);
  and and_a7_b27 (and_27[7], i0[7], i1[27]);
  and and_a7_b28 (and_28[7], i0[7], i1[28]);
  and and_a7_b29 (and_29[7], i0[7], i1[29]);
  and and_a7_b3 (and_3[7], i0[7], i1[3]);
  and and_a7_b30 (and_30[7], i0[7], i1[30]);
  and and_a7_b31 (and_31[7], i0[7], i1[31]);
  and and_a7_b32 (nand_32[7], i0[7], i1[32]);
  and and_a7_b4 (and_4[7], i0[7], i1[4]);
  and and_a7_b5 (and_5[7], i0[7], i1[5]);
  and and_a7_b6 (and_6[7], i0[7], i1[6]);
  and and_a7_b7 (and_7[7], i0[7], i1[7]);
  and and_a7_b8 (and_8[7], i0[7], i1[8]);
  and and_a7_b9 (and_9[7], i0[7], i1[9]);
  and and_a8_b0 (and_0[8], i0[8], i1[0]);
  and and_a8_b1 (and_1[8], i0[8], i1[1]);
  and and_a8_b10 (and_10[8], i0[8], i1[10]);
  and and_a8_b11 (and_11[8], i0[8], i1[11]);
  and and_a8_b12 (and_12[8], i0[8], i1[12]);
  and and_a8_b13 (and_13[8], i0[8], i1[13]);
  and and_a8_b14 (and_14[8], i0[8], i1[14]);
  and and_a8_b15 (and_15[8], i0[8], i1[15]);
  and and_a8_b16 (and_16[8], i0[8], i1[16]);
  and and_a8_b17 (and_17[8], i0[8], i1[17]);
  and and_a8_b18 (and_18[8], i0[8], i1[18]);
  and and_a8_b19 (and_19[8], i0[8], i1[19]);
  and and_a8_b2 (and_2[8], i0[8], i1[2]);
  and and_a8_b20 (and_20[8], i0[8], i1[20]);
  and and_a8_b21 (and_21[8], i0[8], i1[21]);
  and and_a8_b22 (and_22[8], i0[8], i1[22]);
  and and_a8_b23 (and_23[8], i0[8], i1[23]);
  and and_a8_b24 (and_24[8], i0[8], i1[24]);
  and and_a8_b25 (and_25[8], i0[8], i1[25]);
  and and_a8_b26 (and_26[8], i0[8], i1[26]);
  and and_a8_b27 (and_27[8], i0[8], i1[27]);
  and and_a8_b28 (and_28[8], i0[8], i1[28]);
  and and_a8_b29 (and_29[8], i0[8], i1[29]);
  and and_a8_b3 (and_3[8], i0[8], i1[3]);
  and and_a8_b30 (and_30[8], i0[8], i1[30]);
  and and_a8_b31 (and_31[8], i0[8], i1[31]);
  and and_a8_b32 (nand_32[8], i0[8], i1[32]);
  and and_a8_b4 (and_4[8], i0[8], i1[4]);
  and and_a8_b5 (and_5[8], i0[8], i1[5]);
  and and_a8_b6 (and_6[8], i0[8], i1[6]);
  and and_a8_b7 (and_7[8], i0[8], i1[7]);
  and and_a8_b8 (and_8[8], i0[8], i1[8]);
  and and_a8_b9 (and_9[8], i0[8], i1[9]);
  and and_a9_b0 (and_0[9], i0[9], i1[0]);
  and and_a9_b1 (and_1[9], i0[9], i1[1]);
  and and_a9_b10 (and_10[9], i0[9], i1[10]);
  and and_a9_b11 (and_11[9], i0[9], i1[11]);
  and and_a9_b12 (and_12[9], i0[9], i1[12]);
  and and_a9_b13 (and_13[9], i0[9], i1[13]);
  and and_a9_b14 (and_14[9], i0[9], i1[14]);
  and and_a9_b15 (and_15[9], i0[9], i1[15]);
  and and_a9_b16 (and_16[9], i0[9], i1[16]);
  and and_a9_b17 (and_17[9], i0[9], i1[17]);
  and and_a9_b18 (and_18[9], i0[9], i1[18]);
  and and_a9_b19 (and_19[9], i0[9], i1[19]);
  and and_a9_b2 (and_2[9], i0[9], i1[2]);
  and and_a9_b20 (and_20[9], i0[9], i1[20]);
  and and_a9_b21 (and_21[9], i0[9], i1[21]);
  and and_a9_b22 (and_22[9], i0[9], i1[22]);
  and and_a9_b23 (and_23[9], i0[9], i1[23]);
  and and_a9_b24 (and_24[9], i0[9], i1[24]);
  and and_a9_b25 (and_25[9], i0[9], i1[25]);
  and and_a9_b26 (and_26[9], i0[9], i1[26]);
  and and_a9_b27 (and_27[9], i0[9], i1[27]);
  and and_a9_b28 (and_28[9], i0[9], i1[28]);
  and and_a9_b29 (and_29[9], i0[9], i1[29]);
  and and_a9_b3 (and_3[9], i0[9], i1[3]);
  and and_a9_b30 (and_30[9], i0[9], i1[30]);
  and and_a9_b31 (and_31[9], i0[9], i1[31]);
  and and_a9_b32 (nand_32[9], i0[9], i1[32]);
  and and_a9_b4 (and_4[9], i0[9], i1[4]);
  and and_a9_b5 (and_5[9], i0[9], i1[5]);
  and and_a9_b6 (and_6[9], i0[9], i1[6]);
  and and_a9_b7 (and_7[9], i0[9], i1[7]);
  and and_a9_b8 (and_8[9], i0[9], i1[8]);
  and and_a9_b9 (and_9[9], i0[9], i1[9]);
  add_pu64_pu61_pu60_pu59_pu58_pu57_pu56_pu55_pu54_pu53_pu52_pu51_pu50_pu49_pu48_pu47_pu46_pu45_pu44_pu43_pu42_pu41_pu40_pu39_pu38_pu37_pu36_pu35_pu34_pu33_pu32_mu63_mu63_o64 sum (
    .i0({and_32[31],1'b0,and_31[30],and_30[30],and_29[30],and_28[30],and_27[30],and_26[30],and_25[30],and_24[30],and_23[30],and_22[30],and_21[30],and_20[30],and_19[30],and_18[30],and_17[30],and_16[30],and_15[30],and_14[30],and_13[30],and_12[30],and_11[30],and_10[30],and_9[30],and_8[30],and_7[30],and_6[30],and_5[30],and_4[30],and_3[30],and_2[30],and_1[30],and_0[30:0]}),
    .i1({and_31[29],and_30[29],and_29[29],and_28[29],and_27[29],and_26[29],and_25[29],and_24[29],and_23[29],and_22[29],and_21[29],and_20[29],and_19[29],and_18[29],and_17[29],and_16[29],and_15[29],and_14[29],and_13[29],and_12[29],and_11[29],and_10[29],and_9[29],and_8[29],and_7[29],and_6[29],and_5[29],and_4[29],and_3[29],and_2[29],and_1[29:0],1'b0}),
    .i10({and_31[20],and_30[20],and_29[20],and_28[20],and_27[20],and_26[20],and_25[20],and_24[20],and_23[20],and_22[20],and_21[20],and_20[20],and_19[20],and_18[20],and_17[20],and_16[20],and_15[20],and_14[20],and_13[20],and_12[20],and_11[20],and_10[20:0],10'b0000000000}),
    .i11({and_31[19],and_30[19],and_29[19],and_28[19],and_27[19],and_26[19],and_25[19],and_24[19],and_23[19],and_22[19],and_21[19],and_20[19],and_19[19],and_18[19],and_17[19],and_16[19],and_15[19],and_14[19],and_13[19],and_12[19],and_11[19:0],11'b00000000000}),
    .i12({and_31[18],and_30[18],and_29[18],and_28[18],and_27[18],and_26[18],and_25[18],and_24[18],and_23[18],and_22[18],and_21[18],and_20[18],and_19[18],and_18[18],and_17[18],and_16[18],and_15[18],and_14[18],and_13[18],and_12[18:0],12'b000000000000}),
    .i13({and_31[17],and_30[17],and_29[17],and_28[17],and_27[17],and_26[17],and_25[17],and_24[17],and_23[17],and_22[17],and_21[17],and_20[17],and_19[17],and_18[17],and_17[17],and_16[17],and_15[17],and_14[17],and_13[17:0],13'b0000000000000}),
    .i14({and_31[16],and_30[16],and_29[16],and_28[16],and_27[16],and_26[16],and_25[16],and_24[16],and_23[16],and_22[16],and_21[16],and_20[16],and_19[16],and_18[16],and_17[16],and_16[16],and_15[16],and_14[16:0],14'b00000000000000}),
    .i15({and_31[15],and_30[15],and_29[15],and_28[15],and_27[15],and_26[15],and_25[15],and_24[15],and_23[15],and_22[15],and_21[15],and_20[15],and_19[15],and_18[15],and_17[15],and_16[15],and_15[15:0],15'b000000000000000}),
    .i16({and_31[14],and_30[14],and_29[14],and_28[14],and_27[14],and_26[14],and_25[14],and_24[14],and_23[14],and_22[14],and_21[14],and_20[14],and_19[14],and_18[14],and_17[14],and_16[14:0],16'b0000000000000000}),
    .i17({and_31[13],and_30[13],and_29[13],and_28[13],and_27[13],and_26[13],and_25[13],and_24[13],and_23[13],and_22[13],and_21[13],and_20[13],and_19[13],and_18[13],and_17[13:0],17'b00000000000000000}),
    .i18({and_31[12],and_30[12],and_29[12],and_28[12],and_27[12],and_26[12],and_25[12],and_24[12],and_23[12],and_22[12],and_21[12],and_20[12],and_19[12],and_18[12:0],18'b000000000000000000}),
    .i19({and_31[11],and_30[11],and_29[11],and_28[11],and_27[11],and_26[11],and_25[11],and_24[11],and_23[11],and_22[11],and_21[11],and_20[11],and_19[11:0],19'b0000000000000000000}),
    .i2({and_31[28],and_30[28],and_29[28],and_28[28],and_27[28],and_26[28],and_25[28],and_24[28],and_23[28],and_22[28],and_21[28],and_20[28],and_19[28],and_18[28],and_17[28],and_16[28],and_15[28],and_14[28],and_13[28],and_12[28],and_11[28],and_10[28],and_9[28],and_8[28],and_7[28],and_6[28],and_5[28],and_4[28],and_3[28],and_2[28:0],2'b00}),
    .i20({and_31[10],and_30[10],and_29[10],and_28[10],and_27[10],and_26[10],and_25[10],and_24[10],and_23[10],and_22[10],and_21[10],and_20[10:0],20'b00000000000000000000}),
    .i21({and_31[9],and_30[9],and_29[9],and_28[9],and_27[9],and_26[9],and_25[9],and_24[9],and_23[9],and_22[9],and_21[9:0],21'b000000000000000000000}),
    .i22({and_31[8],and_30[8],and_29[8],and_28[8],and_27[8],and_26[8],and_25[8],and_24[8],and_23[8],and_22[8:0],22'b0000000000000000000000}),
    .i23({and_31[7],and_30[7],and_29[7],and_28[7],and_27[7],and_26[7],and_25[7],and_24[7],and_23[7:0],23'b00000000000000000000000}),
    .i24({and_31[6],and_30[6],and_29[6],and_28[6],and_27[6],and_26[6],and_25[6],and_24[6:0],24'b000000000000000000000000}),
    .i25({and_31[5],and_30[5],and_29[5],and_28[5],and_27[5],and_26[5],and_25[5:0],25'b0000000000000000000000000}),
    .i26({and_31[4],and_30[4],and_29[4],and_28[4],and_27[4],and_26[4:0],26'b00000000000000000000000000}),
    .i27({and_31[3],and_30[3],and_29[3],and_28[3],and_27[3:0],27'b000000000000000000000000000}),
    .i28({and_31[2],and_30[2],and_29[2],and_28[2:0],28'b0000000000000000000000000000}),
    .i29({and_31[1],and_30[1],and_29[1:0],29'b00000000000000000000000000000}),
    .i3({and_31[27],and_30[27],and_29[27],and_28[27],and_27[27],and_26[27],and_25[27],and_24[27],and_23[27],and_22[27],and_21[27],and_20[27],and_19[27],and_18[27],and_17[27],and_16[27],and_15[27],and_14[27],and_13[27],and_12[27],and_11[27],and_10[27],and_9[27],and_8[27],and_7[27],and_6[27],and_5[27],and_4[27],and_3[27:0],3'b000}),
    .i30({and_31[0],and_30[0],30'b000000000000000000000000000000}),
    .i31({nand_31[31],nand_30[31],nand_29[31],nand_28[31],nand_27[31],nand_26[31],nand_25[31],nand_24[31],nand_23[31],nand_22[31],nand_21[31],nand_20[31],nand_19[31],nand_18[31],nand_17[31],nand_16[31],nand_15[31],nand_14[31],nand_13[31],nand_12[31],nand_11[31],nand_10[31],nand_9[31],nand_8[31],nand_7[31],nand_6[31],nand_5[31],nand_4[31],nand_3[31],nand_2[31],nand_1[31],nand_0[31],31'b0000000000000000000000000000000}),
    .i32({nand_32[30:0],32'b00000000000000000000000000000000}),
    .i4({and_31[26],and_30[26],and_29[26],and_28[26],and_27[26],and_26[26],and_25[26],and_24[26],and_23[26],and_22[26],and_21[26],and_20[26],and_19[26],and_18[26],and_17[26],and_16[26],and_15[26],and_14[26],and_13[26],and_12[26],and_11[26],and_10[26],and_9[26],and_8[26],and_7[26],and_6[26],and_5[26],and_4[26:0],4'b0000}),
    .i5({and_31[25],and_30[25],and_29[25],and_28[25],and_27[25],and_26[25],and_25[25],and_24[25],and_23[25],and_22[25],and_21[25],and_20[25],and_19[25],and_18[25],and_17[25],and_16[25],and_15[25],and_14[25],and_13[25],and_12[25],and_11[25],and_10[25],and_9[25],and_8[25],and_7[25],and_6[25],and_5[25:0],5'b00000}),
    .i6({and_31[24],and_30[24],and_29[24],and_28[24],and_27[24],and_26[24],and_25[24],and_24[24],and_23[24],and_22[24],and_21[24],and_20[24],and_19[24],and_18[24],and_17[24],and_16[24],and_15[24],and_14[24],and_13[24],and_12[24],and_11[24],and_10[24],and_9[24],and_8[24],and_7[24],and_6[24:0],6'b000000}),
    .i7({and_31[23],and_30[23],and_29[23],and_28[23],and_27[23],and_26[23],and_25[23],and_24[23],and_23[23],and_22[23],and_21[23],and_20[23],and_19[23],and_18[23],and_17[23],and_16[23],and_15[23],and_14[23],and_13[23],and_12[23],and_11[23],and_10[23],and_9[23],and_8[23],and_7[23:0],7'b0000000}),
    .i8({and_31[22],and_30[22],and_29[22],and_28[22],and_27[22],and_26[22],and_25[22],and_24[22],and_23[22],and_22[22],and_21[22],and_20[22],and_19[22],and_18[22],and_17[22],and_16[22],and_15[22],and_14[22],and_13[22],and_12[22],and_11[22],and_10[22],and_9[22],and_8[22:0],8'b00000000}),
    .i9({and_31[21],and_30[21],and_29[21],and_28[21],and_27[21],and_26[21],and_25[21],and_24[21],and_23[21],and_22[21],and_21[21],and_20[21],and_19[21],and_18[21],and_17[21],and_16[21],and_15[21],and_14[21],and_13[21],and_12[21],and_11[21],and_10[21],and_9[21:0],9'b000000000}),
    .o(o));

endmodule 

module add_mu32_o32
  (
  i0,
  o
  );

  input [31:0] i0;
  output [31:0] o;

  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b23;
  wire net_b24;
  wire net_b25;
  wire net_b26;
  wire net_b27;
  wire net_b28;
  wire net_b29;
  wire net_b3;
  wire net_b30;
  wire net_b31;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout23;
  wire net_cout24;
  wire net_cout25;
  wire net_cout26;
  wire net_cout27;
  wire net_cout28;
  wire net_cout29;
  wire net_cout3;
  wire net_cout30;
  wire net_cout31;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_nb0;
  wire net_nb1;
  wire net_nb10;
  wire net_nb11;
  wire net_nb12;
  wire net_nb13;
  wire net_nb14;
  wire net_nb15;
  wire net_nb16;
  wire net_nb17;
  wire net_nb18;
  wire net_nb19;
  wire net_nb2;
  wire net_nb20;
  wire net_nb21;
  wire net_nb22;
  wire net_nb23;
  wire net_nb24;
  wire net_nb25;
  wire net_nb26;
  wire net_nb27;
  wire net_nb28;
  wire net_nb29;
  wire net_nb3;
  wire net_nb30;
  wire net_nb31;
  wire net_nb4;
  wire net_nb5;
  wire net_nb6;
  wire net_nb7;
  wire net_nb8;
  wire net_nb9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum23;
  wire net_sum24;
  wire net_sum25;
  wire net_sum26;
  wire net_sum27;
  wire net_sum28;
  wire net_sum29;
  wire net_sum3;
  wire net_sum30;
  wire net_sum31;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_b31 = i0[31];
  assign net_b30 = i0[30];
  assign net_b29 = i0[29];
  assign net_b28 = i0[28];
  assign net_b27 = i0[27];
  assign net_b26 = i0[26];
  assign net_b25 = i0[25];
  assign net_b24 = i0[24];
  assign net_b23 = i0[23];
  assign net_b22 = i0[22];
  assign net_b21 = i0[21];
  assign net_b20 = i0[20];
  assign net_b19 = i0[19];
  assign net_b18 = i0[18];
  assign net_b17 = i0[17];
  assign net_b16 = i0[16];
  assign net_b15 = i0[15];
  assign net_b14 = i0[14];
  assign net_b13 = i0[13];
  assign net_b12 = i0[12];
  assign net_b11 = i0[11];
  assign net_b10 = i0[10];
  assign net_b9 = i0[9];
  assign net_b8 = i0[8];
  assign net_b7 = i0[7];
  assign net_b6 = i0[6];
  assign net_b5 = i0[5];
  assign net_b4 = i0[4];
  assign net_b3 = i0[3];
  assign net_b2 = i0[2];
  assign net_b1 = i0[1];
  assign net_b0 = i0[0];
  assign o[31] = net_sum31;
  assign o[30] = net_sum30;
  assign o[29] = net_sum29;
  assign o[28] = net_sum28;
  assign o[27] = net_sum27;
  assign o[26] = net_sum26;
  assign o[25] = net_sum25;
  assign o[24] = net_sum24;
  assign o[23] = net_sum23;
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(1'b0),
    .b(net_nb0),
    .c(1'b1),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(1'b0),
    .b(net_nb1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(1'b0),
    .b(net_nb10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(1'b0),
    .b(net_nb11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(1'b0),
    .b(net_nb12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(1'b0),
    .b(net_nb13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(1'b0),
    .b(net_nb14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(1'b0),
    .b(net_nb15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(1'b0),
    .b(net_nb16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(1'b0),
    .b(net_nb17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(1'b0),
    .b(net_nb18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(1'b0),
    .b(net_nb19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(1'b0),
    .b(net_nb2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(1'b0),
    .b(net_nb20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(1'b0),
    .b(net_nb21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(1'b0),
    .b(net_nb22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_23 (
    .a(1'b0),
    .b(net_nb23),
    .c(net_cout22),
    .cout(net_cout23),
    .sum(net_sum23));
  AL_FADD comp_24 (
    .a(1'b0),
    .b(net_nb24),
    .c(net_cout23),
    .cout(net_cout24),
    .sum(net_sum24));
  AL_FADD comp_25 (
    .a(1'b0),
    .b(net_nb25),
    .c(net_cout24),
    .cout(net_cout25),
    .sum(net_sum25));
  AL_FADD comp_26 (
    .a(1'b0),
    .b(net_nb26),
    .c(net_cout25),
    .cout(net_cout26),
    .sum(net_sum26));
  AL_FADD comp_27 (
    .a(1'b0),
    .b(net_nb27),
    .c(net_cout26),
    .cout(net_cout27),
    .sum(net_sum27));
  AL_FADD comp_28 (
    .a(1'b0),
    .b(net_nb28),
    .c(net_cout27),
    .cout(net_cout28),
    .sum(net_sum28));
  AL_FADD comp_29 (
    .a(1'b0),
    .b(net_nb29),
    .c(net_cout28),
    .cout(net_cout29),
    .sum(net_sum29));
  AL_FADD comp_3 (
    .a(1'b0),
    .b(net_nb3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_30 (
    .a(1'b0),
    .b(net_nb30),
    .c(net_cout29),
    .cout(net_cout30),
    .sum(net_sum30));
  AL_FADD comp_31 (
    .a(1'b0),
    .b(net_nb31),
    .c(net_cout30),
    .cout(net_cout31),
    .sum(net_sum31));
  AL_FADD comp_4 (
    .a(1'b0),
    .b(net_nb4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(1'b0),
    .b(net_nb5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(1'b0),
    .b(net_nb6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(1'b0),
    .b(net_nb7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(1'b0),
    .b(net_nb8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(1'b0),
    .b(net_nb9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));
  not inv_b0 (net_nb0, net_b0);
  not inv_b1 (net_nb1, net_b1);
  not inv_b10 (net_nb10, net_b10);
  not inv_b11 (net_nb11, net_b11);
  not inv_b12 (net_nb12, net_b12);
  not inv_b13 (net_nb13, net_b13);
  not inv_b14 (net_nb14, net_b14);
  not inv_b15 (net_nb15, net_b15);
  not inv_b16 (net_nb16, net_b16);
  not inv_b17 (net_nb17, net_b17);
  not inv_b18 (net_nb18, net_b18);
  not inv_b19 (net_nb19, net_b19);
  not inv_b2 (net_nb2, net_b2);
  not inv_b20 (net_nb20, net_b20);
  not inv_b21 (net_nb21, net_b21);
  not inv_b22 (net_nb22, net_b22);
  not inv_b23 (net_nb23, net_b23);
  not inv_b24 (net_nb24, net_b24);
  not inv_b25 (net_nb25, net_b25);
  not inv_b26 (net_nb26, net_b26);
  not inv_b27 (net_nb27, net_b27);
  not inv_b28 (net_nb28, net_b28);
  not inv_b29 (net_nb29, net_b29);
  not inv_b3 (net_nb3, net_b3);
  not inv_b30 (net_nb30, net_b30);
  not inv_b31 (net_nb31, net_b31);
  not inv_b4 (net_nb4, net_b4);
  not inv_b5 (net_nb5, net_b5);
  not inv_b6 (net_nb6, net_b6);
  not inv_b7 (net_nb7, net_b7);
  not inv_b8 (net_nb8, net_b8);
  not inv_b9 (net_nb9, net_b9);

endmodule 

module add_pu23_pu23_o23_1
  (
  i0,
  i1,
  o
  );

  input [22:0] i0;
  input [22:0] i1;
  output [22:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module eq_w24_1
  (
  i0,
  i1,
  o
  );

  input [23:0] i0;
  input [23:0] i1;
  output o;

  wire \or_or_or_or_xor_i0[0_o ;
  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_or_xor_i0[12]__o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[12]_i1[_o ;
  wire \or_or_xor_i0[18]_i1[_o ;
  wire \or_or_xor_i0[6]_i1[6_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[10]_i1[10]_o ;
  wire \or_xor_i0[12]_i1[12]_o ;
  wire \or_xor_i0[13]_i1[13]_o ;
  wire \or_xor_i0[15]_i1[15]_o ;
  wire \or_xor_i0[16]_i1[16]_o ;
  wire \or_xor_i0[18]_i1[18]_o ;
  wire \or_xor_i0[19]_i1[19]_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[21]_i1[21]_o ;
  wire \or_xor_i0[22]_i1[22]_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[7]_i1[7]_o_o ;
  wire \or_xor_i0[9]_i1[9]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[12]_i1[12]_o ;
  wire \xor_i0[13]_i1[13]_o ;
  wire \xor_i0[14]_i1[14]_o ;
  wire \xor_i0[15]_i1[15]_o ;
  wire \xor_i0[16]_i1[16]_o ;
  wire \xor_i0[17]_i1[17]_o ;
  wire \xor_i0[18]_i1[18]_o ;
  wire \xor_i0[19]_i1[19]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[20]_i1[20]_o ;
  wire \xor_i0[21]_i1[21]_o ;
  wire \xor_i0[22]_i1[22]_o ;
  wire \xor_i0[23]_i1[23]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, \or_or_or_or_xor_i0[0_o );
  or \or_or_or_or_xor_i0[0  (\or_or_or_or_xor_i0[0_o , \or_or_or_xor_i0[0]_i_o , \or_or_or_xor_i0[12]__o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[6]_i1[6_o );
  or \or_or_or_xor_i0[12]_  (\or_or_or_xor_i0[12]__o , \or_or_xor_i0[12]_i1[_o , \or_or_xor_i0[18]_i1[_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_or_xor_i0[12]_i1[  (\or_or_xor_i0[12]_i1[_o , \or_xor_i0[12]_i1[12]_o , \or_xor_i0[15]_i1[15]_o );
  or \or_or_xor_i0[18]_i1[  (\or_or_xor_i0[18]_i1[_o , \or_xor_i0[18]_i1[18]_o , \or_xor_i0[21]_i1[21]_o );
  or \or_or_xor_i0[6]_i1[6  (\or_or_xor_i0[6]_i1[6_o , \or_xor_i0[6]_i1[6]_o_o , \or_xor_i0[9]_i1[9]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[10]_i1[10]  (\or_xor_i0[10]_i1[10]_o , \xor_i0[10]_i1[10]_o , \xor_i0[11]_i1[11]_o );
  or \or_xor_i0[12]_i1[12]  (\or_xor_i0[12]_i1[12]_o , \xor_i0[12]_i1[12]_o , \or_xor_i0[13]_i1[13]_o );
  or \or_xor_i0[13]_i1[13]  (\or_xor_i0[13]_i1[13]_o , \xor_i0[13]_i1[13]_o , \xor_i0[14]_i1[14]_o );
  or \or_xor_i0[15]_i1[15]  (\or_xor_i0[15]_i1[15]_o , \xor_i0[15]_i1[15]_o , \or_xor_i0[16]_i1[16]_o );
  or \or_xor_i0[16]_i1[16]  (\or_xor_i0[16]_i1[16]_o , \xor_i0[16]_i1[16]_o , \xor_i0[17]_i1[17]_o );
  or \or_xor_i0[18]_i1[18]  (\or_xor_i0[18]_i1[18]_o , \xor_i0[18]_i1[18]_o , \or_xor_i0[19]_i1[19]_o );
  or \or_xor_i0[19]_i1[19]  (\or_xor_i0[19]_i1[19]_o , \xor_i0[19]_i1[19]_o , \xor_i0[20]_i1[20]_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[21]_i1[21]  (\or_xor_i0[21]_i1[21]_o , \xor_i0[21]_i1[21]_o , \or_xor_i0[22]_i1[22]_o );
  or \or_xor_i0[22]_i1[22]  (\or_xor_i0[22]_i1[22]_o , \xor_i0[22]_i1[22]_o , \xor_i0[23]_i1[23]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \or_xor_i0[4]_i1[4]_o_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \or_xor_i0[7]_i1[7]_o_o );
  or \or_xor_i0[7]_i1[7]_o  (\or_xor_i0[7]_i1[7]_o_o , \xor_i0[7]_i1[7]_o , \xor_i0[8]_i1[8]_o );
  or \or_xor_i0[9]_i1[9]_o  (\or_xor_i0[9]_i1[9]_o_o , \xor_i0[9]_i1[9]_o , \or_xor_i0[10]_i1[10]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (\xor_i0[12]_i1[12]_o , i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (\xor_i0[13]_i1[13]_o , i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (\xor_i0[14]_i1[14]_o , i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (\xor_i0[15]_i1[15]_o , i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (\xor_i0[16]_i1[16]_o , i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (\xor_i0[17]_i1[17]_o , i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (\xor_i0[18]_i1[18]_o , i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (\xor_i0[19]_i1[19]_o , i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (\xor_i0[20]_i1[20]_o , i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (\xor_i0[21]_i1[21]_o , i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (\xor_i0[22]_i1[22]_o , i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (\xor_i0[23]_i1[23]_o , i0[23], i1[23]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module add_pu47_pu46_pu45_pu44_pu43_pu42_pu41_pu40_pu39_pu38_pu37_pu36_pu35_pu34_pu33_pu32_pu31_pu30_pu29_pu28_pu27_pu26_pu25_pu24_o48
  (
  i0,
  i1,
  i10,
  i11,
  i12,
  i13,
  i14,
  i15,
  i16,
  i17,
  i18,
  i19,
  i2,
  i20,
  i21,
  i22,
  i23,
  i3,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  o
  );

  input [46:0] i0;
  input [45:0] i1;
  input [36:0] i10;
  input [35:0] i11;
  input [34:0] i12;
  input [33:0] i13;
  input [32:0] i14;
  input [31:0] i15;
  input [30:0] i16;
  input [29:0] i17;
  input [28:0] i18;
  input [27:0] i19;
  input [44:0] i2;
  input [26:0] i20;
  input [25:0] i21;
  input [24:0] i22;
  input [23:0] i23;
  input [43:0] i3;
  input [42:0] i4;
  input [41:0] i5;
  input [40:0] i6;
  input [39:0] i7;
  input [38:0] i8;
  input [37:0] i9;
  output [47:0] o;

  wire [46:0] cout_1;
  wire [47:0] cout_10;
  wire [47:0] cout_11;
  wire [47:0] cout_12;
  wire [47:0] cout_13;
  wire [47:0] cout_14;
  wire [47:0] cout_15;
  wire [47:0] cout_16;
  wire [47:0] cout_17;
  wire [47:0] cout_18;
  wire [47:0] cout_19;
  wire [47:0] cout_2;
  wire [47:0] cout_20;
  wire [47:0] cout_21;
  wire [47:0] cout_22;
  wire [47:0] cout_23;
  wire [47:0] cout_3;
  wire [47:0] cout_4;
  wire [47:0] cout_5;
  wire [47:0] cout_6;
  wire [47:0] cout_7;
  wire [47:0] cout_8;
  wire [47:0] cout_9;
  wire [46:0] sum_1;
  wire [47:0] sum_10;
  wire [47:0] sum_11;
  wire [47:0] sum_12;
  wire [47:0] sum_13;
  wire [47:0] sum_14;
  wire [47:0] sum_15;
  wire [47:0] sum_16;
  wire [47:0] sum_17;
  wire [47:0] sum_18;
  wire [47:0] sum_19;
  wire [47:0] sum_2;
  wire [47:0] sum_20;
  wire [47:0] sum_21;
  wire [47:0] sum_22;
  wire [47:0] sum_23;
  wire [47:0] sum_3;
  wire [47:0] sum_4;
  wire [47:0] sum_5;
  wire [47:0] sum_6;
  wire [47:0] sum_7;
  wire [47:0] sum_8;
  wire [47:0] sum_9;

  assign o[47] = sum_23[47];
  assign o[46] = sum_23[46];
  assign o[45] = sum_23[45];
  assign o[44] = sum_23[44];
  assign o[43] = sum_23[43];
  assign o[42] = sum_23[42];
  assign o[41] = sum_23[41];
  assign o[40] = sum_23[40];
  assign o[39] = sum_23[39];
  assign o[38] = sum_23[38];
  assign o[37] = sum_23[37];
  assign o[36] = sum_23[36];
  assign o[35] = sum_23[35];
  assign o[34] = sum_23[34];
  assign o[33] = sum_23[33];
  assign o[32] = sum_23[32];
  assign o[31] = sum_23[31];
  assign o[30] = sum_23[30];
  assign o[29] = sum_23[29];
  assign o[28] = sum_23[28];
  assign o[27] = sum_23[27];
  assign o[26] = sum_23[26];
  assign o[25] = sum_23[25];
  assign o[24] = sum_23[24];
  assign o[23] = sum_23[23];
  assign o[22] = sum_23[22];
  assign o[21] = sum_23[21];
  assign o[20] = sum_23[20];
  assign o[19] = sum_23[19];
  assign o[18] = sum_23[18];
  assign o[17] = sum_23[17];
  assign o[16] = sum_23[16];
  assign o[15] = sum_23[15];
  assign o[14] = sum_23[14];
  assign o[13] = sum_23[13];
  assign o[12] = sum_23[12];
  assign o[11] = sum_23[11];
  assign o[10] = sum_23[10];
  assign o[9] = sum_23[9];
  assign o[8] = sum_23[8];
  assign o[7] = sum_23[7];
  assign o[6] = sum_23[6];
  assign o[5] = sum_23[5];
  assign o[4] = sum_23[4];
  assign o[3] = sum_23[3];
  assign o[2] = sum_23[2];
  assign o[1] = sum_23[1];
  assign o[0] = sum_23[0];
  AL_FADD comp10_0 (
    .a(i10[0]),
    .b(sum_9[0]),
    .c(1'b0),
    .cout(cout_10[0]),
    .sum(sum_10[0]));
  AL_FADD comp10_1 (
    .a(i10[1]),
    .b(sum_9[1]),
    .c(cout_10[0]),
    .cout(cout_10[1]),
    .sum(sum_10[1]));
  AL_FADD comp10_10 (
    .a(i10[10]),
    .b(sum_9[10]),
    .c(cout_10[9]),
    .cout(cout_10[10]),
    .sum(sum_10[10]));
  AL_FADD comp10_11 (
    .a(i10[11]),
    .b(sum_9[11]),
    .c(cout_10[10]),
    .cout(cout_10[11]),
    .sum(sum_10[11]));
  AL_FADD comp10_12 (
    .a(i10[12]),
    .b(sum_9[12]),
    .c(cout_10[11]),
    .cout(cout_10[12]),
    .sum(sum_10[12]));
  AL_FADD comp10_13 (
    .a(i10[13]),
    .b(sum_9[13]),
    .c(cout_10[12]),
    .cout(cout_10[13]),
    .sum(sum_10[13]));
  AL_FADD comp10_14 (
    .a(i10[14]),
    .b(sum_9[14]),
    .c(cout_10[13]),
    .cout(cout_10[14]),
    .sum(sum_10[14]));
  AL_FADD comp10_15 (
    .a(i10[15]),
    .b(sum_9[15]),
    .c(cout_10[14]),
    .cout(cout_10[15]),
    .sum(sum_10[15]));
  AL_FADD comp10_16 (
    .a(i10[16]),
    .b(sum_9[16]),
    .c(cout_10[15]),
    .cout(cout_10[16]),
    .sum(sum_10[16]));
  AL_FADD comp10_17 (
    .a(i10[17]),
    .b(sum_9[17]),
    .c(cout_10[16]),
    .cout(cout_10[17]),
    .sum(sum_10[17]));
  AL_FADD comp10_18 (
    .a(i10[18]),
    .b(sum_9[18]),
    .c(cout_10[17]),
    .cout(cout_10[18]),
    .sum(sum_10[18]));
  AL_FADD comp10_19 (
    .a(i10[19]),
    .b(sum_9[19]),
    .c(cout_10[18]),
    .cout(cout_10[19]),
    .sum(sum_10[19]));
  AL_FADD comp10_2 (
    .a(i10[2]),
    .b(sum_9[2]),
    .c(cout_10[1]),
    .cout(cout_10[2]),
    .sum(sum_10[2]));
  AL_FADD comp10_20 (
    .a(i10[20]),
    .b(sum_9[20]),
    .c(cout_10[19]),
    .cout(cout_10[20]),
    .sum(sum_10[20]));
  AL_FADD comp10_21 (
    .a(i10[21]),
    .b(sum_9[21]),
    .c(cout_10[20]),
    .cout(cout_10[21]),
    .sum(sum_10[21]));
  AL_FADD comp10_22 (
    .a(i10[22]),
    .b(sum_9[22]),
    .c(cout_10[21]),
    .cout(cout_10[22]),
    .sum(sum_10[22]));
  AL_FADD comp10_23 (
    .a(i10[23]),
    .b(sum_9[23]),
    .c(cout_10[22]),
    .cout(cout_10[23]),
    .sum(sum_10[23]));
  AL_FADD comp10_24 (
    .a(i10[24]),
    .b(sum_9[24]),
    .c(cout_10[23]),
    .cout(cout_10[24]),
    .sum(sum_10[24]));
  AL_FADD comp10_25 (
    .a(i10[25]),
    .b(sum_9[25]),
    .c(cout_10[24]),
    .cout(cout_10[25]),
    .sum(sum_10[25]));
  AL_FADD comp10_26 (
    .a(i10[26]),
    .b(sum_9[26]),
    .c(cout_10[25]),
    .cout(cout_10[26]),
    .sum(sum_10[26]));
  AL_FADD comp10_27 (
    .a(i10[27]),
    .b(sum_9[27]),
    .c(cout_10[26]),
    .cout(cout_10[27]),
    .sum(sum_10[27]));
  AL_FADD comp10_28 (
    .a(i10[28]),
    .b(sum_9[28]),
    .c(cout_10[27]),
    .cout(cout_10[28]),
    .sum(sum_10[28]));
  AL_FADD comp10_29 (
    .a(i10[29]),
    .b(sum_9[29]),
    .c(cout_10[28]),
    .cout(cout_10[29]),
    .sum(sum_10[29]));
  AL_FADD comp10_3 (
    .a(i10[3]),
    .b(sum_9[3]),
    .c(cout_10[2]),
    .cout(cout_10[3]),
    .sum(sum_10[3]));
  AL_FADD comp10_30 (
    .a(i10[30]),
    .b(sum_9[30]),
    .c(cout_10[29]),
    .cout(cout_10[30]),
    .sum(sum_10[30]));
  AL_FADD comp10_31 (
    .a(i10[31]),
    .b(sum_9[31]),
    .c(cout_10[30]),
    .cout(cout_10[31]),
    .sum(sum_10[31]));
  AL_FADD comp10_32 (
    .a(i10[32]),
    .b(sum_9[32]),
    .c(cout_10[31]),
    .cout(cout_10[32]),
    .sum(sum_10[32]));
  AL_FADD comp10_33 (
    .a(i10[33]),
    .b(sum_9[33]),
    .c(cout_10[32]),
    .cout(cout_10[33]),
    .sum(sum_10[33]));
  AL_FADD comp10_34 (
    .a(i10[34]),
    .b(sum_9[34]),
    .c(cout_10[33]),
    .cout(cout_10[34]),
    .sum(sum_10[34]));
  AL_FADD comp10_35 (
    .a(i10[35]),
    .b(sum_9[35]),
    .c(cout_10[34]),
    .cout(cout_10[35]),
    .sum(sum_10[35]));
  AL_FADD comp10_36 (
    .a(i10[36]),
    .b(sum_9[36]),
    .c(cout_10[35]),
    .cout(cout_10[36]),
    .sum(sum_10[36]));
  AL_FADD comp10_37 (
    .a(1'b0),
    .b(sum_9[37]),
    .c(cout_10[36]),
    .cout(cout_10[37]),
    .sum(sum_10[37]));
  AL_FADD comp10_38 (
    .a(1'b0),
    .b(sum_9[38]),
    .c(cout_10[37]),
    .cout(cout_10[38]),
    .sum(sum_10[38]));
  AL_FADD comp10_39 (
    .a(1'b0),
    .b(sum_9[39]),
    .c(cout_10[38]),
    .cout(cout_10[39]),
    .sum(sum_10[39]));
  AL_FADD comp10_4 (
    .a(i10[4]),
    .b(sum_9[4]),
    .c(cout_10[3]),
    .cout(cout_10[4]),
    .sum(sum_10[4]));
  AL_FADD comp10_40 (
    .a(1'b0),
    .b(sum_9[40]),
    .c(cout_10[39]),
    .cout(cout_10[40]),
    .sum(sum_10[40]));
  AL_FADD comp10_41 (
    .a(1'b0),
    .b(sum_9[41]),
    .c(cout_10[40]),
    .cout(cout_10[41]),
    .sum(sum_10[41]));
  AL_FADD comp10_42 (
    .a(1'b0),
    .b(sum_9[42]),
    .c(cout_10[41]),
    .cout(cout_10[42]),
    .sum(sum_10[42]));
  AL_FADD comp10_43 (
    .a(1'b0),
    .b(sum_9[43]),
    .c(cout_10[42]),
    .cout(cout_10[43]),
    .sum(sum_10[43]));
  AL_FADD comp10_44 (
    .a(1'b0),
    .b(sum_9[44]),
    .c(cout_10[43]),
    .cout(cout_10[44]),
    .sum(sum_10[44]));
  AL_FADD comp10_45 (
    .a(1'b0),
    .b(sum_9[45]),
    .c(cout_10[44]),
    .cout(cout_10[45]),
    .sum(sum_10[45]));
  AL_FADD comp10_46 (
    .a(1'b0),
    .b(sum_9[46]),
    .c(cout_10[45]),
    .cout(cout_10[46]),
    .sum(sum_10[46]));
  AL_FADD comp10_47 (
    .a(1'b0),
    .b(sum_9[47]),
    .c(cout_10[46]),
    .cout(cout_10[47]),
    .sum(sum_10[47]));
  AL_FADD comp10_5 (
    .a(i10[5]),
    .b(sum_9[5]),
    .c(cout_10[4]),
    .cout(cout_10[5]),
    .sum(sum_10[5]));
  AL_FADD comp10_6 (
    .a(i10[6]),
    .b(sum_9[6]),
    .c(cout_10[5]),
    .cout(cout_10[6]),
    .sum(sum_10[6]));
  AL_FADD comp10_7 (
    .a(i10[7]),
    .b(sum_9[7]),
    .c(cout_10[6]),
    .cout(cout_10[7]),
    .sum(sum_10[7]));
  AL_FADD comp10_8 (
    .a(i10[8]),
    .b(sum_9[8]),
    .c(cout_10[7]),
    .cout(cout_10[8]),
    .sum(sum_10[8]));
  AL_FADD comp10_9 (
    .a(i10[9]),
    .b(sum_9[9]),
    .c(cout_10[8]),
    .cout(cout_10[9]),
    .sum(sum_10[9]));
  AL_FADD comp11_0 (
    .a(i11[0]),
    .b(sum_10[0]),
    .c(1'b0),
    .cout(cout_11[0]),
    .sum(sum_11[0]));
  AL_FADD comp11_1 (
    .a(i11[1]),
    .b(sum_10[1]),
    .c(cout_11[0]),
    .cout(cout_11[1]),
    .sum(sum_11[1]));
  AL_FADD comp11_10 (
    .a(i11[10]),
    .b(sum_10[10]),
    .c(cout_11[9]),
    .cout(cout_11[10]),
    .sum(sum_11[10]));
  AL_FADD comp11_11 (
    .a(i11[11]),
    .b(sum_10[11]),
    .c(cout_11[10]),
    .cout(cout_11[11]),
    .sum(sum_11[11]));
  AL_FADD comp11_12 (
    .a(i11[12]),
    .b(sum_10[12]),
    .c(cout_11[11]),
    .cout(cout_11[12]),
    .sum(sum_11[12]));
  AL_FADD comp11_13 (
    .a(i11[13]),
    .b(sum_10[13]),
    .c(cout_11[12]),
    .cout(cout_11[13]),
    .sum(sum_11[13]));
  AL_FADD comp11_14 (
    .a(i11[14]),
    .b(sum_10[14]),
    .c(cout_11[13]),
    .cout(cout_11[14]),
    .sum(sum_11[14]));
  AL_FADD comp11_15 (
    .a(i11[15]),
    .b(sum_10[15]),
    .c(cout_11[14]),
    .cout(cout_11[15]),
    .sum(sum_11[15]));
  AL_FADD comp11_16 (
    .a(i11[16]),
    .b(sum_10[16]),
    .c(cout_11[15]),
    .cout(cout_11[16]),
    .sum(sum_11[16]));
  AL_FADD comp11_17 (
    .a(i11[17]),
    .b(sum_10[17]),
    .c(cout_11[16]),
    .cout(cout_11[17]),
    .sum(sum_11[17]));
  AL_FADD comp11_18 (
    .a(i11[18]),
    .b(sum_10[18]),
    .c(cout_11[17]),
    .cout(cout_11[18]),
    .sum(sum_11[18]));
  AL_FADD comp11_19 (
    .a(i11[19]),
    .b(sum_10[19]),
    .c(cout_11[18]),
    .cout(cout_11[19]),
    .sum(sum_11[19]));
  AL_FADD comp11_2 (
    .a(i11[2]),
    .b(sum_10[2]),
    .c(cout_11[1]),
    .cout(cout_11[2]),
    .sum(sum_11[2]));
  AL_FADD comp11_20 (
    .a(i11[20]),
    .b(sum_10[20]),
    .c(cout_11[19]),
    .cout(cout_11[20]),
    .sum(sum_11[20]));
  AL_FADD comp11_21 (
    .a(i11[21]),
    .b(sum_10[21]),
    .c(cout_11[20]),
    .cout(cout_11[21]),
    .sum(sum_11[21]));
  AL_FADD comp11_22 (
    .a(i11[22]),
    .b(sum_10[22]),
    .c(cout_11[21]),
    .cout(cout_11[22]),
    .sum(sum_11[22]));
  AL_FADD comp11_23 (
    .a(i11[23]),
    .b(sum_10[23]),
    .c(cout_11[22]),
    .cout(cout_11[23]),
    .sum(sum_11[23]));
  AL_FADD comp11_24 (
    .a(i11[24]),
    .b(sum_10[24]),
    .c(cout_11[23]),
    .cout(cout_11[24]),
    .sum(sum_11[24]));
  AL_FADD comp11_25 (
    .a(i11[25]),
    .b(sum_10[25]),
    .c(cout_11[24]),
    .cout(cout_11[25]),
    .sum(sum_11[25]));
  AL_FADD comp11_26 (
    .a(i11[26]),
    .b(sum_10[26]),
    .c(cout_11[25]),
    .cout(cout_11[26]),
    .sum(sum_11[26]));
  AL_FADD comp11_27 (
    .a(i11[27]),
    .b(sum_10[27]),
    .c(cout_11[26]),
    .cout(cout_11[27]),
    .sum(sum_11[27]));
  AL_FADD comp11_28 (
    .a(i11[28]),
    .b(sum_10[28]),
    .c(cout_11[27]),
    .cout(cout_11[28]),
    .sum(sum_11[28]));
  AL_FADD comp11_29 (
    .a(i11[29]),
    .b(sum_10[29]),
    .c(cout_11[28]),
    .cout(cout_11[29]),
    .sum(sum_11[29]));
  AL_FADD comp11_3 (
    .a(i11[3]),
    .b(sum_10[3]),
    .c(cout_11[2]),
    .cout(cout_11[3]),
    .sum(sum_11[3]));
  AL_FADD comp11_30 (
    .a(i11[30]),
    .b(sum_10[30]),
    .c(cout_11[29]),
    .cout(cout_11[30]),
    .sum(sum_11[30]));
  AL_FADD comp11_31 (
    .a(i11[31]),
    .b(sum_10[31]),
    .c(cout_11[30]),
    .cout(cout_11[31]),
    .sum(sum_11[31]));
  AL_FADD comp11_32 (
    .a(i11[32]),
    .b(sum_10[32]),
    .c(cout_11[31]),
    .cout(cout_11[32]),
    .sum(sum_11[32]));
  AL_FADD comp11_33 (
    .a(i11[33]),
    .b(sum_10[33]),
    .c(cout_11[32]),
    .cout(cout_11[33]),
    .sum(sum_11[33]));
  AL_FADD comp11_34 (
    .a(i11[34]),
    .b(sum_10[34]),
    .c(cout_11[33]),
    .cout(cout_11[34]),
    .sum(sum_11[34]));
  AL_FADD comp11_35 (
    .a(i11[35]),
    .b(sum_10[35]),
    .c(cout_11[34]),
    .cout(cout_11[35]),
    .sum(sum_11[35]));
  AL_FADD comp11_36 (
    .a(1'b0),
    .b(sum_10[36]),
    .c(cout_11[35]),
    .cout(cout_11[36]),
    .sum(sum_11[36]));
  AL_FADD comp11_37 (
    .a(1'b0),
    .b(sum_10[37]),
    .c(cout_11[36]),
    .cout(cout_11[37]),
    .sum(sum_11[37]));
  AL_FADD comp11_38 (
    .a(1'b0),
    .b(sum_10[38]),
    .c(cout_11[37]),
    .cout(cout_11[38]),
    .sum(sum_11[38]));
  AL_FADD comp11_39 (
    .a(1'b0),
    .b(sum_10[39]),
    .c(cout_11[38]),
    .cout(cout_11[39]),
    .sum(sum_11[39]));
  AL_FADD comp11_4 (
    .a(i11[4]),
    .b(sum_10[4]),
    .c(cout_11[3]),
    .cout(cout_11[4]),
    .sum(sum_11[4]));
  AL_FADD comp11_40 (
    .a(1'b0),
    .b(sum_10[40]),
    .c(cout_11[39]),
    .cout(cout_11[40]),
    .sum(sum_11[40]));
  AL_FADD comp11_41 (
    .a(1'b0),
    .b(sum_10[41]),
    .c(cout_11[40]),
    .cout(cout_11[41]),
    .sum(sum_11[41]));
  AL_FADD comp11_42 (
    .a(1'b0),
    .b(sum_10[42]),
    .c(cout_11[41]),
    .cout(cout_11[42]),
    .sum(sum_11[42]));
  AL_FADD comp11_43 (
    .a(1'b0),
    .b(sum_10[43]),
    .c(cout_11[42]),
    .cout(cout_11[43]),
    .sum(sum_11[43]));
  AL_FADD comp11_44 (
    .a(1'b0),
    .b(sum_10[44]),
    .c(cout_11[43]),
    .cout(cout_11[44]),
    .sum(sum_11[44]));
  AL_FADD comp11_45 (
    .a(1'b0),
    .b(sum_10[45]),
    .c(cout_11[44]),
    .cout(cout_11[45]),
    .sum(sum_11[45]));
  AL_FADD comp11_46 (
    .a(1'b0),
    .b(sum_10[46]),
    .c(cout_11[45]),
    .cout(cout_11[46]),
    .sum(sum_11[46]));
  AL_FADD comp11_47 (
    .a(1'b0),
    .b(sum_10[47]),
    .c(cout_11[46]),
    .cout(cout_11[47]),
    .sum(sum_11[47]));
  AL_FADD comp11_5 (
    .a(i11[5]),
    .b(sum_10[5]),
    .c(cout_11[4]),
    .cout(cout_11[5]),
    .sum(sum_11[5]));
  AL_FADD comp11_6 (
    .a(i11[6]),
    .b(sum_10[6]),
    .c(cout_11[5]),
    .cout(cout_11[6]),
    .sum(sum_11[6]));
  AL_FADD comp11_7 (
    .a(i11[7]),
    .b(sum_10[7]),
    .c(cout_11[6]),
    .cout(cout_11[7]),
    .sum(sum_11[7]));
  AL_FADD comp11_8 (
    .a(i11[8]),
    .b(sum_10[8]),
    .c(cout_11[7]),
    .cout(cout_11[8]),
    .sum(sum_11[8]));
  AL_FADD comp11_9 (
    .a(i11[9]),
    .b(sum_10[9]),
    .c(cout_11[8]),
    .cout(cout_11[9]),
    .sum(sum_11[9]));
  AL_FADD comp12_0 (
    .a(i12[0]),
    .b(sum_11[0]),
    .c(1'b0),
    .cout(cout_12[0]),
    .sum(sum_12[0]));
  AL_FADD comp12_1 (
    .a(i12[1]),
    .b(sum_11[1]),
    .c(cout_12[0]),
    .cout(cout_12[1]),
    .sum(sum_12[1]));
  AL_FADD comp12_10 (
    .a(i12[10]),
    .b(sum_11[10]),
    .c(cout_12[9]),
    .cout(cout_12[10]),
    .sum(sum_12[10]));
  AL_FADD comp12_11 (
    .a(i12[11]),
    .b(sum_11[11]),
    .c(cout_12[10]),
    .cout(cout_12[11]),
    .sum(sum_12[11]));
  AL_FADD comp12_12 (
    .a(i12[12]),
    .b(sum_11[12]),
    .c(cout_12[11]),
    .cout(cout_12[12]),
    .sum(sum_12[12]));
  AL_FADD comp12_13 (
    .a(i12[13]),
    .b(sum_11[13]),
    .c(cout_12[12]),
    .cout(cout_12[13]),
    .sum(sum_12[13]));
  AL_FADD comp12_14 (
    .a(i12[14]),
    .b(sum_11[14]),
    .c(cout_12[13]),
    .cout(cout_12[14]),
    .sum(sum_12[14]));
  AL_FADD comp12_15 (
    .a(i12[15]),
    .b(sum_11[15]),
    .c(cout_12[14]),
    .cout(cout_12[15]),
    .sum(sum_12[15]));
  AL_FADD comp12_16 (
    .a(i12[16]),
    .b(sum_11[16]),
    .c(cout_12[15]),
    .cout(cout_12[16]),
    .sum(sum_12[16]));
  AL_FADD comp12_17 (
    .a(i12[17]),
    .b(sum_11[17]),
    .c(cout_12[16]),
    .cout(cout_12[17]),
    .sum(sum_12[17]));
  AL_FADD comp12_18 (
    .a(i12[18]),
    .b(sum_11[18]),
    .c(cout_12[17]),
    .cout(cout_12[18]),
    .sum(sum_12[18]));
  AL_FADD comp12_19 (
    .a(i12[19]),
    .b(sum_11[19]),
    .c(cout_12[18]),
    .cout(cout_12[19]),
    .sum(sum_12[19]));
  AL_FADD comp12_2 (
    .a(i12[2]),
    .b(sum_11[2]),
    .c(cout_12[1]),
    .cout(cout_12[2]),
    .sum(sum_12[2]));
  AL_FADD comp12_20 (
    .a(i12[20]),
    .b(sum_11[20]),
    .c(cout_12[19]),
    .cout(cout_12[20]),
    .sum(sum_12[20]));
  AL_FADD comp12_21 (
    .a(i12[21]),
    .b(sum_11[21]),
    .c(cout_12[20]),
    .cout(cout_12[21]),
    .sum(sum_12[21]));
  AL_FADD comp12_22 (
    .a(i12[22]),
    .b(sum_11[22]),
    .c(cout_12[21]),
    .cout(cout_12[22]),
    .sum(sum_12[22]));
  AL_FADD comp12_23 (
    .a(i12[23]),
    .b(sum_11[23]),
    .c(cout_12[22]),
    .cout(cout_12[23]),
    .sum(sum_12[23]));
  AL_FADD comp12_24 (
    .a(i12[24]),
    .b(sum_11[24]),
    .c(cout_12[23]),
    .cout(cout_12[24]),
    .sum(sum_12[24]));
  AL_FADD comp12_25 (
    .a(i12[25]),
    .b(sum_11[25]),
    .c(cout_12[24]),
    .cout(cout_12[25]),
    .sum(sum_12[25]));
  AL_FADD comp12_26 (
    .a(i12[26]),
    .b(sum_11[26]),
    .c(cout_12[25]),
    .cout(cout_12[26]),
    .sum(sum_12[26]));
  AL_FADD comp12_27 (
    .a(i12[27]),
    .b(sum_11[27]),
    .c(cout_12[26]),
    .cout(cout_12[27]),
    .sum(sum_12[27]));
  AL_FADD comp12_28 (
    .a(i12[28]),
    .b(sum_11[28]),
    .c(cout_12[27]),
    .cout(cout_12[28]),
    .sum(sum_12[28]));
  AL_FADD comp12_29 (
    .a(i12[29]),
    .b(sum_11[29]),
    .c(cout_12[28]),
    .cout(cout_12[29]),
    .sum(sum_12[29]));
  AL_FADD comp12_3 (
    .a(i12[3]),
    .b(sum_11[3]),
    .c(cout_12[2]),
    .cout(cout_12[3]),
    .sum(sum_12[3]));
  AL_FADD comp12_30 (
    .a(i12[30]),
    .b(sum_11[30]),
    .c(cout_12[29]),
    .cout(cout_12[30]),
    .sum(sum_12[30]));
  AL_FADD comp12_31 (
    .a(i12[31]),
    .b(sum_11[31]),
    .c(cout_12[30]),
    .cout(cout_12[31]),
    .sum(sum_12[31]));
  AL_FADD comp12_32 (
    .a(i12[32]),
    .b(sum_11[32]),
    .c(cout_12[31]),
    .cout(cout_12[32]),
    .sum(sum_12[32]));
  AL_FADD comp12_33 (
    .a(i12[33]),
    .b(sum_11[33]),
    .c(cout_12[32]),
    .cout(cout_12[33]),
    .sum(sum_12[33]));
  AL_FADD comp12_34 (
    .a(i12[34]),
    .b(sum_11[34]),
    .c(cout_12[33]),
    .cout(cout_12[34]),
    .sum(sum_12[34]));
  AL_FADD comp12_35 (
    .a(1'b0),
    .b(sum_11[35]),
    .c(cout_12[34]),
    .cout(cout_12[35]),
    .sum(sum_12[35]));
  AL_FADD comp12_36 (
    .a(1'b0),
    .b(sum_11[36]),
    .c(cout_12[35]),
    .cout(cout_12[36]),
    .sum(sum_12[36]));
  AL_FADD comp12_37 (
    .a(1'b0),
    .b(sum_11[37]),
    .c(cout_12[36]),
    .cout(cout_12[37]),
    .sum(sum_12[37]));
  AL_FADD comp12_38 (
    .a(1'b0),
    .b(sum_11[38]),
    .c(cout_12[37]),
    .cout(cout_12[38]),
    .sum(sum_12[38]));
  AL_FADD comp12_39 (
    .a(1'b0),
    .b(sum_11[39]),
    .c(cout_12[38]),
    .cout(cout_12[39]),
    .sum(sum_12[39]));
  AL_FADD comp12_4 (
    .a(i12[4]),
    .b(sum_11[4]),
    .c(cout_12[3]),
    .cout(cout_12[4]),
    .sum(sum_12[4]));
  AL_FADD comp12_40 (
    .a(1'b0),
    .b(sum_11[40]),
    .c(cout_12[39]),
    .cout(cout_12[40]),
    .sum(sum_12[40]));
  AL_FADD comp12_41 (
    .a(1'b0),
    .b(sum_11[41]),
    .c(cout_12[40]),
    .cout(cout_12[41]),
    .sum(sum_12[41]));
  AL_FADD comp12_42 (
    .a(1'b0),
    .b(sum_11[42]),
    .c(cout_12[41]),
    .cout(cout_12[42]),
    .sum(sum_12[42]));
  AL_FADD comp12_43 (
    .a(1'b0),
    .b(sum_11[43]),
    .c(cout_12[42]),
    .cout(cout_12[43]),
    .sum(sum_12[43]));
  AL_FADD comp12_44 (
    .a(1'b0),
    .b(sum_11[44]),
    .c(cout_12[43]),
    .cout(cout_12[44]),
    .sum(sum_12[44]));
  AL_FADD comp12_45 (
    .a(1'b0),
    .b(sum_11[45]),
    .c(cout_12[44]),
    .cout(cout_12[45]),
    .sum(sum_12[45]));
  AL_FADD comp12_46 (
    .a(1'b0),
    .b(sum_11[46]),
    .c(cout_12[45]),
    .cout(cout_12[46]),
    .sum(sum_12[46]));
  AL_FADD comp12_47 (
    .a(1'b0),
    .b(sum_11[47]),
    .c(cout_12[46]),
    .cout(cout_12[47]),
    .sum(sum_12[47]));
  AL_FADD comp12_5 (
    .a(i12[5]),
    .b(sum_11[5]),
    .c(cout_12[4]),
    .cout(cout_12[5]),
    .sum(sum_12[5]));
  AL_FADD comp12_6 (
    .a(i12[6]),
    .b(sum_11[6]),
    .c(cout_12[5]),
    .cout(cout_12[6]),
    .sum(sum_12[6]));
  AL_FADD comp12_7 (
    .a(i12[7]),
    .b(sum_11[7]),
    .c(cout_12[6]),
    .cout(cout_12[7]),
    .sum(sum_12[7]));
  AL_FADD comp12_8 (
    .a(i12[8]),
    .b(sum_11[8]),
    .c(cout_12[7]),
    .cout(cout_12[8]),
    .sum(sum_12[8]));
  AL_FADD comp12_9 (
    .a(i12[9]),
    .b(sum_11[9]),
    .c(cout_12[8]),
    .cout(cout_12[9]),
    .sum(sum_12[9]));
  AL_FADD comp13_0 (
    .a(i13[0]),
    .b(sum_12[0]),
    .c(1'b0),
    .cout(cout_13[0]),
    .sum(sum_13[0]));
  AL_FADD comp13_1 (
    .a(i13[1]),
    .b(sum_12[1]),
    .c(cout_13[0]),
    .cout(cout_13[1]),
    .sum(sum_13[1]));
  AL_FADD comp13_10 (
    .a(i13[10]),
    .b(sum_12[10]),
    .c(cout_13[9]),
    .cout(cout_13[10]),
    .sum(sum_13[10]));
  AL_FADD comp13_11 (
    .a(i13[11]),
    .b(sum_12[11]),
    .c(cout_13[10]),
    .cout(cout_13[11]),
    .sum(sum_13[11]));
  AL_FADD comp13_12 (
    .a(i13[12]),
    .b(sum_12[12]),
    .c(cout_13[11]),
    .cout(cout_13[12]),
    .sum(sum_13[12]));
  AL_FADD comp13_13 (
    .a(i13[13]),
    .b(sum_12[13]),
    .c(cout_13[12]),
    .cout(cout_13[13]),
    .sum(sum_13[13]));
  AL_FADD comp13_14 (
    .a(i13[14]),
    .b(sum_12[14]),
    .c(cout_13[13]),
    .cout(cout_13[14]),
    .sum(sum_13[14]));
  AL_FADD comp13_15 (
    .a(i13[15]),
    .b(sum_12[15]),
    .c(cout_13[14]),
    .cout(cout_13[15]),
    .sum(sum_13[15]));
  AL_FADD comp13_16 (
    .a(i13[16]),
    .b(sum_12[16]),
    .c(cout_13[15]),
    .cout(cout_13[16]),
    .sum(sum_13[16]));
  AL_FADD comp13_17 (
    .a(i13[17]),
    .b(sum_12[17]),
    .c(cout_13[16]),
    .cout(cout_13[17]),
    .sum(sum_13[17]));
  AL_FADD comp13_18 (
    .a(i13[18]),
    .b(sum_12[18]),
    .c(cout_13[17]),
    .cout(cout_13[18]),
    .sum(sum_13[18]));
  AL_FADD comp13_19 (
    .a(i13[19]),
    .b(sum_12[19]),
    .c(cout_13[18]),
    .cout(cout_13[19]),
    .sum(sum_13[19]));
  AL_FADD comp13_2 (
    .a(i13[2]),
    .b(sum_12[2]),
    .c(cout_13[1]),
    .cout(cout_13[2]),
    .sum(sum_13[2]));
  AL_FADD comp13_20 (
    .a(i13[20]),
    .b(sum_12[20]),
    .c(cout_13[19]),
    .cout(cout_13[20]),
    .sum(sum_13[20]));
  AL_FADD comp13_21 (
    .a(i13[21]),
    .b(sum_12[21]),
    .c(cout_13[20]),
    .cout(cout_13[21]),
    .sum(sum_13[21]));
  AL_FADD comp13_22 (
    .a(i13[22]),
    .b(sum_12[22]),
    .c(cout_13[21]),
    .cout(cout_13[22]),
    .sum(sum_13[22]));
  AL_FADD comp13_23 (
    .a(i13[23]),
    .b(sum_12[23]),
    .c(cout_13[22]),
    .cout(cout_13[23]),
    .sum(sum_13[23]));
  AL_FADD comp13_24 (
    .a(i13[24]),
    .b(sum_12[24]),
    .c(cout_13[23]),
    .cout(cout_13[24]),
    .sum(sum_13[24]));
  AL_FADD comp13_25 (
    .a(i13[25]),
    .b(sum_12[25]),
    .c(cout_13[24]),
    .cout(cout_13[25]),
    .sum(sum_13[25]));
  AL_FADD comp13_26 (
    .a(i13[26]),
    .b(sum_12[26]),
    .c(cout_13[25]),
    .cout(cout_13[26]),
    .sum(sum_13[26]));
  AL_FADD comp13_27 (
    .a(i13[27]),
    .b(sum_12[27]),
    .c(cout_13[26]),
    .cout(cout_13[27]),
    .sum(sum_13[27]));
  AL_FADD comp13_28 (
    .a(i13[28]),
    .b(sum_12[28]),
    .c(cout_13[27]),
    .cout(cout_13[28]),
    .sum(sum_13[28]));
  AL_FADD comp13_29 (
    .a(i13[29]),
    .b(sum_12[29]),
    .c(cout_13[28]),
    .cout(cout_13[29]),
    .sum(sum_13[29]));
  AL_FADD comp13_3 (
    .a(i13[3]),
    .b(sum_12[3]),
    .c(cout_13[2]),
    .cout(cout_13[3]),
    .sum(sum_13[3]));
  AL_FADD comp13_30 (
    .a(i13[30]),
    .b(sum_12[30]),
    .c(cout_13[29]),
    .cout(cout_13[30]),
    .sum(sum_13[30]));
  AL_FADD comp13_31 (
    .a(i13[31]),
    .b(sum_12[31]),
    .c(cout_13[30]),
    .cout(cout_13[31]),
    .sum(sum_13[31]));
  AL_FADD comp13_32 (
    .a(i13[32]),
    .b(sum_12[32]),
    .c(cout_13[31]),
    .cout(cout_13[32]),
    .sum(sum_13[32]));
  AL_FADD comp13_33 (
    .a(i13[33]),
    .b(sum_12[33]),
    .c(cout_13[32]),
    .cout(cout_13[33]),
    .sum(sum_13[33]));
  AL_FADD comp13_34 (
    .a(1'b0),
    .b(sum_12[34]),
    .c(cout_13[33]),
    .cout(cout_13[34]),
    .sum(sum_13[34]));
  AL_FADD comp13_35 (
    .a(1'b0),
    .b(sum_12[35]),
    .c(cout_13[34]),
    .cout(cout_13[35]),
    .sum(sum_13[35]));
  AL_FADD comp13_36 (
    .a(1'b0),
    .b(sum_12[36]),
    .c(cout_13[35]),
    .cout(cout_13[36]),
    .sum(sum_13[36]));
  AL_FADD comp13_37 (
    .a(1'b0),
    .b(sum_12[37]),
    .c(cout_13[36]),
    .cout(cout_13[37]),
    .sum(sum_13[37]));
  AL_FADD comp13_38 (
    .a(1'b0),
    .b(sum_12[38]),
    .c(cout_13[37]),
    .cout(cout_13[38]),
    .sum(sum_13[38]));
  AL_FADD comp13_39 (
    .a(1'b0),
    .b(sum_12[39]),
    .c(cout_13[38]),
    .cout(cout_13[39]),
    .sum(sum_13[39]));
  AL_FADD comp13_4 (
    .a(i13[4]),
    .b(sum_12[4]),
    .c(cout_13[3]),
    .cout(cout_13[4]),
    .sum(sum_13[4]));
  AL_FADD comp13_40 (
    .a(1'b0),
    .b(sum_12[40]),
    .c(cout_13[39]),
    .cout(cout_13[40]),
    .sum(sum_13[40]));
  AL_FADD comp13_41 (
    .a(1'b0),
    .b(sum_12[41]),
    .c(cout_13[40]),
    .cout(cout_13[41]),
    .sum(sum_13[41]));
  AL_FADD comp13_42 (
    .a(1'b0),
    .b(sum_12[42]),
    .c(cout_13[41]),
    .cout(cout_13[42]),
    .sum(sum_13[42]));
  AL_FADD comp13_43 (
    .a(1'b0),
    .b(sum_12[43]),
    .c(cout_13[42]),
    .cout(cout_13[43]),
    .sum(sum_13[43]));
  AL_FADD comp13_44 (
    .a(1'b0),
    .b(sum_12[44]),
    .c(cout_13[43]),
    .cout(cout_13[44]),
    .sum(sum_13[44]));
  AL_FADD comp13_45 (
    .a(1'b0),
    .b(sum_12[45]),
    .c(cout_13[44]),
    .cout(cout_13[45]),
    .sum(sum_13[45]));
  AL_FADD comp13_46 (
    .a(1'b0),
    .b(sum_12[46]),
    .c(cout_13[45]),
    .cout(cout_13[46]),
    .sum(sum_13[46]));
  AL_FADD comp13_47 (
    .a(1'b0),
    .b(sum_12[47]),
    .c(cout_13[46]),
    .cout(cout_13[47]),
    .sum(sum_13[47]));
  AL_FADD comp13_5 (
    .a(i13[5]),
    .b(sum_12[5]),
    .c(cout_13[4]),
    .cout(cout_13[5]),
    .sum(sum_13[5]));
  AL_FADD comp13_6 (
    .a(i13[6]),
    .b(sum_12[6]),
    .c(cout_13[5]),
    .cout(cout_13[6]),
    .sum(sum_13[6]));
  AL_FADD comp13_7 (
    .a(i13[7]),
    .b(sum_12[7]),
    .c(cout_13[6]),
    .cout(cout_13[7]),
    .sum(sum_13[7]));
  AL_FADD comp13_8 (
    .a(i13[8]),
    .b(sum_12[8]),
    .c(cout_13[7]),
    .cout(cout_13[8]),
    .sum(sum_13[8]));
  AL_FADD comp13_9 (
    .a(i13[9]),
    .b(sum_12[9]),
    .c(cout_13[8]),
    .cout(cout_13[9]),
    .sum(sum_13[9]));
  AL_FADD comp14_0 (
    .a(i14[0]),
    .b(sum_13[0]),
    .c(1'b0),
    .cout(cout_14[0]),
    .sum(sum_14[0]));
  AL_FADD comp14_1 (
    .a(i14[1]),
    .b(sum_13[1]),
    .c(cout_14[0]),
    .cout(cout_14[1]),
    .sum(sum_14[1]));
  AL_FADD comp14_10 (
    .a(i14[10]),
    .b(sum_13[10]),
    .c(cout_14[9]),
    .cout(cout_14[10]),
    .sum(sum_14[10]));
  AL_FADD comp14_11 (
    .a(i14[11]),
    .b(sum_13[11]),
    .c(cout_14[10]),
    .cout(cout_14[11]),
    .sum(sum_14[11]));
  AL_FADD comp14_12 (
    .a(i14[12]),
    .b(sum_13[12]),
    .c(cout_14[11]),
    .cout(cout_14[12]),
    .sum(sum_14[12]));
  AL_FADD comp14_13 (
    .a(i14[13]),
    .b(sum_13[13]),
    .c(cout_14[12]),
    .cout(cout_14[13]),
    .sum(sum_14[13]));
  AL_FADD comp14_14 (
    .a(i14[14]),
    .b(sum_13[14]),
    .c(cout_14[13]),
    .cout(cout_14[14]),
    .sum(sum_14[14]));
  AL_FADD comp14_15 (
    .a(i14[15]),
    .b(sum_13[15]),
    .c(cout_14[14]),
    .cout(cout_14[15]),
    .sum(sum_14[15]));
  AL_FADD comp14_16 (
    .a(i14[16]),
    .b(sum_13[16]),
    .c(cout_14[15]),
    .cout(cout_14[16]),
    .sum(sum_14[16]));
  AL_FADD comp14_17 (
    .a(i14[17]),
    .b(sum_13[17]),
    .c(cout_14[16]),
    .cout(cout_14[17]),
    .sum(sum_14[17]));
  AL_FADD comp14_18 (
    .a(i14[18]),
    .b(sum_13[18]),
    .c(cout_14[17]),
    .cout(cout_14[18]),
    .sum(sum_14[18]));
  AL_FADD comp14_19 (
    .a(i14[19]),
    .b(sum_13[19]),
    .c(cout_14[18]),
    .cout(cout_14[19]),
    .sum(sum_14[19]));
  AL_FADD comp14_2 (
    .a(i14[2]),
    .b(sum_13[2]),
    .c(cout_14[1]),
    .cout(cout_14[2]),
    .sum(sum_14[2]));
  AL_FADD comp14_20 (
    .a(i14[20]),
    .b(sum_13[20]),
    .c(cout_14[19]),
    .cout(cout_14[20]),
    .sum(sum_14[20]));
  AL_FADD comp14_21 (
    .a(i14[21]),
    .b(sum_13[21]),
    .c(cout_14[20]),
    .cout(cout_14[21]),
    .sum(sum_14[21]));
  AL_FADD comp14_22 (
    .a(i14[22]),
    .b(sum_13[22]),
    .c(cout_14[21]),
    .cout(cout_14[22]),
    .sum(sum_14[22]));
  AL_FADD comp14_23 (
    .a(i14[23]),
    .b(sum_13[23]),
    .c(cout_14[22]),
    .cout(cout_14[23]),
    .sum(sum_14[23]));
  AL_FADD comp14_24 (
    .a(i14[24]),
    .b(sum_13[24]),
    .c(cout_14[23]),
    .cout(cout_14[24]),
    .sum(sum_14[24]));
  AL_FADD comp14_25 (
    .a(i14[25]),
    .b(sum_13[25]),
    .c(cout_14[24]),
    .cout(cout_14[25]),
    .sum(sum_14[25]));
  AL_FADD comp14_26 (
    .a(i14[26]),
    .b(sum_13[26]),
    .c(cout_14[25]),
    .cout(cout_14[26]),
    .sum(sum_14[26]));
  AL_FADD comp14_27 (
    .a(i14[27]),
    .b(sum_13[27]),
    .c(cout_14[26]),
    .cout(cout_14[27]),
    .sum(sum_14[27]));
  AL_FADD comp14_28 (
    .a(i14[28]),
    .b(sum_13[28]),
    .c(cout_14[27]),
    .cout(cout_14[28]),
    .sum(sum_14[28]));
  AL_FADD comp14_29 (
    .a(i14[29]),
    .b(sum_13[29]),
    .c(cout_14[28]),
    .cout(cout_14[29]),
    .sum(sum_14[29]));
  AL_FADD comp14_3 (
    .a(i14[3]),
    .b(sum_13[3]),
    .c(cout_14[2]),
    .cout(cout_14[3]),
    .sum(sum_14[3]));
  AL_FADD comp14_30 (
    .a(i14[30]),
    .b(sum_13[30]),
    .c(cout_14[29]),
    .cout(cout_14[30]),
    .sum(sum_14[30]));
  AL_FADD comp14_31 (
    .a(i14[31]),
    .b(sum_13[31]),
    .c(cout_14[30]),
    .cout(cout_14[31]),
    .sum(sum_14[31]));
  AL_FADD comp14_32 (
    .a(i14[32]),
    .b(sum_13[32]),
    .c(cout_14[31]),
    .cout(cout_14[32]),
    .sum(sum_14[32]));
  AL_FADD comp14_33 (
    .a(1'b0),
    .b(sum_13[33]),
    .c(cout_14[32]),
    .cout(cout_14[33]),
    .sum(sum_14[33]));
  AL_FADD comp14_34 (
    .a(1'b0),
    .b(sum_13[34]),
    .c(cout_14[33]),
    .cout(cout_14[34]),
    .sum(sum_14[34]));
  AL_FADD comp14_35 (
    .a(1'b0),
    .b(sum_13[35]),
    .c(cout_14[34]),
    .cout(cout_14[35]),
    .sum(sum_14[35]));
  AL_FADD comp14_36 (
    .a(1'b0),
    .b(sum_13[36]),
    .c(cout_14[35]),
    .cout(cout_14[36]),
    .sum(sum_14[36]));
  AL_FADD comp14_37 (
    .a(1'b0),
    .b(sum_13[37]),
    .c(cout_14[36]),
    .cout(cout_14[37]),
    .sum(sum_14[37]));
  AL_FADD comp14_38 (
    .a(1'b0),
    .b(sum_13[38]),
    .c(cout_14[37]),
    .cout(cout_14[38]),
    .sum(sum_14[38]));
  AL_FADD comp14_39 (
    .a(1'b0),
    .b(sum_13[39]),
    .c(cout_14[38]),
    .cout(cout_14[39]),
    .sum(sum_14[39]));
  AL_FADD comp14_4 (
    .a(i14[4]),
    .b(sum_13[4]),
    .c(cout_14[3]),
    .cout(cout_14[4]),
    .sum(sum_14[4]));
  AL_FADD comp14_40 (
    .a(1'b0),
    .b(sum_13[40]),
    .c(cout_14[39]),
    .cout(cout_14[40]),
    .sum(sum_14[40]));
  AL_FADD comp14_41 (
    .a(1'b0),
    .b(sum_13[41]),
    .c(cout_14[40]),
    .cout(cout_14[41]),
    .sum(sum_14[41]));
  AL_FADD comp14_42 (
    .a(1'b0),
    .b(sum_13[42]),
    .c(cout_14[41]),
    .cout(cout_14[42]),
    .sum(sum_14[42]));
  AL_FADD comp14_43 (
    .a(1'b0),
    .b(sum_13[43]),
    .c(cout_14[42]),
    .cout(cout_14[43]),
    .sum(sum_14[43]));
  AL_FADD comp14_44 (
    .a(1'b0),
    .b(sum_13[44]),
    .c(cout_14[43]),
    .cout(cout_14[44]),
    .sum(sum_14[44]));
  AL_FADD comp14_45 (
    .a(1'b0),
    .b(sum_13[45]),
    .c(cout_14[44]),
    .cout(cout_14[45]),
    .sum(sum_14[45]));
  AL_FADD comp14_46 (
    .a(1'b0),
    .b(sum_13[46]),
    .c(cout_14[45]),
    .cout(cout_14[46]),
    .sum(sum_14[46]));
  AL_FADD comp14_47 (
    .a(1'b0),
    .b(sum_13[47]),
    .c(cout_14[46]),
    .cout(cout_14[47]),
    .sum(sum_14[47]));
  AL_FADD comp14_5 (
    .a(i14[5]),
    .b(sum_13[5]),
    .c(cout_14[4]),
    .cout(cout_14[5]),
    .sum(sum_14[5]));
  AL_FADD comp14_6 (
    .a(i14[6]),
    .b(sum_13[6]),
    .c(cout_14[5]),
    .cout(cout_14[6]),
    .sum(sum_14[6]));
  AL_FADD comp14_7 (
    .a(i14[7]),
    .b(sum_13[7]),
    .c(cout_14[6]),
    .cout(cout_14[7]),
    .sum(sum_14[7]));
  AL_FADD comp14_8 (
    .a(i14[8]),
    .b(sum_13[8]),
    .c(cout_14[7]),
    .cout(cout_14[8]),
    .sum(sum_14[8]));
  AL_FADD comp14_9 (
    .a(i14[9]),
    .b(sum_13[9]),
    .c(cout_14[8]),
    .cout(cout_14[9]),
    .sum(sum_14[9]));
  AL_FADD comp15_0 (
    .a(i15[0]),
    .b(sum_14[0]),
    .c(1'b0),
    .cout(cout_15[0]),
    .sum(sum_15[0]));
  AL_FADD comp15_1 (
    .a(i15[1]),
    .b(sum_14[1]),
    .c(cout_15[0]),
    .cout(cout_15[1]),
    .sum(sum_15[1]));
  AL_FADD comp15_10 (
    .a(i15[10]),
    .b(sum_14[10]),
    .c(cout_15[9]),
    .cout(cout_15[10]),
    .sum(sum_15[10]));
  AL_FADD comp15_11 (
    .a(i15[11]),
    .b(sum_14[11]),
    .c(cout_15[10]),
    .cout(cout_15[11]),
    .sum(sum_15[11]));
  AL_FADD comp15_12 (
    .a(i15[12]),
    .b(sum_14[12]),
    .c(cout_15[11]),
    .cout(cout_15[12]),
    .sum(sum_15[12]));
  AL_FADD comp15_13 (
    .a(i15[13]),
    .b(sum_14[13]),
    .c(cout_15[12]),
    .cout(cout_15[13]),
    .sum(sum_15[13]));
  AL_FADD comp15_14 (
    .a(i15[14]),
    .b(sum_14[14]),
    .c(cout_15[13]),
    .cout(cout_15[14]),
    .sum(sum_15[14]));
  AL_FADD comp15_15 (
    .a(i15[15]),
    .b(sum_14[15]),
    .c(cout_15[14]),
    .cout(cout_15[15]),
    .sum(sum_15[15]));
  AL_FADD comp15_16 (
    .a(i15[16]),
    .b(sum_14[16]),
    .c(cout_15[15]),
    .cout(cout_15[16]),
    .sum(sum_15[16]));
  AL_FADD comp15_17 (
    .a(i15[17]),
    .b(sum_14[17]),
    .c(cout_15[16]),
    .cout(cout_15[17]),
    .sum(sum_15[17]));
  AL_FADD comp15_18 (
    .a(i15[18]),
    .b(sum_14[18]),
    .c(cout_15[17]),
    .cout(cout_15[18]),
    .sum(sum_15[18]));
  AL_FADD comp15_19 (
    .a(i15[19]),
    .b(sum_14[19]),
    .c(cout_15[18]),
    .cout(cout_15[19]),
    .sum(sum_15[19]));
  AL_FADD comp15_2 (
    .a(i15[2]),
    .b(sum_14[2]),
    .c(cout_15[1]),
    .cout(cout_15[2]),
    .sum(sum_15[2]));
  AL_FADD comp15_20 (
    .a(i15[20]),
    .b(sum_14[20]),
    .c(cout_15[19]),
    .cout(cout_15[20]),
    .sum(sum_15[20]));
  AL_FADD comp15_21 (
    .a(i15[21]),
    .b(sum_14[21]),
    .c(cout_15[20]),
    .cout(cout_15[21]),
    .sum(sum_15[21]));
  AL_FADD comp15_22 (
    .a(i15[22]),
    .b(sum_14[22]),
    .c(cout_15[21]),
    .cout(cout_15[22]),
    .sum(sum_15[22]));
  AL_FADD comp15_23 (
    .a(i15[23]),
    .b(sum_14[23]),
    .c(cout_15[22]),
    .cout(cout_15[23]),
    .sum(sum_15[23]));
  AL_FADD comp15_24 (
    .a(i15[24]),
    .b(sum_14[24]),
    .c(cout_15[23]),
    .cout(cout_15[24]),
    .sum(sum_15[24]));
  AL_FADD comp15_25 (
    .a(i15[25]),
    .b(sum_14[25]),
    .c(cout_15[24]),
    .cout(cout_15[25]),
    .sum(sum_15[25]));
  AL_FADD comp15_26 (
    .a(i15[26]),
    .b(sum_14[26]),
    .c(cout_15[25]),
    .cout(cout_15[26]),
    .sum(sum_15[26]));
  AL_FADD comp15_27 (
    .a(i15[27]),
    .b(sum_14[27]),
    .c(cout_15[26]),
    .cout(cout_15[27]),
    .sum(sum_15[27]));
  AL_FADD comp15_28 (
    .a(i15[28]),
    .b(sum_14[28]),
    .c(cout_15[27]),
    .cout(cout_15[28]),
    .sum(sum_15[28]));
  AL_FADD comp15_29 (
    .a(i15[29]),
    .b(sum_14[29]),
    .c(cout_15[28]),
    .cout(cout_15[29]),
    .sum(sum_15[29]));
  AL_FADD comp15_3 (
    .a(i15[3]),
    .b(sum_14[3]),
    .c(cout_15[2]),
    .cout(cout_15[3]),
    .sum(sum_15[3]));
  AL_FADD comp15_30 (
    .a(i15[30]),
    .b(sum_14[30]),
    .c(cout_15[29]),
    .cout(cout_15[30]),
    .sum(sum_15[30]));
  AL_FADD comp15_31 (
    .a(i15[31]),
    .b(sum_14[31]),
    .c(cout_15[30]),
    .cout(cout_15[31]),
    .sum(sum_15[31]));
  AL_FADD comp15_32 (
    .a(1'b0),
    .b(sum_14[32]),
    .c(cout_15[31]),
    .cout(cout_15[32]),
    .sum(sum_15[32]));
  AL_FADD comp15_33 (
    .a(1'b0),
    .b(sum_14[33]),
    .c(cout_15[32]),
    .cout(cout_15[33]),
    .sum(sum_15[33]));
  AL_FADD comp15_34 (
    .a(1'b0),
    .b(sum_14[34]),
    .c(cout_15[33]),
    .cout(cout_15[34]),
    .sum(sum_15[34]));
  AL_FADD comp15_35 (
    .a(1'b0),
    .b(sum_14[35]),
    .c(cout_15[34]),
    .cout(cout_15[35]),
    .sum(sum_15[35]));
  AL_FADD comp15_36 (
    .a(1'b0),
    .b(sum_14[36]),
    .c(cout_15[35]),
    .cout(cout_15[36]),
    .sum(sum_15[36]));
  AL_FADD comp15_37 (
    .a(1'b0),
    .b(sum_14[37]),
    .c(cout_15[36]),
    .cout(cout_15[37]),
    .sum(sum_15[37]));
  AL_FADD comp15_38 (
    .a(1'b0),
    .b(sum_14[38]),
    .c(cout_15[37]),
    .cout(cout_15[38]),
    .sum(sum_15[38]));
  AL_FADD comp15_39 (
    .a(1'b0),
    .b(sum_14[39]),
    .c(cout_15[38]),
    .cout(cout_15[39]),
    .sum(sum_15[39]));
  AL_FADD comp15_4 (
    .a(i15[4]),
    .b(sum_14[4]),
    .c(cout_15[3]),
    .cout(cout_15[4]),
    .sum(sum_15[4]));
  AL_FADD comp15_40 (
    .a(1'b0),
    .b(sum_14[40]),
    .c(cout_15[39]),
    .cout(cout_15[40]),
    .sum(sum_15[40]));
  AL_FADD comp15_41 (
    .a(1'b0),
    .b(sum_14[41]),
    .c(cout_15[40]),
    .cout(cout_15[41]),
    .sum(sum_15[41]));
  AL_FADD comp15_42 (
    .a(1'b0),
    .b(sum_14[42]),
    .c(cout_15[41]),
    .cout(cout_15[42]),
    .sum(sum_15[42]));
  AL_FADD comp15_43 (
    .a(1'b0),
    .b(sum_14[43]),
    .c(cout_15[42]),
    .cout(cout_15[43]),
    .sum(sum_15[43]));
  AL_FADD comp15_44 (
    .a(1'b0),
    .b(sum_14[44]),
    .c(cout_15[43]),
    .cout(cout_15[44]),
    .sum(sum_15[44]));
  AL_FADD comp15_45 (
    .a(1'b0),
    .b(sum_14[45]),
    .c(cout_15[44]),
    .cout(cout_15[45]),
    .sum(sum_15[45]));
  AL_FADD comp15_46 (
    .a(1'b0),
    .b(sum_14[46]),
    .c(cout_15[45]),
    .cout(cout_15[46]),
    .sum(sum_15[46]));
  AL_FADD comp15_47 (
    .a(1'b0),
    .b(sum_14[47]),
    .c(cout_15[46]),
    .cout(cout_15[47]),
    .sum(sum_15[47]));
  AL_FADD comp15_5 (
    .a(i15[5]),
    .b(sum_14[5]),
    .c(cout_15[4]),
    .cout(cout_15[5]),
    .sum(sum_15[5]));
  AL_FADD comp15_6 (
    .a(i15[6]),
    .b(sum_14[6]),
    .c(cout_15[5]),
    .cout(cout_15[6]),
    .sum(sum_15[6]));
  AL_FADD comp15_7 (
    .a(i15[7]),
    .b(sum_14[7]),
    .c(cout_15[6]),
    .cout(cout_15[7]),
    .sum(sum_15[7]));
  AL_FADD comp15_8 (
    .a(i15[8]),
    .b(sum_14[8]),
    .c(cout_15[7]),
    .cout(cout_15[8]),
    .sum(sum_15[8]));
  AL_FADD comp15_9 (
    .a(i15[9]),
    .b(sum_14[9]),
    .c(cout_15[8]),
    .cout(cout_15[9]),
    .sum(sum_15[9]));
  AL_FADD comp16_0 (
    .a(i16[0]),
    .b(sum_15[0]),
    .c(1'b0),
    .cout(cout_16[0]),
    .sum(sum_16[0]));
  AL_FADD comp16_1 (
    .a(i16[1]),
    .b(sum_15[1]),
    .c(cout_16[0]),
    .cout(cout_16[1]),
    .sum(sum_16[1]));
  AL_FADD comp16_10 (
    .a(i16[10]),
    .b(sum_15[10]),
    .c(cout_16[9]),
    .cout(cout_16[10]),
    .sum(sum_16[10]));
  AL_FADD comp16_11 (
    .a(i16[11]),
    .b(sum_15[11]),
    .c(cout_16[10]),
    .cout(cout_16[11]),
    .sum(sum_16[11]));
  AL_FADD comp16_12 (
    .a(i16[12]),
    .b(sum_15[12]),
    .c(cout_16[11]),
    .cout(cout_16[12]),
    .sum(sum_16[12]));
  AL_FADD comp16_13 (
    .a(i16[13]),
    .b(sum_15[13]),
    .c(cout_16[12]),
    .cout(cout_16[13]),
    .sum(sum_16[13]));
  AL_FADD comp16_14 (
    .a(i16[14]),
    .b(sum_15[14]),
    .c(cout_16[13]),
    .cout(cout_16[14]),
    .sum(sum_16[14]));
  AL_FADD comp16_15 (
    .a(i16[15]),
    .b(sum_15[15]),
    .c(cout_16[14]),
    .cout(cout_16[15]),
    .sum(sum_16[15]));
  AL_FADD comp16_16 (
    .a(i16[16]),
    .b(sum_15[16]),
    .c(cout_16[15]),
    .cout(cout_16[16]),
    .sum(sum_16[16]));
  AL_FADD comp16_17 (
    .a(i16[17]),
    .b(sum_15[17]),
    .c(cout_16[16]),
    .cout(cout_16[17]),
    .sum(sum_16[17]));
  AL_FADD comp16_18 (
    .a(i16[18]),
    .b(sum_15[18]),
    .c(cout_16[17]),
    .cout(cout_16[18]),
    .sum(sum_16[18]));
  AL_FADD comp16_19 (
    .a(i16[19]),
    .b(sum_15[19]),
    .c(cout_16[18]),
    .cout(cout_16[19]),
    .sum(sum_16[19]));
  AL_FADD comp16_2 (
    .a(i16[2]),
    .b(sum_15[2]),
    .c(cout_16[1]),
    .cout(cout_16[2]),
    .sum(sum_16[2]));
  AL_FADD comp16_20 (
    .a(i16[20]),
    .b(sum_15[20]),
    .c(cout_16[19]),
    .cout(cout_16[20]),
    .sum(sum_16[20]));
  AL_FADD comp16_21 (
    .a(i16[21]),
    .b(sum_15[21]),
    .c(cout_16[20]),
    .cout(cout_16[21]),
    .sum(sum_16[21]));
  AL_FADD comp16_22 (
    .a(i16[22]),
    .b(sum_15[22]),
    .c(cout_16[21]),
    .cout(cout_16[22]),
    .sum(sum_16[22]));
  AL_FADD comp16_23 (
    .a(i16[23]),
    .b(sum_15[23]),
    .c(cout_16[22]),
    .cout(cout_16[23]),
    .sum(sum_16[23]));
  AL_FADD comp16_24 (
    .a(i16[24]),
    .b(sum_15[24]),
    .c(cout_16[23]),
    .cout(cout_16[24]),
    .sum(sum_16[24]));
  AL_FADD comp16_25 (
    .a(i16[25]),
    .b(sum_15[25]),
    .c(cout_16[24]),
    .cout(cout_16[25]),
    .sum(sum_16[25]));
  AL_FADD comp16_26 (
    .a(i16[26]),
    .b(sum_15[26]),
    .c(cout_16[25]),
    .cout(cout_16[26]),
    .sum(sum_16[26]));
  AL_FADD comp16_27 (
    .a(i16[27]),
    .b(sum_15[27]),
    .c(cout_16[26]),
    .cout(cout_16[27]),
    .sum(sum_16[27]));
  AL_FADD comp16_28 (
    .a(i16[28]),
    .b(sum_15[28]),
    .c(cout_16[27]),
    .cout(cout_16[28]),
    .sum(sum_16[28]));
  AL_FADD comp16_29 (
    .a(i16[29]),
    .b(sum_15[29]),
    .c(cout_16[28]),
    .cout(cout_16[29]),
    .sum(sum_16[29]));
  AL_FADD comp16_3 (
    .a(i16[3]),
    .b(sum_15[3]),
    .c(cout_16[2]),
    .cout(cout_16[3]),
    .sum(sum_16[3]));
  AL_FADD comp16_30 (
    .a(i16[30]),
    .b(sum_15[30]),
    .c(cout_16[29]),
    .cout(cout_16[30]),
    .sum(sum_16[30]));
  AL_FADD comp16_31 (
    .a(1'b0),
    .b(sum_15[31]),
    .c(cout_16[30]),
    .cout(cout_16[31]),
    .sum(sum_16[31]));
  AL_FADD comp16_32 (
    .a(1'b0),
    .b(sum_15[32]),
    .c(cout_16[31]),
    .cout(cout_16[32]),
    .sum(sum_16[32]));
  AL_FADD comp16_33 (
    .a(1'b0),
    .b(sum_15[33]),
    .c(cout_16[32]),
    .cout(cout_16[33]),
    .sum(sum_16[33]));
  AL_FADD comp16_34 (
    .a(1'b0),
    .b(sum_15[34]),
    .c(cout_16[33]),
    .cout(cout_16[34]),
    .sum(sum_16[34]));
  AL_FADD comp16_35 (
    .a(1'b0),
    .b(sum_15[35]),
    .c(cout_16[34]),
    .cout(cout_16[35]),
    .sum(sum_16[35]));
  AL_FADD comp16_36 (
    .a(1'b0),
    .b(sum_15[36]),
    .c(cout_16[35]),
    .cout(cout_16[36]),
    .sum(sum_16[36]));
  AL_FADD comp16_37 (
    .a(1'b0),
    .b(sum_15[37]),
    .c(cout_16[36]),
    .cout(cout_16[37]),
    .sum(sum_16[37]));
  AL_FADD comp16_38 (
    .a(1'b0),
    .b(sum_15[38]),
    .c(cout_16[37]),
    .cout(cout_16[38]),
    .sum(sum_16[38]));
  AL_FADD comp16_39 (
    .a(1'b0),
    .b(sum_15[39]),
    .c(cout_16[38]),
    .cout(cout_16[39]),
    .sum(sum_16[39]));
  AL_FADD comp16_4 (
    .a(i16[4]),
    .b(sum_15[4]),
    .c(cout_16[3]),
    .cout(cout_16[4]),
    .sum(sum_16[4]));
  AL_FADD comp16_40 (
    .a(1'b0),
    .b(sum_15[40]),
    .c(cout_16[39]),
    .cout(cout_16[40]),
    .sum(sum_16[40]));
  AL_FADD comp16_41 (
    .a(1'b0),
    .b(sum_15[41]),
    .c(cout_16[40]),
    .cout(cout_16[41]),
    .sum(sum_16[41]));
  AL_FADD comp16_42 (
    .a(1'b0),
    .b(sum_15[42]),
    .c(cout_16[41]),
    .cout(cout_16[42]),
    .sum(sum_16[42]));
  AL_FADD comp16_43 (
    .a(1'b0),
    .b(sum_15[43]),
    .c(cout_16[42]),
    .cout(cout_16[43]),
    .sum(sum_16[43]));
  AL_FADD comp16_44 (
    .a(1'b0),
    .b(sum_15[44]),
    .c(cout_16[43]),
    .cout(cout_16[44]),
    .sum(sum_16[44]));
  AL_FADD comp16_45 (
    .a(1'b0),
    .b(sum_15[45]),
    .c(cout_16[44]),
    .cout(cout_16[45]),
    .sum(sum_16[45]));
  AL_FADD comp16_46 (
    .a(1'b0),
    .b(sum_15[46]),
    .c(cout_16[45]),
    .cout(cout_16[46]),
    .sum(sum_16[46]));
  AL_FADD comp16_47 (
    .a(1'b0),
    .b(sum_15[47]),
    .c(cout_16[46]),
    .cout(cout_16[47]),
    .sum(sum_16[47]));
  AL_FADD comp16_5 (
    .a(i16[5]),
    .b(sum_15[5]),
    .c(cout_16[4]),
    .cout(cout_16[5]),
    .sum(sum_16[5]));
  AL_FADD comp16_6 (
    .a(i16[6]),
    .b(sum_15[6]),
    .c(cout_16[5]),
    .cout(cout_16[6]),
    .sum(sum_16[6]));
  AL_FADD comp16_7 (
    .a(i16[7]),
    .b(sum_15[7]),
    .c(cout_16[6]),
    .cout(cout_16[7]),
    .sum(sum_16[7]));
  AL_FADD comp16_8 (
    .a(i16[8]),
    .b(sum_15[8]),
    .c(cout_16[7]),
    .cout(cout_16[8]),
    .sum(sum_16[8]));
  AL_FADD comp16_9 (
    .a(i16[9]),
    .b(sum_15[9]),
    .c(cout_16[8]),
    .cout(cout_16[9]),
    .sum(sum_16[9]));
  AL_FADD comp17_0 (
    .a(i17[0]),
    .b(sum_16[0]),
    .c(1'b0),
    .cout(cout_17[0]),
    .sum(sum_17[0]));
  AL_FADD comp17_1 (
    .a(i17[1]),
    .b(sum_16[1]),
    .c(cout_17[0]),
    .cout(cout_17[1]),
    .sum(sum_17[1]));
  AL_FADD comp17_10 (
    .a(i17[10]),
    .b(sum_16[10]),
    .c(cout_17[9]),
    .cout(cout_17[10]),
    .sum(sum_17[10]));
  AL_FADD comp17_11 (
    .a(i17[11]),
    .b(sum_16[11]),
    .c(cout_17[10]),
    .cout(cout_17[11]),
    .sum(sum_17[11]));
  AL_FADD comp17_12 (
    .a(i17[12]),
    .b(sum_16[12]),
    .c(cout_17[11]),
    .cout(cout_17[12]),
    .sum(sum_17[12]));
  AL_FADD comp17_13 (
    .a(i17[13]),
    .b(sum_16[13]),
    .c(cout_17[12]),
    .cout(cout_17[13]),
    .sum(sum_17[13]));
  AL_FADD comp17_14 (
    .a(i17[14]),
    .b(sum_16[14]),
    .c(cout_17[13]),
    .cout(cout_17[14]),
    .sum(sum_17[14]));
  AL_FADD comp17_15 (
    .a(i17[15]),
    .b(sum_16[15]),
    .c(cout_17[14]),
    .cout(cout_17[15]),
    .sum(sum_17[15]));
  AL_FADD comp17_16 (
    .a(i17[16]),
    .b(sum_16[16]),
    .c(cout_17[15]),
    .cout(cout_17[16]),
    .sum(sum_17[16]));
  AL_FADD comp17_17 (
    .a(i17[17]),
    .b(sum_16[17]),
    .c(cout_17[16]),
    .cout(cout_17[17]),
    .sum(sum_17[17]));
  AL_FADD comp17_18 (
    .a(i17[18]),
    .b(sum_16[18]),
    .c(cout_17[17]),
    .cout(cout_17[18]),
    .sum(sum_17[18]));
  AL_FADD comp17_19 (
    .a(i17[19]),
    .b(sum_16[19]),
    .c(cout_17[18]),
    .cout(cout_17[19]),
    .sum(sum_17[19]));
  AL_FADD comp17_2 (
    .a(i17[2]),
    .b(sum_16[2]),
    .c(cout_17[1]),
    .cout(cout_17[2]),
    .sum(sum_17[2]));
  AL_FADD comp17_20 (
    .a(i17[20]),
    .b(sum_16[20]),
    .c(cout_17[19]),
    .cout(cout_17[20]),
    .sum(sum_17[20]));
  AL_FADD comp17_21 (
    .a(i17[21]),
    .b(sum_16[21]),
    .c(cout_17[20]),
    .cout(cout_17[21]),
    .sum(sum_17[21]));
  AL_FADD comp17_22 (
    .a(i17[22]),
    .b(sum_16[22]),
    .c(cout_17[21]),
    .cout(cout_17[22]),
    .sum(sum_17[22]));
  AL_FADD comp17_23 (
    .a(i17[23]),
    .b(sum_16[23]),
    .c(cout_17[22]),
    .cout(cout_17[23]),
    .sum(sum_17[23]));
  AL_FADD comp17_24 (
    .a(i17[24]),
    .b(sum_16[24]),
    .c(cout_17[23]),
    .cout(cout_17[24]),
    .sum(sum_17[24]));
  AL_FADD comp17_25 (
    .a(i17[25]),
    .b(sum_16[25]),
    .c(cout_17[24]),
    .cout(cout_17[25]),
    .sum(sum_17[25]));
  AL_FADD comp17_26 (
    .a(i17[26]),
    .b(sum_16[26]),
    .c(cout_17[25]),
    .cout(cout_17[26]),
    .sum(sum_17[26]));
  AL_FADD comp17_27 (
    .a(i17[27]),
    .b(sum_16[27]),
    .c(cout_17[26]),
    .cout(cout_17[27]),
    .sum(sum_17[27]));
  AL_FADD comp17_28 (
    .a(i17[28]),
    .b(sum_16[28]),
    .c(cout_17[27]),
    .cout(cout_17[28]),
    .sum(sum_17[28]));
  AL_FADD comp17_29 (
    .a(i17[29]),
    .b(sum_16[29]),
    .c(cout_17[28]),
    .cout(cout_17[29]),
    .sum(sum_17[29]));
  AL_FADD comp17_3 (
    .a(i17[3]),
    .b(sum_16[3]),
    .c(cout_17[2]),
    .cout(cout_17[3]),
    .sum(sum_17[3]));
  AL_FADD comp17_30 (
    .a(1'b0),
    .b(sum_16[30]),
    .c(cout_17[29]),
    .cout(cout_17[30]),
    .sum(sum_17[30]));
  AL_FADD comp17_31 (
    .a(1'b0),
    .b(sum_16[31]),
    .c(cout_17[30]),
    .cout(cout_17[31]),
    .sum(sum_17[31]));
  AL_FADD comp17_32 (
    .a(1'b0),
    .b(sum_16[32]),
    .c(cout_17[31]),
    .cout(cout_17[32]),
    .sum(sum_17[32]));
  AL_FADD comp17_33 (
    .a(1'b0),
    .b(sum_16[33]),
    .c(cout_17[32]),
    .cout(cout_17[33]),
    .sum(sum_17[33]));
  AL_FADD comp17_34 (
    .a(1'b0),
    .b(sum_16[34]),
    .c(cout_17[33]),
    .cout(cout_17[34]),
    .sum(sum_17[34]));
  AL_FADD comp17_35 (
    .a(1'b0),
    .b(sum_16[35]),
    .c(cout_17[34]),
    .cout(cout_17[35]),
    .sum(sum_17[35]));
  AL_FADD comp17_36 (
    .a(1'b0),
    .b(sum_16[36]),
    .c(cout_17[35]),
    .cout(cout_17[36]),
    .sum(sum_17[36]));
  AL_FADD comp17_37 (
    .a(1'b0),
    .b(sum_16[37]),
    .c(cout_17[36]),
    .cout(cout_17[37]),
    .sum(sum_17[37]));
  AL_FADD comp17_38 (
    .a(1'b0),
    .b(sum_16[38]),
    .c(cout_17[37]),
    .cout(cout_17[38]),
    .sum(sum_17[38]));
  AL_FADD comp17_39 (
    .a(1'b0),
    .b(sum_16[39]),
    .c(cout_17[38]),
    .cout(cout_17[39]),
    .sum(sum_17[39]));
  AL_FADD comp17_4 (
    .a(i17[4]),
    .b(sum_16[4]),
    .c(cout_17[3]),
    .cout(cout_17[4]),
    .sum(sum_17[4]));
  AL_FADD comp17_40 (
    .a(1'b0),
    .b(sum_16[40]),
    .c(cout_17[39]),
    .cout(cout_17[40]),
    .sum(sum_17[40]));
  AL_FADD comp17_41 (
    .a(1'b0),
    .b(sum_16[41]),
    .c(cout_17[40]),
    .cout(cout_17[41]),
    .sum(sum_17[41]));
  AL_FADD comp17_42 (
    .a(1'b0),
    .b(sum_16[42]),
    .c(cout_17[41]),
    .cout(cout_17[42]),
    .sum(sum_17[42]));
  AL_FADD comp17_43 (
    .a(1'b0),
    .b(sum_16[43]),
    .c(cout_17[42]),
    .cout(cout_17[43]),
    .sum(sum_17[43]));
  AL_FADD comp17_44 (
    .a(1'b0),
    .b(sum_16[44]),
    .c(cout_17[43]),
    .cout(cout_17[44]),
    .sum(sum_17[44]));
  AL_FADD comp17_45 (
    .a(1'b0),
    .b(sum_16[45]),
    .c(cout_17[44]),
    .cout(cout_17[45]),
    .sum(sum_17[45]));
  AL_FADD comp17_46 (
    .a(1'b0),
    .b(sum_16[46]),
    .c(cout_17[45]),
    .cout(cout_17[46]),
    .sum(sum_17[46]));
  AL_FADD comp17_47 (
    .a(1'b0),
    .b(sum_16[47]),
    .c(cout_17[46]),
    .cout(cout_17[47]),
    .sum(sum_17[47]));
  AL_FADD comp17_5 (
    .a(i17[5]),
    .b(sum_16[5]),
    .c(cout_17[4]),
    .cout(cout_17[5]),
    .sum(sum_17[5]));
  AL_FADD comp17_6 (
    .a(i17[6]),
    .b(sum_16[6]),
    .c(cout_17[5]),
    .cout(cout_17[6]),
    .sum(sum_17[6]));
  AL_FADD comp17_7 (
    .a(i17[7]),
    .b(sum_16[7]),
    .c(cout_17[6]),
    .cout(cout_17[7]),
    .sum(sum_17[7]));
  AL_FADD comp17_8 (
    .a(i17[8]),
    .b(sum_16[8]),
    .c(cout_17[7]),
    .cout(cout_17[8]),
    .sum(sum_17[8]));
  AL_FADD comp17_9 (
    .a(i17[9]),
    .b(sum_16[9]),
    .c(cout_17[8]),
    .cout(cout_17[9]),
    .sum(sum_17[9]));
  AL_FADD comp18_0 (
    .a(i18[0]),
    .b(sum_17[0]),
    .c(1'b0),
    .cout(cout_18[0]),
    .sum(sum_18[0]));
  AL_FADD comp18_1 (
    .a(i18[1]),
    .b(sum_17[1]),
    .c(cout_18[0]),
    .cout(cout_18[1]),
    .sum(sum_18[1]));
  AL_FADD comp18_10 (
    .a(i18[10]),
    .b(sum_17[10]),
    .c(cout_18[9]),
    .cout(cout_18[10]),
    .sum(sum_18[10]));
  AL_FADD comp18_11 (
    .a(i18[11]),
    .b(sum_17[11]),
    .c(cout_18[10]),
    .cout(cout_18[11]),
    .sum(sum_18[11]));
  AL_FADD comp18_12 (
    .a(i18[12]),
    .b(sum_17[12]),
    .c(cout_18[11]),
    .cout(cout_18[12]),
    .sum(sum_18[12]));
  AL_FADD comp18_13 (
    .a(i18[13]),
    .b(sum_17[13]),
    .c(cout_18[12]),
    .cout(cout_18[13]),
    .sum(sum_18[13]));
  AL_FADD comp18_14 (
    .a(i18[14]),
    .b(sum_17[14]),
    .c(cout_18[13]),
    .cout(cout_18[14]),
    .sum(sum_18[14]));
  AL_FADD comp18_15 (
    .a(i18[15]),
    .b(sum_17[15]),
    .c(cout_18[14]),
    .cout(cout_18[15]),
    .sum(sum_18[15]));
  AL_FADD comp18_16 (
    .a(i18[16]),
    .b(sum_17[16]),
    .c(cout_18[15]),
    .cout(cout_18[16]),
    .sum(sum_18[16]));
  AL_FADD comp18_17 (
    .a(i18[17]),
    .b(sum_17[17]),
    .c(cout_18[16]),
    .cout(cout_18[17]),
    .sum(sum_18[17]));
  AL_FADD comp18_18 (
    .a(i18[18]),
    .b(sum_17[18]),
    .c(cout_18[17]),
    .cout(cout_18[18]),
    .sum(sum_18[18]));
  AL_FADD comp18_19 (
    .a(i18[19]),
    .b(sum_17[19]),
    .c(cout_18[18]),
    .cout(cout_18[19]),
    .sum(sum_18[19]));
  AL_FADD comp18_2 (
    .a(i18[2]),
    .b(sum_17[2]),
    .c(cout_18[1]),
    .cout(cout_18[2]),
    .sum(sum_18[2]));
  AL_FADD comp18_20 (
    .a(i18[20]),
    .b(sum_17[20]),
    .c(cout_18[19]),
    .cout(cout_18[20]),
    .sum(sum_18[20]));
  AL_FADD comp18_21 (
    .a(i18[21]),
    .b(sum_17[21]),
    .c(cout_18[20]),
    .cout(cout_18[21]),
    .sum(sum_18[21]));
  AL_FADD comp18_22 (
    .a(i18[22]),
    .b(sum_17[22]),
    .c(cout_18[21]),
    .cout(cout_18[22]),
    .sum(sum_18[22]));
  AL_FADD comp18_23 (
    .a(i18[23]),
    .b(sum_17[23]),
    .c(cout_18[22]),
    .cout(cout_18[23]),
    .sum(sum_18[23]));
  AL_FADD comp18_24 (
    .a(i18[24]),
    .b(sum_17[24]),
    .c(cout_18[23]),
    .cout(cout_18[24]),
    .sum(sum_18[24]));
  AL_FADD comp18_25 (
    .a(i18[25]),
    .b(sum_17[25]),
    .c(cout_18[24]),
    .cout(cout_18[25]),
    .sum(sum_18[25]));
  AL_FADD comp18_26 (
    .a(i18[26]),
    .b(sum_17[26]),
    .c(cout_18[25]),
    .cout(cout_18[26]),
    .sum(sum_18[26]));
  AL_FADD comp18_27 (
    .a(i18[27]),
    .b(sum_17[27]),
    .c(cout_18[26]),
    .cout(cout_18[27]),
    .sum(sum_18[27]));
  AL_FADD comp18_28 (
    .a(i18[28]),
    .b(sum_17[28]),
    .c(cout_18[27]),
    .cout(cout_18[28]),
    .sum(sum_18[28]));
  AL_FADD comp18_29 (
    .a(1'b0),
    .b(sum_17[29]),
    .c(cout_18[28]),
    .cout(cout_18[29]),
    .sum(sum_18[29]));
  AL_FADD comp18_3 (
    .a(i18[3]),
    .b(sum_17[3]),
    .c(cout_18[2]),
    .cout(cout_18[3]),
    .sum(sum_18[3]));
  AL_FADD comp18_30 (
    .a(1'b0),
    .b(sum_17[30]),
    .c(cout_18[29]),
    .cout(cout_18[30]),
    .sum(sum_18[30]));
  AL_FADD comp18_31 (
    .a(1'b0),
    .b(sum_17[31]),
    .c(cout_18[30]),
    .cout(cout_18[31]),
    .sum(sum_18[31]));
  AL_FADD comp18_32 (
    .a(1'b0),
    .b(sum_17[32]),
    .c(cout_18[31]),
    .cout(cout_18[32]),
    .sum(sum_18[32]));
  AL_FADD comp18_33 (
    .a(1'b0),
    .b(sum_17[33]),
    .c(cout_18[32]),
    .cout(cout_18[33]),
    .sum(sum_18[33]));
  AL_FADD comp18_34 (
    .a(1'b0),
    .b(sum_17[34]),
    .c(cout_18[33]),
    .cout(cout_18[34]),
    .sum(sum_18[34]));
  AL_FADD comp18_35 (
    .a(1'b0),
    .b(sum_17[35]),
    .c(cout_18[34]),
    .cout(cout_18[35]),
    .sum(sum_18[35]));
  AL_FADD comp18_36 (
    .a(1'b0),
    .b(sum_17[36]),
    .c(cout_18[35]),
    .cout(cout_18[36]),
    .sum(sum_18[36]));
  AL_FADD comp18_37 (
    .a(1'b0),
    .b(sum_17[37]),
    .c(cout_18[36]),
    .cout(cout_18[37]),
    .sum(sum_18[37]));
  AL_FADD comp18_38 (
    .a(1'b0),
    .b(sum_17[38]),
    .c(cout_18[37]),
    .cout(cout_18[38]),
    .sum(sum_18[38]));
  AL_FADD comp18_39 (
    .a(1'b0),
    .b(sum_17[39]),
    .c(cout_18[38]),
    .cout(cout_18[39]),
    .sum(sum_18[39]));
  AL_FADD comp18_4 (
    .a(i18[4]),
    .b(sum_17[4]),
    .c(cout_18[3]),
    .cout(cout_18[4]),
    .sum(sum_18[4]));
  AL_FADD comp18_40 (
    .a(1'b0),
    .b(sum_17[40]),
    .c(cout_18[39]),
    .cout(cout_18[40]),
    .sum(sum_18[40]));
  AL_FADD comp18_41 (
    .a(1'b0),
    .b(sum_17[41]),
    .c(cout_18[40]),
    .cout(cout_18[41]),
    .sum(sum_18[41]));
  AL_FADD comp18_42 (
    .a(1'b0),
    .b(sum_17[42]),
    .c(cout_18[41]),
    .cout(cout_18[42]),
    .sum(sum_18[42]));
  AL_FADD comp18_43 (
    .a(1'b0),
    .b(sum_17[43]),
    .c(cout_18[42]),
    .cout(cout_18[43]),
    .sum(sum_18[43]));
  AL_FADD comp18_44 (
    .a(1'b0),
    .b(sum_17[44]),
    .c(cout_18[43]),
    .cout(cout_18[44]),
    .sum(sum_18[44]));
  AL_FADD comp18_45 (
    .a(1'b0),
    .b(sum_17[45]),
    .c(cout_18[44]),
    .cout(cout_18[45]),
    .sum(sum_18[45]));
  AL_FADD comp18_46 (
    .a(1'b0),
    .b(sum_17[46]),
    .c(cout_18[45]),
    .cout(cout_18[46]),
    .sum(sum_18[46]));
  AL_FADD comp18_47 (
    .a(1'b0),
    .b(sum_17[47]),
    .c(cout_18[46]),
    .cout(cout_18[47]),
    .sum(sum_18[47]));
  AL_FADD comp18_5 (
    .a(i18[5]),
    .b(sum_17[5]),
    .c(cout_18[4]),
    .cout(cout_18[5]),
    .sum(sum_18[5]));
  AL_FADD comp18_6 (
    .a(i18[6]),
    .b(sum_17[6]),
    .c(cout_18[5]),
    .cout(cout_18[6]),
    .sum(sum_18[6]));
  AL_FADD comp18_7 (
    .a(i18[7]),
    .b(sum_17[7]),
    .c(cout_18[6]),
    .cout(cout_18[7]),
    .sum(sum_18[7]));
  AL_FADD comp18_8 (
    .a(i18[8]),
    .b(sum_17[8]),
    .c(cout_18[7]),
    .cout(cout_18[8]),
    .sum(sum_18[8]));
  AL_FADD comp18_9 (
    .a(i18[9]),
    .b(sum_17[9]),
    .c(cout_18[8]),
    .cout(cout_18[9]),
    .sum(sum_18[9]));
  AL_FADD comp19_0 (
    .a(i19[0]),
    .b(sum_18[0]),
    .c(1'b0),
    .cout(cout_19[0]),
    .sum(sum_19[0]));
  AL_FADD comp19_1 (
    .a(i19[1]),
    .b(sum_18[1]),
    .c(cout_19[0]),
    .cout(cout_19[1]),
    .sum(sum_19[1]));
  AL_FADD comp19_10 (
    .a(i19[10]),
    .b(sum_18[10]),
    .c(cout_19[9]),
    .cout(cout_19[10]),
    .sum(sum_19[10]));
  AL_FADD comp19_11 (
    .a(i19[11]),
    .b(sum_18[11]),
    .c(cout_19[10]),
    .cout(cout_19[11]),
    .sum(sum_19[11]));
  AL_FADD comp19_12 (
    .a(i19[12]),
    .b(sum_18[12]),
    .c(cout_19[11]),
    .cout(cout_19[12]),
    .sum(sum_19[12]));
  AL_FADD comp19_13 (
    .a(i19[13]),
    .b(sum_18[13]),
    .c(cout_19[12]),
    .cout(cout_19[13]),
    .sum(sum_19[13]));
  AL_FADD comp19_14 (
    .a(i19[14]),
    .b(sum_18[14]),
    .c(cout_19[13]),
    .cout(cout_19[14]),
    .sum(sum_19[14]));
  AL_FADD comp19_15 (
    .a(i19[15]),
    .b(sum_18[15]),
    .c(cout_19[14]),
    .cout(cout_19[15]),
    .sum(sum_19[15]));
  AL_FADD comp19_16 (
    .a(i19[16]),
    .b(sum_18[16]),
    .c(cout_19[15]),
    .cout(cout_19[16]),
    .sum(sum_19[16]));
  AL_FADD comp19_17 (
    .a(i19[17]),
    .b(sum_18[17]),
    .c(cout_19[16]),
    .cout(cout_19[17]),
    .sum(sum_19[17]));
  AL_FADD comp19_18 (
    .a(i19[18]),
    .b(sum_18[18]),
    .c(cout_19[17]),
    .cout(cout_19[18]),
    .sum(sum_19[18]));
  AL_FADD comp19_19 (
    .a(i19[19]),
    .b(sum_18[19]),
    .c(cout_19[18]),
    .cout(cout_19[19]),
    .sum(sum_19[19]));
  AL_FADD comp19_2 (
    .a(i19[2]),
    .b(sum_18[2]),
    .c(cout_19[1]),
    .cout(cout_19[2]),
    .sum(sum_19[2]));
  AL_FADD comp19_20 (
    .a(i19[20]),
    .b(sum_18[20]),
    .c(cout_19[19]),
    .cout(cout_19[20]),
    .sum(sum_19[20]));
  AL_FADD comp19_21 (
    .a(i19[21]),
    .b(sum_18[21]),
    .c(cout_19[20]),
    .cout(cout_19[21]),
    .sum(sum_19[21]));
  AL_FADD comp19_22 (
    .a(i19[22]),
    .b(sum_18[22]),
    .c(cout_19[21]),
    .cout(cout_19[22]),
    .sum(sum_19[22]));
  AL_FADD comp19_23 (
    .a(i19[23]),
    .b(sum_18[23]),
    .c(cout_19[22]),
    .cout(cout_19[23]),
    .sum(sum_19[23]));
  AL_FADD comp19_24 (
    .a(i19[24]),
    .b(sum_18[24]),
    .c(cout_19[23]),
    .cout(cout_19[24]),
    .sum(sum_19[24]));
  AL_FADD comp19_25 (
    .a(i19[25]),
    .b(sum_18[25]),
    .c(cout_19[24]),
    .cout(cout_19[25]),
    .sum(sum_19[25]));
  AL_FADD comp19_26 (
    .a(i19[26]),
    .b(sum_18[26]),
    .c(cout_19[25]),
    .cout(cout_19[26]),
    .sum(sum_19[26]));
  AL_FADD comp19_27 (
    .a(i19[27]),
    .b(sum_18[27]),
    .c(cout_19[26]),
    .cout(cout_19[27]),
    .sum(sum_19[27]));
  AL_FADD comp19_28 (
    .a(1'b0),
    .b(sum_18[28]),
    .c(cout_19[27]),
    .cout(cout_19[28]),
    .sum(sum_19[28]));
  AL_FADD comp19_29 (
    .a(1'b0),
    .b(sum_18[29]),
    .c(cout_19[28]),
    .cout(cout_19[29]),
    .sum(sum_19[29]));
  AL_FADD comp19_3 (
    .a(i19[3]),
    .b(sum_18[3]),
    .c(cout_19[2]),
    .cout(cout_19[3]),
    .sum(sum_19[3]));
  AL_FADD comp19_30 (
    .a(1'b0),
    .b(sum_18[30]),
    .c(cout_19[29]),
    .cout(cout_19[30]),
    .sum(sum_19[30]));
  AL_FADD comp19_31 (
    .a(1'b0),
    .b(sum_18[31]),
    .c(cout_19[30]),
    .cout(cout_19[31]),
    .sum(sum_19[31]));
  AL_FADD comp19_32 (
    .a(1'b0),
    .b(sum_18[32]),
    .c(cout_19[31]),
    .cout(cout_19[32]),
    .sum(sum_19[32]));
  AL_FADD comp19_33 (
    .a(1'b0),
    .b(sum_18[33]),
    .c(cout_19[32]),
    .cout(cout_19[33]),
    .sum(sum_19[33]));
  AL_FADD comp19_34 (
    .a(1'b0),
    .b(sum_18[34]),
    .c(cout_19[33]),
    .cout(cout_19[34]),
    .sum(sum_19[34]));
  AL_FADD comp19_35 (
    .a(1'b0),
    .b(sum_18[35]),
    .c(cout_19[34]),
    .cout(cout_19[35]),
    .sum(sum_19[35]));
  AL_FADD comp19_36 (
    .a(1'b0),
    .b(sum_18[36]),
    .c(cout_19[35]),
    .cout(cout_19[36]),
    .sum(sum_19[36]));
  AL_FADD comp19_37 (
    .a(1'b0),
    .b(sum_18[37]),
    .c(cout_19[36]),
    .cout(cout_19[37]),
    .sum(sum_19[37]));
  AL_FADD comp19_38 (
    .a(1'b0),
    .b(sum_18[38]),
    .c(cout_19[37]),
    .cout(cout_19[38]),
    .sum(sum_19[38]));
  AL_FADD comp19_39 (
    .a(1'b0),
    .b(sum_18[39]),
    .c(cout_19[38]),
    .cout(cout_19[39]),
    .sum(sum_19[39]));
  AL_FADD comp19_4 (
    .a(i19[4]),
    .b(sum_18[4]),
    .c(cout_19[3]),
    .cout(cout_19[4]),
    .sum(sum_19[4]));
  AL_FADD comp19_40 (
    .a(1'b0),
    .b(sum_18[40]),
    .c(cout_19[39]),
    .cout(cout_19[40]),
    .sum(sum_19[40]));
  AL_FADD comp19_41 (
    .a(1'b0),
    .b(sum_18[41]),
    .c(cout_19[40]),
    .cout(cout_19[41]),
    .sum(sum_19[41]));
  AL_FADD comp19_42 (
    .a(1'b0),
    .b(sum_18[42]),
    .c(cout_19[41]),
    .cout(cout_19[42]),
    .sum(sum_19[42]));
  AL_FADD comp19_43 (
    .a(1'b0),
    .b(sum_18[43]),
    .c(cout_19[42]),
    .cout(cout_19[43]),
    .sum(sum_19[43]));
  AL_FADD comp19_44 (
    .a(1'b0),
    .b(sum_18[44]),
    .c(cout_19[43]),
    .cout(cout_19[44]),
    .sum(sum_19[44]));
  AL_FADD comp19_45 (
    .a(1'b0),
    .b(sum_18[45]),
    .c(cout_19[44]),
    .cout(cout_19[45]),
    .sum(sum_19[45]));
  AL_FADD comp19_46 (
    .a(1'b0),
    .b(sum_18[46]),
    .c(cout_19[45]),
    .cout(cout_19[46]),
    .sum(sum_19[46]));
  AL_FADD comp19_47 (
    .a(1'b0),
    .b(sum_18[47]),
    .c(cout_19[46]),
    .cout(cout_19[47]),
    .sum(sum_19[47]));
  AL_FADD comp19_5 (
    .a(i19[5]),
    .b(sum_18[5]),
    .c(cout_19[4]),
    .cout(cout_19[5]),
    .sum(sum_19[5]));
  AL_FADD comp19_6 (
    .a(i19[6]),
    .b(sum_18[6]),
    .c(cout_19[5]),
    .cout(cout_19[6]),
    .sum(sum_19[6]));
  AL_FADD comp19_7 (
    .a(i19[7]),
    .b(sum_18[7]),
    .c(cout_19[6]),
    .cout(cout_19[7]),
    .sum(sum_19[7]));
  AL_FADD comp19_8 (
    .a(i19[8]),
    .b(sum_18[8]),
    .c(cout_19[7]),
    .cout(cout_19[8]),
    .sum(sum_19[8]));
  AL_FADD comp19_9 (
    .a(i19[9]),
    .b(sum_18[9]),
    .c(cout_19[8]),
    .cout(cout_19[9]),
    .sum(sum_19[9]));
  AL_FADD comp1_0 (
    .a(i1[0]),
    .b(i0[0]),
    .c(1'b0),
    .cout(cout_1[0]),
    .sum(sum_1[0]));
  AL_FADD comp1_1 (
    .a(i1[1]),
    .b(i0[1]),
    .c(cout_1[0]),
    .cout(cout_1[1]),
    .sum(sum_1[1]));
  AL_FADD comp1_10 (
    .a(i1[10]),
    .b(i0[10]),
    .c(cout_1[9]),
    .cout(cout_1[10]),
    .sum(sum_1[10]));
  AL_FADD comp1_11 (
    .a(i1[11]),
    .b(i0[11]),
    .c(cout_1[10]),
    .cout(cout_1[11]),
    .sum(sum_1[11]));
  AL_FADD comp1_12 (
    .a(i1[12]),
    .b(i0[12]),
    .c(cout_1[11]),
    .cout(cout_1[12]),
    .sum(sum_1[12]));
  AL_FADD comp1_13 (
    .a(i1[13]),
    .b(i0[13]),
    .c(cout_1[12]),
    .cout(cout_1[13]),
    .sum(sum_1[13]));
  AL_FADD comp1_14 (
    .a(i1[14]),
    .b(i0[14]),
    .c(cout_1[13]),
    .cout(cout_1[14]),
    .sum(sum_1[14]));
  AL_FADD comp1_15 (
    .a(i1[15]),
    .b(i0[15]),
    .c(cout_1[14]),
    .cout(cout_1[15]),
    .sum(sum_1[15]));
  AL_FADD comp1_16 (
    .a(i1[16]),
    .b(i0[16]),
    .c(cout_1[15]),
    .cout(cout_1[16]),
    .sum(sum_1[16]));
  AL_FADD comp1_17 (
    .a(i1[17]),
    .b(i0[17]),
    .c(cout_1[16]),
    .cout(cout_1[17]),
    .sum(sum_1[17]));
  AL_FADD comp1_18 (
    .a(i1[18]),
    .b(i0[18]),
    .c(cout_1[17]),
    .cout(cout_1[18]),
    .sum(sum_1[18]));
  AL_FADD comp1_19 (
    .a(i1[19]),
    .b(i0[19]),
    .c(cout_1[18]),
    .cout(cout_1[19]),
    .sum(sum_1[19]));
  AL_FADD comp1_2 (
    .a(i1[2]),
    .b(i0[2]),
    .c(cout_1[1]),
    .cout(cout_1[2]),
    .sum(sum_1[2]));
  AL_FADD comp1_20 (
    .a(i1[20]),
    .b(i0[20]),
    .c(cout_1[19]),
    .cout(cout_1[20]),
    .sum(sum_1[20]));
  AL_FADD comp1_21 (
    .a(i1[21]),
    .b(i0[21]),
    .c(cout_1[20]),
    .cout(cout_1[21]),
    .sum(sum_1[21]));
  AL_FADD comp1_22 (
    .a(i1[22]),
    .b(i0[22]),
    .c(cout_1[21]),
    .cout(cout_1[22]),
    .sum(sum_1[22]));
  AL_FADD comp1_23 (
    .a(i1[23]),
    .b(i0[23]),
    .c(cout_1[22]),
    .cout(cout_1[23]),
    .sum(sum_1[23]));
  AL_FADD comp1_24 (
    .a(i1[24]),
    .b(i0[24]),
    .c(cout_1[23]),
    .cout(cout_1[24]),
    .sum(sum_1[24]));
  AL_FADD comp1_25 (
    .a(i1[25]),
    .b(i0[25]),
    .c(cout_1[24]),
    .cout(cout_1[25]),
    .sum(sum_1[25]));
  AL_FADD comp1_26 (
    .a(i1[26]),
    .b(i0[26]),
    .c(cout_1[25]),
    .cout(cout_1[26]),
    .sum(sum_1[26]));
  AL_FADD comp1_27 (
    .a(i1[27]),
    .b(i0[27]),
    .c(cout_1[26]),
    .cout(cout_1[27]),
    .sum(sum_1[27]));
  AL_FADD comp1_28 (
    .a(i1[28]),
    .b(i0[28]),
    .c(cout_1[27]),
    .cout(cout_1[28]),
    .sum(sum_1[28]));
  AL_FADD comp1_29 (
    .a(i1[29]),
    .b(i0[29]),
    .c(cout_1[28]),
    .cout(cout_1[29]),
    .sum(sum_1[29]));
  AL_FADD comp1_3 (
    .a(i1[3]),
    .b(i0[3]),
    .c(cout_1[2]),
    .cout(cout_1[3]),
    .sum(sum_1[3]));
  AL_FADD comp1_30 (
    .a(i1[30]),
    .b(i0[30]),
    .c(cout_1[29]),
    .cout(cout_1[30]),
    .sum(sum_1[30]));
  AL_FADD comp1_31 (
    .a(i1[31]),
    .b(i0[31]),
    .c(cout_1[30]),
    .cout(cout_1[31]),
    .sum(sum_1[31]));
  AL_FADD comp1_32 (
    .a(i1[32]),
    .b(i0[32]),
    .c(cout_1[31]),
    .cout(cout_1[32]),
    .sum(sum_1[32]));
  AL_FADD comp1_33 (
    .a(i1[33]),
    .b(i0[33]),
    .c(cout_1[32]),
    .cout(cout_1[33]),
    .sum(sum_1[33]));
  AL_FADD comp1_34 (
    .a(i1[34]),
    .b(i0[34]),
    .c(cout_1[33]),
    .cout(cout_1[34]),
    .sum(sum_1[34]));
  AL_FADD comp1_35 (
    .a(i1[35]),
    .b(i0[35]),
    .c(cout_1[34]),
    .cout(cout_1[35]),
    .sum(sum_1[35]));
  AL_FADD comp1_36 (
    .a(i1[36]),
    .b(i0[36]),
    .c(cout_1[35]),
    .cout(cout_1[36]),
    .sum(sum_1[36]));
  AL_FADD comp1_37 (
    .a(i1[37]),
    .b(i0[37]),
    .c(cout_1[36]),
    .cout(cout_1[37]),
    .sum(sum_1[37]));
  AL_FADD comp1_38 (
    .a(i1[38]),
    .b(i0[38]),
    .c(cout_1[37]),
    .cout(cout_1[38]),
    .sum(sum_1[38]));
  AL_FADD comp1_39 (
    .a(i1[39]),
    .b(i0[39]),
    .c(cout_1[38]),
    .cout(cout_1[39]),
    .sum(sum_1[39]));
  AL_FADD comp1_4 (
    .a(i1[4]),
    .b(i0[4]),
    .c(cout_1[3]),
    .cout(cout_1[4]),
    .sum(sum_1[4]));
  AL_FADD comp1_40 (
    .a(i1[40]),
    .b(i0[40]),
    .c(cout_1[39]),
    .cout(cout_1[40]),
    .sum(sum_1[40]));
  AL_FADD comp1_41 (
    .a(i1[41]),
    .b(i0[41]),
    .c(cout_1[40]),
    .cout(cout_1[41]),
    .sum(sum_1[41]));
  AL_FADD comp1_42 (
    .a(i1[42]),
    .b(i0[42]),
    .c(cout_1[41]),
    .cout(cout_1[42]),
    .sum(sum_1[42]));
  AL_FADD comp1_43 (
    .a(i1[43]),
    .b(i0[43]),
    .c(cout_1[42]),
    .cout(cout_1[43]),
    .sum(sum_1[43]));
  AL_FADD comp1_44 (
    .a(i1[44]),
    .b(i0[44]),
    .c(cout_1[43]),
    .cout(cout_1[44]),
    .sum(sum_1[44]));
  AL_FADD comp1_45 (
    .a(i1[45]),
    .b(i0[45]),
    .c(cout_1[44]),
    .cout(cout_1[45]),
    .sum(sum_1[45]));
  AL_FADD comp1_46 (
    .a(1'b0),
    .b(i0[46]),
    .c(cout_1[45]),
    .cout(cout_1[46]),
    .sum(sum_1[46]));
  AL_FADD comp1_5 (
    .a(i1[5]),
    .b(i0[5]),
    .c(cout_1[4]),
    .cout(cout_1[5]),
    .sum(sum_1[5]));
  AL_FADD comp1_6 (
    .a(i1[6]),
    .b(i0[6]),
    .c(cout_1[5]),
    .cout(cout_1[6]),
    .sum(sum_1[6]));
  AL_FADD comp1_7 (
    .a(i1[7]),
    .b(i0[7]),
    .c(cout_1[6]),
    .cout(cout_1[7]),
    .sum(sum_1[7]));
  AL_FADD comp1_8 (
    .a(i1[8]),
    .b(i0[8]),
    .c(cout_1[7]),
    .cout(cout_1[8]),
    .sum(sum_1[8]));
  AL_FADD comp1_9 (
    .a(i1[9]),
    .b(i0[9]),
    .c(cout_1[8]),
    .cout(cout_1[9]),
    .sum(sum_1[9]));
  AL_FADD comp20_0 (
    .a(i20[0]),
    .b(sum_19[0]),
    .c(1'b0),
    .cout(cout_20[0]),
    .sum(sum_20[0]));
  AL_FADD comp20_1 (
    .a(i20[1]),
    .b(sum_19[1]),
    .c(cout_20[0]),
    .cout(cout_20[1]),
    .sum(sum_20[1]));
  AL_FADD comp20_10 (
    .a(i20[10]),
    .b(sum_19[10]),
    .c(cout_20[9]),
    .cout(cout_20[10]),
    .sum(sum_20[10]));
  AL_FADD comp20_11 (
    .a(i20[11]),
    .b(sum_19[11]),
    .c(cout_20[10]),
    .cout(cout_20[11]),
    .sum(sum_20[11]));
  AL_FADD comp20_12 (
    .a(i20[12]),
    .b(sum_19[12]),
    .c(cout_20[11]),
    .cout(cout_20[12]),
    .sum(sum_20[12]));
  AL_FADD comp20_13 (
    .a(i20[13]),
    .b(sum_19[13]),
    .c(cout_20[12]),
    .cout(cout_20[13]),
    .sum(sum_20[13]));
  AL_FADD comp20_14 (
    .a(i20[14]),
    .b(sum_19[14]),
    .c(cout_20[13]),
    .cout(cout_20[14]),
    .sum(sum_20[14]));
  AL_FADD comp20_15 (
    .a(i20[15]),
    .b(sum_19[15]),
    .c(cout_20[14]),
    .cout(cout_20[15]),
    .sum(sum_20[15]));
  AL_FADD comp20_16 (
    .a(i20[16]),
    .b(sum_19[16]),
    .c(cout_20[15]),
    .cout(cout_20[16]),
    .sum(sum_20[16]));
  AL_FADD comp20_17 (
    .a(i20[17]),
    .b(sum_19[17]),
    .c(cout_20[16]),
    .cout(cout_20[17]),
    .sum(sum_20[17]));
  AL_FADD comp20_18 (
    .a(i20[18]),
    .b(sum_19[18]),
    .c(cout_20[17]),
    .cout(cout_20[18]),
    .sum(sum_20[18]));
  AL_FADD comp20_19 (
    .a(i20[19]),
    .b(sum_19[19]),
    .c(cout_20[18]),
    .cout(cout_20[19]),
    .sum(sum_20[19]));
  AL_FADD comp20_2 (
    .a(i20[2]),
    .b(sum_19[2]),
    .c(cout_20[1]),
    .cout(cout_20[2]),
    .sum(sum_20[2]));
  AL_FADD comp20_20 (
    .a(i20[20]),
    .b(sum_19[20]),
    .c(cout_20[19]),
    .cout(cout_20[20]),
    .sum(sum_20[20]));
  AL_FADD comp20_21 (
    .a(i20[21]),
    .b(sum_19[21]),
    .c(cout_20[20]),
    .cout(cout_20[21]),
    .sum(sum_20[21]));
  AL_FADD comp20_22 (
    .a(i20[22]),
    .b(sum_19[22]),
    .c(cout_20[21]),
    .cout(cout_20[22]),
    .sum(sum_20[22]));
  AL_FADD comp20_23 (
    .a(i20[23]),
    .b(sum_19[23]),
    .c(cout_20[22]),
    .cout(cout_20[23]),
    .sum(sum_20[23]));
  AL_FADD comp20_24 (
    .a(i20[24]),
    .b(sum_19[24]),
    .c(cout_20[23]),
    .cout(cout_20[24]),
    .sum(sum_20[24]));
  AL_FADD comp20_25 (
    .a(i20[25]),
    .b(sum_19[25]),
    .c(cout_20[24]),
    .cout(cout_20[25]),
    .sum(sum_20[25]));
  AL_FADD comp20_26 (
    .a(i20[26]),
    .b(sum_19[26]),
    .c(cout_20[25]),
    .cout(cout_20[26]),
    .sum(sum_20[26]));
  AL_FADD comp20_27 (
    .a(1'b0),
    .b(sum_19[27]),
    .c(cout_20[26]),
    .cout(cout_20[27]),
    .sum(sum_20[27]));
  AL_FADD comp20_28 (
    .a(1'b0),
    .b(sum_19[28]),
    .c(cout_20[27]),
    .cout(cout_20[28]),
    .sum(sum_20[28]));
  AL_FADD comp20_29 (
    .a(1'b0),
    .b(sum_19[29]),
    .c(cout_20[28]),
    .cout(cout_20[29]),
    .sum(sum_20[29]));
  AL_FADD comp20_3 (
    .a(i20[3]),
    .b(sum_19[3]),
    .c(cout_20[2]),
    .cout(cout_20[3]),
    .sum(sum_20[3]));
  AL_FADD comp20_30 (
    .a(1'b0),
    .b(sum_19[30]),
    .c(cout_20[29]),
    .cout(cout_20[30]),
    .sum(sum_20[30]));
  AL_FADD comp20_31 (
    .a(1'b0),
    .b(sum_19[31]),
    .c(cout_20[30]),
    .cout(cout_20[31]),
    .sum(sum_20[31]));
  AL_FADD comp20_32 (
    .a(1'b0),
    .b(sum_19[32]),
    .c(cout_20[31]),
    .cout(cout_20[32]),
    .sum(sum_20[32]));
  AL_FADD comp20_33 (
    .a(1'b0),
    .b(sum_19[33]),
    .c(cout_20[32]),
    .cout(cout_20[33]),
    .sum(sum_20[33]));
  AL_FADD comp20_34 (
    .a(1'b0),
    .b(sum_19[34]),
    .c(cout_20[33]),
    .cout(cout_20[34]),
    .sum(sum_20[34]));
  AL_FADD comp20_35 (
    .a(1'b0),
    .b(sum_19[35]),
    .c(cout_20[34]),
    .cout(cout_20[35]),
    .sum(sum_20[35]));
  AL_FADD comp20_36 (
    .a(1'b0),
    .b(sum_19[36]),
    .c(cout_20[35]),
    .cout(cout_20[36]),
    .sum(sum_20[36]));
  AL_FADD comp20_37 (
    .a(1'b0),
    .b(sum_19[37]),
    .c(cout_20[36]),
    .cout(cout_20[37]),
    .sum(sum_20[37]));
  AL_FADD comp20_38 (
    .a(1'b0),
    .b(sum_19[38]),
    .c(cout_20[37]),
    .cout(cout_20[38]),
    .sum(sum_20[38]));
  AL_FADD comp20_39 (
    .a(1'b0),
    .b(sum_19[39]),
    .c(cout_20[38]),
    .cout(cout_20[39]),
    .sum(sum_20[39]));
  AL_FADD comp20_4 (
    .a(i20[4]),
    .b(sum_19[4]),
    .c(cout_20[3]),
    .cout(cout_20[4]),
    .sum(sum_20[4]));
  AL_FADD comp20_40 (
    .a(1'b0),
    .b(sum_19[40]),
    .c(cout_20[39]),
    .cout(cout_20[40]),
    .sum(sum_20[40]));
  AL_FADD comp20_41 (
    .a(1'b0),
    .b(sum_19[41]),
    .c(cout_20[40]),
    .cout(cout_20[41]),
    .sum(sum_20[41]));
  AL_FADD comp20_42 (
    .a(1'b0),
    .b(sum_19[42]),
    .c(cout_20[41]),
    .cout(cout_20[42]),
    .sum(sum_20[42]));
  AL_FADD comp20_43 (
    .a(1'b0),
    .b(sum_19[43]),
    .c(cout_20[42]),
    .cout(cout_20[43]),
    .sum(sum_20[43]));
  AL_FADD comp20_44 (
    .a(1'b0),
    .b(sum_19[44]),
    .c(cout_20[43]),
    .cout(cout_20[44]),
    .sum(sum_20[44]));
  AL_FADD comp20_45 (
    .a(1'b0),
    .b(sum_19[45]),
    .c(cout_20[44]),
    .cout(cout_20[45]),
    .sum(sum_20[45]));
  AL_FADD comp20_46 (
    .a(1'b0),
    .b(sum_19[46]),
    .c(cout_20[45]),
    .cout(cout_20[46]),
    .sum(sum_20[46]));
  AL_FADD comp20_47 (
    .a(1'b0),
    .b(sum_19[47]),
    .c(cout_20[46]),
    .cout(cout_20[47]),
    .sum(sum_20[47]));
  AL_FADD comp20_5 (
    .a(i20[5]),
    .b(sum_19[5]),
    .c(cout_20[4]),
    .cout(cout_20[5]),
    .sum(sum_20[5]));
  AL_FADD comp20_6 (
    .a(i20[6]),
    .b(sum_19[6]),
    .c(cout_20[5]),
    .cout(cout_20[6]),
    .sum(sum_20[6]));
  AL_FADD comp20_7 (
    .a(i20[7]),
    .b(sum_19[7]),
    .c(cout_20[6]),
    .cout(cout_20[7]),
    .sum(sum_20[7]));
  AL_FADD comp20_8 (
    .a(i20[8]),
    .b(sum_19[8]),
    .c(cout_20[7]),
    .cout(cout_20[8]),
    .sum(sum_20[8]));
  AL_FADD comp20_9 (
    .a(i20[9]),
    .b(sum_19[9]),
    .c(cout_20[8]),
    .cout(cout_20[9]),
    .sum(sum_20[9]));
  AL_FADD comp21_0 (
    .a(i21[0]),
    .b(sum_20[0]),
    .c(1'b0),
    .cout(cout_21[0]),
    .sum(sum_21[0]));
  AL_FADD comp21_1 (
    .a(i21[1]),
    .b(sum_20[1]),
    .c(cout_21[0]),
    .cout(cout_21[1]),
    .sum(sum_21[1]));
  AL_FADD comp21_10 (
    .a(i21[10]),
    .b(sum_20[10]),
    .c(cout_21[9]),
    .cout(cout_21[10]),
    .sum(sum_21[10]));
  AL_FADD comp21_11 (
    .a(i21[11]),
    .b(sum_20[11]),
    .c(cout_21[10]),
    .cout(cout_21[11]),
    .sum(sum_21[11]));
  AL_FADD comp21_12 (
    .a(i21[12]),
    .b(sum_20[12]),
    .c(cout_21[11]),
    .cout(cout_21[12]),
    .sum(sum_21[12]));
  AL_FADD comp21_13 (
    .a(i21[13]),
    .b(sum_20[13]),
    .c(cout_21[12]),
    .cout(cout_21[13]),
    .sum(sum_21[13]));
  AL_FADD comp21_14 (
    .a(i21[14]),
    .b(sum_20[14]),
    .c(cout_21[13]),
    .cout(cout_21[14]),
    .sum(sum_21[14]));
  AL_FADD comp21_15 (
    .a(i21[15]),
    .b(sum_20[15]),
    .c(cout_21[14]),
    .cout(cout_21[15]),
    .sum(sum_21[15]));
  AL_FADD comp21_16 (
    .a(i21[16]),
    .b(sum_20[16]),
    .c(cout_21[15]),
    .cout(cout_21[16]),
    .sum(sum_21[16]));
  AL_FADD comp21_17 (
    .a(i21[17]),
    .b(sum_20[17]),
    .c(cout_21[16]),
    .cout(cout_21[17]),
    .sum(sum_21[17]));
  AL_FADD comp21_18 (
    .a(i21[18]),
    .b(sum_20[18]),
    .c(cout_21[17]),
    .cout(cout_21[18]),
    .sum(sum_21[18]));
  AL_FADD comp21_19 (
    .a(i21[19]),
    .b(sum_20[19]),
    .c(cout_21[18]),
    .cout(cout_21[19]),
    .sum(sum_21[19]));
  AL_FADD comp21_2 (
    .a(i21[2]),
    .b(sum_20[2]),
    .c(cout_21[1]),
    .cout(cout_21[2]),
    .sum(sum_21[2]));
  AL_FADD comp21_20 (
    .a(i21[20]),
    .b(sum_20[20]),
    .c(cout_21[19]),
    .cout(cout_21[20]),
    .sum(sum_21[20]));
  AL_FADD comp21_21 (
    .a(i21[21]),
    .b(sum_20[21]),
    .c(cout_21[20]),
    .cout(cout_21[21]),
    .sum(sum_21[21]));
  AL_FADD comp21_22 (
    .a(i21[22]),
    .b(sum_20[22]),
    .c(cout_21[21]),
    .cout(cout_21[22]),
    .sum(sum_21[22]));
  AL_FADD comp21_23 (
    .a(i21[23]),
    .b(sum_20[23]),
    .c(cout_21[22]),
    .cout(cout_21[23]),
    .sum(sum_21[23]));
  AL_FADD comp21_24 (
    .a(i21[24]),
    .b(sum_20[24]),
    .c(cout_21[23]),
    .cout(cout_21[24]),
    .sum(sum_21[24]));
  AL_FADD comp21_25 (
    .a(i21[25]),
    .b(sum_20[25]),
    .c(cout_21[24]),
    .cout(cout_21[25]),
    .sum(sum_21[25]));
  AL_FADD comp21_26 (
    .a(1'b0),
    .b(sum_20[26]),
    .c(cout_21[25]),
    .cout(cout_21[26]),
    .sum(sum_21[26]));
  AL_FADD comp21_27 (
    .a(1'b0),
    .b(sum_20[27]),
    .c(cout_21[26]),
    .cout(cout_21[27]),
    .sum(sum_21[27]));
  AL_FADD comp21_28 (
    .a(1'b0),
    .b(sum_20[28]),
    .c(cout_21[27]),
    .cout(cout_21[28]),
    .sum(sum_21[28]));
  AL_FADD comp21_29 (
    .a(1'b0),
    .b(sum_20[29]),
    .c(cout_21[28]),
    .cout(cout_21[29]),
    .sum(sum_21[29]));
  AL_FADD comp21_3 (
    .a(i21[3]),
    .b(sum_20[3]),
    .c(cout_21[2]),
    .cout(cout_21[3]),
    .sum(sum_21[3]));
  AL_FADD comp21_30 (
    .a(1'b0),
    .b(sum_20[30]),
    .c(cout_21[29]),
    .cout(cout_21[30]),
    .sum(sum_21[30]));
  AL_FADD comp21_31 (
    .a(1'b0),
    .b(sum_20[31]),
    .c(cout_21[30]),
    .cout(cout_21[31]),
    .sum(sum_21[31]));
  AL_FADD comp21_32 (
    .a(1'b0),
    .b(sum_20[32]),
    .c(cout_21[31]),
    .cout(cout_21[32]),
    .sum(sum_21[32]));
  AL_FADD comp21_33 (
    .a(1'b0),
    .b(sum_20[33]),
    .c(cout_21[32]),
    .cout(cout_21[33]),
    .sum(sum_21[33]));
  AL_FADD comp21_34 (
    .a(1'b0),
    .b(sum_20[34]),
    .c(cout_21[33]),
    .cout(cout_21[34]),
    .sum(sum_21[34]));
  AL_FADD comp21_35 (
    .a(1'b0),
    .b(sum_20[35]),
    .c(cout_21[34]),
    .cout(cout_21[35]),
    .sum(sum_21[35]));
  AL_FADD comp21_36 (
    .a(1'b0),
    .b(sum_20[36]),
    .c(cout_21[35]),
    .cout(cout_21[36]),
    .sum(sum_21[36]));
  AL_FADD comp21_37 (
    .a(1'b0),
    .b(sum_20[37]),
    .c(cout_21[36]),
    .cout(cout_21[37]),
    .sum(sum_21[37]));
  AL_FADD comp21_38 (
    .a(1'b0),
    .b(sum_20[38]),
    .c(cout_21[37]),
    .cout(cout_21[38]),
    .sum(sum_21[38]));
  AL_FADD comp21_39 (
    .a(1'b0),
    .b(sum_20[39]),
    .c(cout_21[38]),
    .cout(cout_21[39]),
    .sum(sum_21[39]));
  AL_FADD comp21_4 (
    .a(i21[4]),
    .b(sum_20[4]),
    .c(cout_21[3]),
    .cout(cout_21[4]),
    .sum(sum_21[4]));
  AL_FADD comp21_40 (
    .a(1'b0),
    .b(sum_20[40]),
    .c(cout_21[39]),
    .cout(cout_21[40]),
    .sum(sum_21[40]));
  AL_FADD comp21_41 (
    .a(1'b0),
    .b(sum_20[41]),
    .c(cout_21[40]),
    .cout(cout_21[41]),
    .sum(sum_21[41]));
  AL_FADD comp21_42 (
    .a(1'b0),
    .b(sum_20[42]),
    .c(cout_21[41]),
    .cout(cout_21[42]),
    .sum(sum_21[42]));
  AL_FADD comp21_43 (
    .a(1'b0),
    .b(sum_20[43]),
    .c(cout_21[42]),
    .cout(cout_21[43]),
    .sum(sum_21[43]));
  AL_FADD comp21_44 (
    .a(1'b0),
    .b(sum_20[44]),
    .c(cout_21[43]),
    .cout(cout_21[44]),
    .sum(sum_21[44]));
  AL_FADD comp21_45 (
    .a(1'b0),
    .b(sum_20[45]),
    .c(cout_21[44]),
    .cout(cout_21[45]),
    .sum(sum_21[45]));
  AL_FADD comp21_46 (
    .a(1'b0),
    .b(sum_20[46]),
    .c(cout_21[45]),
    .cout(cout_21[46]),
    .sum(sum_21[46]));
  AL_FADD comp21_47 (
    .a(1'b0),
    .b(sum_20[47]),
    .c(cout_21[46]),
    .cout(cout_21[47]),
    .sum(sum_21[47]));
  AL_FADD comp21_5 (
    .a(i21[5]),
    .b(sum_20[5]),
    .c(cout_21[4]),
    .cout(cout_21[5]),
    .sum(sum_21[5]));
  AL_FADD comp21_6 (
    .a(i21[6]),
    .b(sum_20[6]),
    .c(cout_21[5]),
    .cout(cout_21[6]),
    .sum(sum_21[6]));
  AL_FADD comp21_7 (
    .a(i21[7]),
    .b(sum_20[7]),
    .c(cout_21[6]),
    .cout(cout_21[7]),
    .sum(sum_21[7]));
  AL_FADD comp21_8 (
    .a(i21[8]),
    .b(sum_20[8]),
    .c(cout_21[7]),
    .cout(cout_21[8]),
    .sum(sum_21[8]));
  AL_FADD comp21_9 (
    .a(i21[9]),
    .b(sum_20[9]),
    .c(cout_21[8]),
    .cout(cout_21[9]),
    .sum(sum_21[9]));
  AL_FADD comp22_0 (
    .a(i22[0]),
    .b(sum_21[0]),
    .c(1'b0),
    .cout(cout_22[0]),
    .sum(sum_22[0]));
  AL_FADD comp22_1 (
    .a(i22[1]),
    .b(sum_21[1]),
    .c(cout_22[0]),
    .cout(cout_22[1]),
    .sum(sum_22[1]));
  AL_FADD comp22_10 (
    .a(i22[10]),
    .b(sum_21[10]),
    .c(cout_22[9]),
    .cout(cout_22[10]),
    .sum(sum_22[10]));
  AL_FADD comp22_11 (
    .a(i22[11]),
    .b(sum_21[11]),
    .c(cout_22[10]),
    .cout(cout_22[11]),
    .sum(sum_22[11]));
  AL_FADD comp22_12 (
    .a(i22[12]),
    .b(sum_21[12]),
    .c(cout_22[11]),
    .cout(cout_22[12]),
    .sum(sum_22[12]));
  AL_FADD comp22_13 (
    .a(i22[13]),
    .b(sum_21[13]),
    .c(cout_22[12]),
    .cout(cout_22[13]),
    .sum(sum_22[13]));
  AL_FADD comp22_14 (
    .a(i22[14]),
    .b(sum_21[14]),
    .c(cout_22[13]),
    .cout(cout_22[14]),
    .sum(sum_22[14]));
  AL_FADD comp22_15 (
    .a(i22[15]),
    .b(sum_21[15]),
    .c(cout_22[14]),
    .cout(cout_22[15]),
    .sum(sum_22[15]));
  AL_FADD comp22_16 (
    .a(i22[16]),
    .b(sum_21[16]),
    .c(cout_22[15]),
    .cout(cout_22[16]),
    .sum(sum_22[16]));
  AL_FADD comp22_17 (
    .a(i22[17]),
    .b(sum_21[17]),
    .c(cout_22[16]),
    .cout(cout_22[17]),
    .sum(sum_22[17]));
  AL_FADD comp22_18 (
    .a(i22[18]),
    .b(sum_21[18]),
    .c(cout_22[17]),
    .cout(cout_22[18]),
    .sum(sum_22[18]));
  AL_FADD comp22_19 (
    .a(i22[19]),
    .b(sum_21[19]),
    .c(cout_22[18]),
    .cout(cout_22[19]),
    .sum(sum_22[19]));
  AL_FADD comp22_2 (
    .a(i22[2]),
    .b(sum_21[2]),
    .c(cout_22[1]),
    .cout(cout_22[2]),
    .sum(sum_22[2]));
  AL_FADD comp22_20 (
    .a(i22[20]),
    .b(sum_21[20]),
    .c(cout_22[19]),
    .cout(cout_22[20]),
    .sum(sum_22[20]));
  AL_FADD comp22_21 (
    .a(i22[21]),
    .b(sum_21[21]),
    .c(cout_22[20]),
    .cout(cout_22[21]),
    .sum(sum_22[21]));
  AL_FADD comp22_22 (
    .a(i22[22]),
    .b(sum_21[22]),
    .c(cout_22[21]),
    .cout(cout_22[22]),
    .sum(sum_22[22]));
  AL_FADD comp22_23 (
    .a(i22[23]),
    .b(sum_21[23]),
    .c(cout_22[22]),
    .cout(cout_22[23]),
    .sum(sum_22[23]));
  AL_FADD comp22_24 (
    .a(i22[24]),
    .b(sum_21[24]),
    .c(cout_22[23]),
    .cout(cout_22[24]),
    .sum(sum_22[24]));
  AL_FADD comp22_25 (
    .a(1'b0),
    .b(sum_21[25]),
    .c(cout_22[24]),
    .cout(cout_22[25]),
    .sum(sum_22[25]));
  AL_FADD comp22_26 (
    .a(1'b0),
    .b(sum_21[26]),
    .c(cout_22[25]),
    .cout(cout_22[26]),
    .sum(sum_22[26]));
  AL_FADD comp22_27 (
    .a(1'b0),
    .b(sum_21[27]),
    .c(cout_22[26]),
    .cout(cout_22[27]),
    .sum(sum_22[27]));
  AL_FADD comp22_28 (
    .a(1'b0),
    .b(sum_21[28]),
    .c(cout_22[27]),
    .cout(cout_22[28]),
    .sum(sum_22[28]));
  AL_FADD comp22_29 (
    .a(1'b0),
    .b(sum_21[29]),
    .c(cout_22[28]),
    .cout(cout_22[29]),
    .sum(sum_22[29]));
  AL_FADD comp22_3 (
    .a(i22[3]),
    .b(sum_21[3]),
    .c(cout_22[2]),
    .cout(cout_22[3]),
    .sum(sum_22[3]));
  AL_FADD comp22_30 (
    .a(1'b0),
    .b(sum_21[30]),
    .c(cout_22[29]),
    .cout(cout_22[30]),
    .sum(sum_22[30]));
  AL_FADD comp22_31 (
    .a(1'b0),
    .b(sum_21[31]),
    .c(cout_22[30]),
    .cout(cout_22[31]),
    .sum(sum_22[31]));
  AL_FADD comp22_32 (
    .a(1'b0),
    .b(sum_21[32]),
    .c(cout_22[31]),
    .cout(cout_22[32]),
    .sum(sum_22[32]));
  AL_FADD comp22_33 (
    .a(1'b0),
    .b(sum_21[33]),
    .c(cout_22[32]),
    .cout(cout_22[33]),
    .sum(sum_22[33]));
  AL_FADD comp22_34 (
    .a(1'b0),
    .b(sum_21[34]),
    .c(cout_22[33]),
    .cout(cout_22[34]),
    .sum(sum_22[34]));
  AL_FADD comp22_35 (
    .a(1'b0),
    .b(sum_21[35]),
    .c(cout_22[34]),
    .cout(cout_22[35]),
    .sum(sum_22[35]));
  AL_FADD comp22_36 (
    .a(1'b0),
    .b(sum_21[36]),
    .c(cout_22[35]),
    .cout(cout_22[36]),
    .sum(sum_22[36]));
  AL_FADD comp22_37 (
    .a(1'b0),
    .b(sum_21[37]),
    .c(cout_22[36]),
    .cout(cout_22[37]),
    .sum(sum_22[37]));
  AL_FADD comp22_38 (
    .a(1'b0),
    .b(sum_21[38]),
    .c(cout_22[37]),
    .cout(cout_22[38]),
    .sum(sum_22[38]));
  AL_FADD comp22_39 (
    .a(1'b0),
    .b(sum_21[39]),
    .c(cout_22[38]),
    .cout(cout_22[39]),
    .sum(sum_22[39]));
  AL_FADD comp22_4 (
    .a(i22[4]),
    .b(sum_21[4]),
    .c(cout_22[3]),
    .cout(cout_22[4]),
    .sum(sum_22[4]));
  AL_FADD comp22_40 (
    .a(1'b0),
    .b(sum_21[40]),
    .c(cout_22[39]),
    .cout(cout_22[40]),
    .sum(sum_22[40]));
  AL_FADD comp22_41 (
    .a(1'b0),
    .b(sum_21[41]),
    .c(cout_22[40]),
    .cout(cout_22[41]),
    .sum(sum_22[41]));
  AL_FADD comp22_42 (
    .a(1'b0),
    .b(sum_21[42]),
    .c(cout_22[41]),
    .cout(cout_22[42]),
    .sum(sum_22[42]));
  AL_FADD comp22_43 (
    .a(1'b0),
    .b(sum_21[43]),
    .c(cout_22[42]),
    .cout(cout_22[43]),
    .sum(sum_22[43]));
  AL_FADD comp22_44 (
    .a(1'b0),
    .b(sum_21[44]),
    .c(cout_22[43]),
    .cout(cout_22[44]),
    .sum(sum_22[44]));
  AL_FADD comp22_45 (
    .a(1'b0),
    .b(sum_21[45]),
    .c(cout_22[44]),
    .cout(cout_22[45]),
    .sum(sum_22[45]));
  AL_FADD comp22_46 (
    .a(1'b0),
    .b(sum_21[46]),
    .c(cout_22[45]),
    .cout(cout_22[46]),
    .sum(sum_22[46]));
  AL_FADD comp22_47 (
    .a(1'b0),
    .b(sum_21[47]),
    .c(cout_22[46]),
    .cout(cout_22[47]),
    .sum(sum_22[47]));
  AL_FADD comp22_5 (
    .a(i22[5]),
    .b(sum_21[5]),
    .c(cout_22[4]),
    .cout(cout_22[5]),
    .sum(sum_22[5]));
  AL_FADD comp22_6 (
    .a(i22[6]),
    .b(sum_21[6]),
    .c(cout_22[5]),
    .cout(cout_22[6]),
    .sum(sum_22[6]));
  AL_FADD comp22_7 (
    .a(i22[7]),
    .b(sum_21[7]),
    .c(cout_22[6]),
    .cout(cout_22[7]),
    .sum(sum_22[7]));
  AL_FADD comp22_8 (
    .a(i22[8]),
    .b(sum_21[8]),
    .c(cout_22[7]),
    .cout(cout_22[8]),
    .sum(sum_22[8]));
  AL_FADD comp22_9 (
    .a(i22[9]),
    .b(sum_21[9]),
    .c(cout_22[8]),
    .cout(cout_22[9]),
    .sum(sum_22[9]));
  AL_FADD comp23_0 (
    .a(i23[0]),
    .b(sum_22[0]),
    .c(1'b0),
    .cout(cout_23[0]),
    .sum(sum_23[0]));
  AL_FADD comp23_1 (
    .a(i23[1]),
    .b(sum_22[1]),
    .c(cout_23[0]),
    .cout(cout_23[1]),
    .sum(sum_23[1]));
  AL_FADD comp23_10 (
    .a(i23[10]),
    .b(sum_22[10]),
    .c(cout_23[9]),
    .cout(cout_23[10]),
    .sum(sum_23[10]));
  AL_FADD comp23_11 (
    .a(i23[11]),
    .b(sum_22[11]),
    .c(cout_23[10]),
    .cout(cout_23[11]),
    .sum(sum_23[11]));
  AL_FADD comp23_12 (
    .a(i23[12]),
    .b(sum_22[12]),
    .c(cout_23[11]),
    .cout(cout_23[12]),
    .sum(sum_23[12]));
  AL_FADD comp23_13 (
    .a(i23[13]),
    .b(sum_22[13]),
    .c(cout_23[12]),
    .cout(cout_23[13]),
    .sum(sum_23[13]));
  AL_FADD comp23_14 (
    .a(i23[14]),
    .b(sum_22[14]),
    .c(cout_23[13]),
    .cout(cout_23[14]),
    .sum(sum_23[14]));
  AL_FADD comp23_15 (
    .a(i23[15]),
    .b(sum_22[15]),
    .c(cout_23[14]),
    .cout(cout_23[15]),
    .sum(sum_23[15]));
  AL_FADD comp23_16 (
    .a(i23[16]),
    .b(sum_22[16]),
    .c(cout_23[15]),
    .cout(cout_23[16]),
    .sum(sum_23[16]));
  AL_FADD comp23_17 (
    .a(i23[17]),
    .b(sum_22[17]),
    .c(cout_23[16]),
    .cout(cout_23[17]),
    .sum(sum_23[17]));
  AL_FADD comp23_18 (
    .a(i23[18]),
    .b(sum_22[18]),
    .c(cout_23[17]),
    .cout(cout_23[18]),
    .sum(sum_23[18]));
  AL_FADD comp23_19 (
    .a(i23[19]),
    .b(sum_22[19]),
    .c(cout_23[18]),
    .cout(cout_23[19]),
    .sum(sum_23[19]));
  AL_FADD comp23_2 (
    .a(i23[2]),
    .b(sum_22[2]),
    .c(cout_23[1]),
    .cout(cout_23[2]),
    .sum(sum_23[2]));
  AL_FADD comp23_20 (
    .a(i23[20]),
    .b(sum_22[20]),
    .c(cout_23[19]),
    .cout(cout_23[20]),
    .sum(sum_23[20]));
  AL_FADD comp23_21 (
    .a(i23[21]),
    .b(sum_22[21]),
    .c(cout_23[20]),
    .cout(cout_23[21]),
    .sum(sum_23[21]));
  AL_FADD comp23_22 (
    .a(i23[22]),
    .b(sum_22[22]),
    .c(cout_23[21]),
    .cout(cout_23[22]),
    .sum(sum_23[22]));
  AL_FADD comp23_23 (
    .a(i23[23]),
    .b(sum_22[23]),
    .c(cout_23[22]),
    .cout(cout_23[23]),
    .sum(sum_23[23]));
  AL_FADD comp23_24 (
    .a(1'b0),
    .b(sum_22[24]),
    .c(cout_23[23]),
    .cout(cout_23[24]),
    .sum(sum_23[24]));
  AL_FADD comp23_25 (
    .a(1'b0),
    .b(sum_22[25]),
    .c(cout_23[24]),
    .cout(cout_23[25]),
    .sum(sum_23[25]));
  AL_FADD comp23_26 (
    .a(1'b0),
    .b(sum_22[26]),
    .c(cout_23[25]),
    .cout(cout_23[26]),
    .sum(sum_23[26]));
  AL_FADD comp23_27 (
    .a(1'b0),
    .b(sum_22[27]),
    .c(cout_23[26]),
    .cout(cout_23[27]),
    .sum(sum_23[27]));
  AL_FADD comp23_28 (
    .a(1'b0),
    .b(sum_22[28]),
    .c(cout_23[27]),
    .cout(cout_23[28]),
    .sum(sum_23[28]));
  AL_FADD comp23_29 (
    .a(1'b0),
    .b(sum_22[29]),
    .c(cout_23[28]),
    .cout(cout_23[29]),
    .sum(sum_23[29]));
  AL_FADD comp23_3 (
    .a(i23[3]),
    .b(sum_22[3]),
    .c(cout_23[2]),
    .cout(cout_23[3]),
    .sum(sum_23[3]));
  AL_FADD comp23_30 (
    .a(1'b0),
    .b(sum_22[30]),
    .c(cout_23[29]),
    .cout(cout_23[30]),
    .sum(sum_23[30]));
  AL_FADD comp23_31 (
    .a(1'b0),
    .b(sum_22[31]),
    .c(cout_23[30]),
    .cout(cout_23[31]),
    .sum(sum_23[31]));
  AL_FADD comp23_32 (
    .a(1'b0),
    .b(sum_22[32]),
    .c(cout_23[31]),
    .cout(cout_23[32]),
    .sum(sum_23[32]));
  AL_FADD comp23_33 (
    .a(1'b0),
    .b(sum_22[33]),
    .c(cout_23[32]),
    .cout(cout_23[33]),
    .sum(sum_23[33]));
  AL_FADD comp23_34 (
    .a(1'b0),
    .b(sum_22[34]),
    .c(cout_23[33]),
    .cout(cout_23[34]),
    .sum(sum_23[34]));
  AL_FADD comp23_35 (
    .a(1'b0),
    .b(sum_22[35]),
    .c(cout_23[34]),
    .cout(cout_23[35]),
    .sum(sum_23[35]));
  AL_FADD comp23_36 (
    .a(1'b0),
    .b(sum_22[36]),
    .c(cout_23[35]),
    .cout(cout_23[36]),
    .sum(sum_23[36]));
  AL_FADD comp23_37 (
    .a(1'b0),
    .b(sum_22[37]),
    .c(cout_23[36]),
    .cout(cout_23[37]),
    .sum(sum_23[37]));
  AL_FADD comp23_38 (
    .a(1'b0),
    .b(sum_22[38]),
    .c(cout_23[37]),
    .cout(cout_23[38]),
    .sum(sum_23[38]));
  AL_FADD comp23_39 (
    .a(1'b0),
    .b(sum_22[39]),
    .c(cout_23[38]),
    .cout(cout_23[39]),
    .sum(sum_23[39]));
  AL_FADD comp23_4 (
    .a(i23[4]),
    .b(sum_22[4]),
    .c(cout_23[3]),
    .cout(cout_23[4]),
    .sum(sum_23[4]));
  AL_FADD comp23_40 (
    .a(1'b0),
    .b(sum_22[40]),
    .c(cout_23[39]),
    .cout(cout_23[40]),
    .sum(sum_23[40]));
  AL_FADD comp23_41 (
    .a(1'b0),
    .b(sum_22[41]),
    .c(cout_23[40]),
    .cout(cout_23[41]),
    .sum(sum_23[41]));
  AL_FADD comp23_42 (
    .a(1'b0),
    .b(sum_22[42]),
    .c(cout_23[41]),
    .cout(cout_23[42]),
    .sum(sum_23[42]));
  AL_FADD comp23_43 (
    .a(1'b0),
    .b(sum_22[43]),
    .c(cout_23[42]),
    .cout(cout_23[43]),
    .sum(sum_23[43]));
  AL_FADD comp23_44 (
    .a(1'b0),
    .b(sum_22[44]),
    .c(cout_23[43]),
    .cout(cout_23[44]),
    .sum(sum_23[44]));
  AL_FADD comp23_45 (
    .a(1'b0),
    .b(sum_22[45]),
    .c(cout_23[44]),
    .cout(cout_23[45]),
    .sum(sum_23[45]));
  AL_FADD comp23_46 (
    .a(1'b0),
    .b(sum_22[46]),
    .c(cout_23[45]),
    .cout(cout_23[46]),
    .sum(sum_23[46]));
  AL_FADD comp23_47 (
    .a(1'b0),
    .b(sum_22[47]),
    .c(cout_23[46]),
    .cout(cout_23[47]),
    .sum(sum_23[47]));
  AL_FADD comp23_5 (
    .a(i23[5]),
    .b(sum_22[5]),
    .c(cout_23[4]),
    .cout(cout_23[5]),
    .sum(sum_23[5]));
  AL_FADD comp23_6 (
    .a(i23[6]),
    .b(sum_22[6]),
    .c(cout_23[5]),
    .cout(cout_23[6]),
    .sum(sum_23[6]));
  AL_FADD comp23_7 (
    .a(i23[7]),
    .b(sum_22[7]),
    .c(cout_23[6]),
    .cout(cout_23[7]),
    .sum(sum_23[7]));
  AL_FADD comp23_8 (
    .a(i23[8]),
    .b(sum_22[8]),
    .c(cout_23[7]),
    .cout(cout_23[8]),
    .sum(sum_23[8]));
  AL_FADD comp23_9 (
    .a(i23[9]),
    .b(sum_22[9]),
    .c(cout_23[8]),
    .cout(cout_23[9]),
    .sum(sum_23[9]));
  AL_FADD comp2_0 (
    .a(i2[0]),
    .b(sum_1[0]),
    .c(1'b0),
    .cout(cout_2[0]),
    .sum(sum_2[0]));
  AL_FADD comp2_1 (
    .a(i2[1]),
    .b(sum_1[1]),
    .c(cout_2[0]),
    .cout(cout_2[1]),
    .sum(sum_2[1]));
  AL_FADD comp2_10 (
    .a(i2[10]),
    .b(sum_1[10]),
    .c(cout_2[9]),
    .cout(cout_2[10]),
    .sum(sum_2[10]));
  AL_FADD comp2_11 (
    .a(i2[11]),
    .b(sum_1[11]),
    .c(cout_2[10]),
    .cout(cout_2[11]),
    .sum(sum_2[11]));
  AL_FADD comp2_12 (
    .a(i2[12]),
    .b(sum_1[12]),
    .c(cout_2[11]),
    .cout(cout_2[12]),
    .sum(sum_2[12]));
  AL_FADD comp2_13 (
    .a(i2[13]),
    .b(sum_1[13]),
    .c(cout_2[12]),
    .cout(cout_2[13]),
    .sum(sum_2[13]));
  AL_FADD comp2_14 (
    .a(i2[14]),
    .b(sum_1[14]),
    .c(cout_2[13]),
    .cout(cout_2[14]),
    .sum(sum_2[14]));
  AL_FADD comp2_15 (
    .a(i2[15]),
    .b(sum_1[15]),
    .c(cout_2[14]),
    .cout(cout_2[15]),
    .sum(sum_2[15]));
  AL_FADD comp2_16 (
    .a(i2[16]),
    .b(sum_1[16]),
    .c(cout_2[15]),
    .cout(cout_2[16]),
    .sum(sum_2[16]));
  AL_FADD comp2_17 (
    .a(i2[17]),
    .b(sum_1[17]),
    .c(cout_2[16]),
    .cout(cout_2[17]),
    .sum(sum_2[17]));
  AL_FADD comp2_18 (
    .a(i2[18]),
    .b(sum_1[18]),
    .c(cout_2[17]),
    .cout(cout_2[18]),
    .sum(sum_2[18]));
  AL_FADD comp2_19 (
    .a(i2[19]),
    .b(sum_1[19]),
    .c(cout_2[18]),
    .cout(cout_2[19]),
    .sum(sum_2[19]));
  AL_FADD comp2_2 (
    .a(i2[2]),
    .b(sum_1[2]),
    .c(cout_2[1]),
    .cout(cout_2[2]),
    .sum(sum_2[2]));
  AL_FADD comp2_20 (
    .a(i2[20]),
    .b(sum_1[20]),
    .c(cout_2[19]),
    .cout(cout_2[20]),
    .sum(sum_2[20]));
  AL_FADD comp2_21 (
    .a(i2[21]),
    .b(sum_1[21]),
    .c(cout_2[20]),
    .cout(cout_2[21]),
    .sum(sum_2[21]));
  AL_FADD comp2_22 (
    .a(i2[22]),
    .b(sum_1[22]),
    .c(cout_2[21]),
    .cout(cout_2[22]),
    .sum(sum_2[22]));
  AL_FADD comp2_23 (
    .a(i2[23]),
    .b(sum_1[23]),
    .c(cout_2[22]),
    .cout(cout_2[23]),
    .sum(sum_2[23]));
  AL_FADD comp2_24 (
    .a(i2[24]),
    .b(sum_1[24]),
    .c(cout_2[23]),
    .cout(cout_2[24]),
    .sum(sum_2[24]));
  AL_FADD comp2_25 (
    .a(i2[25]),
    .b(sum_1[25]),
    .c(cout_2[24]),
    .cout(cout_2[25]),
    .sum(sum_2[25]));
  AL_FADD comp2_26 (
    .a(i2[26]),
    .b(sum_1[26]),
    .c(cout_2[25]),
    .cout(cout_2[26]),
    .sum(sum_2[26]));
  AL_FADD comp2_27 (
    .a(i2[27]),
    .b(sum_1[27]),
    .c(cout_2[26]),
    .cout(cout_2[27]),
    .sum(sum_2[27]));
  AL_FADD comp2_28 (
    .a(i2[28]),
    .b(sum_1[28]),
    .c(cout_2[27]),
    .cout(cout_2[28]),
    .sum(sum_2[28]));
  AL_FADD comp2_29 (
    .a(i2[29]),
    .b(sum_1[29]),
    .c(cout_2[28]),
    .cout(cout_2[29]),
    .sum(sum_2[29]));
  AL_FADD comp2_3 (
    .a(i2[3]),
    .b(sum_1[3]),
    .c(cout_2[2]),
    .cout(cout_2[3]),
    .sum(sum_2[3]));
  AL_FADD comp2_30 (
    .a(i2[30]),
    .b(sum_1[30]),
    .c(cout_2[29]),
    .cout(cout_2[30]),
    .sum(sum_2[30]));
  AL_FADD comp2_31 (
    .a(i2[31]),
    .b(sum_1[31]),
    .c(cout_2[30]),
    .cout(cout_2[31]),
    .sum(sum_2[31]));
  AL_FADD comp2_32 (
    .a(i2[32]),
    .b(sum_1[32]),
    .c(cout_2[31]),
    .cout(cout_2[32]),
    .sum(sum_2[32]));
  AL_FADD comp2_33 (
    .a(i2[33]),
    .b(sum_1[33]),
    .c(cout_2[32]),
    .cout(cout_2[33]),
    .sum(sum_2[33]));
  AL_FADD comp2_34 (
    .a(i2[34]),
    .b(sum_1[34]),
    .c(cout_2[33]),
    .cout(cout_2[34]),
    .sum(sum_2[34]));
  AL_FADD comp2_35 (
    .a(i2[35]),
    .b(sum_1[35]),
    .c(cout_2[34]),
    .cout(cout_2[35]),
    .sum(sum_2[35]));
  AL_FADD comp2_36 (
    .a(i2[36]),
    .b(sum_1[36]),
    .c(cout_2[35]),
    .cout(cout_2[36]),
    .sum(sum_2[36]));
  AL_FADD comp2_37 (
    .a(i2[37]),
    .b(sum_1[37]),
    .c(cout_2[36]),
    .cout(cout_2[37]),
    .sum(sum_2[37]));
  AL_FADD comp2_38 (
    .a(i2[38]),
    .b(sum_1[38]),
    .c(cout_2[37]),
    .cout(cout_2[38]),
    .sum(sum_2[38]));
  AL_FADD comp2_39 (
    .a(i2[39]),
    .b(sum_1[39]),
    .c(cout_2[38]),
    .cout(cout_2[39]),
    .sum(sum_2[39]));
  AL_FADD comp2_4 (
    .a(i2[4]),
    .b(sum_1[4]),
    .c(cout_2[3]),
    .cout(cout_2[4]),
    .sum(sum_2[4]));
  AL_FADD comp2_40 (
    .a(i2[40]),
    .b(sum_1[40]),
    .c(cout_2[39]),
    .cout(cout_2[40]),
    .sum(sum_2[40]));
  AL_FADD comp2_41 (
    .a(i2[41]),
    .b(sum_1[41]),
    .c(cout_2[40]),
    .cout(cout_2[41]),
    .sum(sum_2[41]));
  AL_FADD comp2_42 (
    .a(i2[42]),
    .b(sum_1[42]),
    .c(cout_2[41]),
    .cout(cout_2[42]),
    .sum(sum_2[42]));
  AL_FADD comp2_43 (
    .a(i2[43]),
    .b(sum_1[43]),
    .c(cout_2[42]),
    .cout(cout_2[43]),
    .sum(sum_2[43]));
  AL_FADD comp2_44 (
    .a(i2[44]),
    .b(sum_1[44]),
    .c(cout_2[43]),
    .cout(cout_2[44]),
    .sum(sum_2[44]));
  AL_FADD comp2_45 (
    .a(1'b0),
    .b(sum_1[45]),
    .c(cout_2[44]),
    .cout(cout_2[45]),
    .sum(sum_2[45]));
  AL_FADD comp2_46 (
    .a(1'b0),
    .b(sum_1[46]),
    .c(cout_2[45]),
    .cout(cout_2[46]),
    .sum(sum_2[46]));
  AL_FADD comp2_47 (
    .a(1'b0),
    .b(cout_1[46]),
    .c(cout_2[46]),
    .cout(cout_2[47]),
    .sum(sum_2[47]));
  AL_FADD comp2_5 (
    .a(i2[5]),
    .b(sum_1[5]),
    .c(cout_2[4]),
    .cout(cout_2[5]),
    .sum(sum_2[5]));
  AL_FADD comp2_6 (
    .a(i2[6]),
    .b(sum_1[6]),
    .c(cout_2[5]),
    .cout(cout_2[6]),
    .sum(sum_2[6]));
  AL_FADD comp2_7 (
    .a(i2[7]),
    .b(sum_1[7]),
    .c(cout_2[6]),
    .cout(cout_2[7]),
    .sum(sum_2[7]));
  AL_FADD comp2_8 (
    .a(i2[8]),
    .b(sum_1[8]),
    .c(cout_2[7]),
    .cout(cout_2[8]),
    .sum(sum_2[8]));
  AL_FADD comp2_9 (
    .a(i2[9]),
    .b(sum_1[9]),
    .c(cout_2[8]),
    .cout(cout_2[9]),
    .sum(sum_2[9]));
  AL_FADD comp3_0 (
    .a(i3[0]),
    .b(sum_2[0]),
    .c(1'b0),
    .cout(cout_3[0]),
    .sum(sum_3[0]));
  AL_FADD comp3_1 (
    .a(i3[1]),
    .b(sum_2[1]),
    .c(cout_3[0]),
    .cout(cout_3[1]),
    .sum(sum_3[1]));
  AL_FADD comp3_10 (
    .a(i3[10]),
    .b(sum_2[10]),
    .c(cout_3[9]),
    .cout(cout_3[10]),
    .sum(sum_3[10]));
  AL_FADD comp3_11 (
    .a(i3[11]),
    .b(sum_2[11]),
    .c(cout_3[10]),
    .cout(cout_3[11]),
    .sum(sum_3[11]));
  AL_FADD comp3_12 (
    .a(i3[12]),
    .b(sum_2[12]),
    .c(cout_3[11]),
    .cout(cout_3[12]),
    .sum(sum_3[12]));
  AL_FADD comp3_13 (
    .a(i3[13]),
    .b(sum_2[13]),
    .c(cout_3[12]),
    .cout(cout_3[13]),
    .sum(sum_3[13]));
  AL_FADD comp3_14 (
    .a(i3[14]),
    .b(sum_2[14]),
    .c(cout_3[13]),
    .cout(cout_3[14]),
    .sum(sum_3[14]));
  AL_FADD comp3_15 (
    .a(i3[15]),
    .b(sum_2[15]),
    .c(cout_3[14]),
    .cout(cout_3[15]),
    .sum(sum_3[15]));
  AL_FADD comp3_16 (
    .a(i3[16]),
    .b(sum_2[16]),
    .c(cout_3[15]),
    .cout(cout_3[16]),
    .sum(sum_3[16]));
  AL_FADD comp3_17 (
    .a(i3[17]),
    .b(sum_2[17]),
    .c(cout_3[16]),
    .cout(cout_3[17]),
    .sum(sum_3[17]));
  AL_FADD comp3_18 (
    .a(i3[18]),
    .b(sum_2[18]),
    .c(cout_3[17]),
    .cout(cout_3[18]),
    .sum(sum_3[18]));
  AL_FADD comp3_19 (
    .a(i3[19]),
    .b(sum_2[19]),
    .c(cout_3[18]),
    .cout(cout_3[19]),
    .sum(sum_3[19]));
  AL_FADD comp3_2 (
    .a(i3[2]),
    .b(sum_2[2]),
    .c(cout_3[1]),
    .cout(cout_3[2]),
    .sum(sum_3[2]));
  AL_FADD comp3_20 (
    .a(i3[20]),
    .b(sum_2[20]),
    .c(cout_3[19]),
    .cout(cout_3[20]),
    .sum(sum_3[20]));
  AL_FADD comp3_21 (
    .a(i3[21]),
    .b(sum_2[21]),
    .c(cout_3[20]),
    .cout(cout_3[21]),
    .sum(sum_3[21]));
  AL_FADD comp3_22 (
    .a(i3[22]),
    .b(sum_2[22]),
    .c(cout_3[21]),
    .cout(cout_3[22]),
    .sum(sum_3[22]));
  AL_FADD comp3_23 (
    .a(i3[23]),
    .b(sum_2[23]),
    .c(cout_3[22]),
    .cout(cout_3[23]),
    .sum(sum_3[23]));
  AL_FADD comp3_24 (
    .a(i3[24]),
    .b(sum_2[24]),
    .c(cout_3[23]),
    .cout(cout_3[24]),
    .sum(sum_3[24]));
  AL_FADD comp3_25 (
    .a(i3[25]),
    .b(sum_2[25]),
    .c(cout_3[24]),
    .cout(cout_3[25]),
    .sum(sum_3[25]));
  AL_FADD comp3_26 (
    .a(i3[26]),
    .b(sum_2[26]),
    .c(cout_3[25]),
    .cout(cout_3[26]),
    .sum(sum_3[26]));
  AL_FADD comp3_27 (
    .a(i3[27]),
    .b(sum_2[27]),
    .c(cout_3[26]),
    .cout(cout_3[27]),
    .sum(sum_3[27]));
  AL_FADD comp3_28 (
    .a(i3[28]),
    .b(sum_2[28]),
    .c(cout_3[27]),
    .cout(cout_3[28]),
    .sum(sum_3[28]));
  AL_FADD comp3_29 (
    .a(i3[29]),
    .b(sum_2[29]),
    .c(cout_3[28]),
    .cout(cout_3[29]),
    .sum(sum_3[29]));
  AL_FADD comp3_3 (
    .a(i3[3]),
    .b(sum_2[3]),
    .c(cout_3[2]),
    .cout(cout_3[3]),
    .sum(sum_3[3]));
  AL_FADD comp3_30 (
    .a(i3[30]),
    .b(sum_2[30]),
    .c(cout_3[29]),
    .cout(cout_3[30]),
    .sum(sum_3[30]));
  AL_FADD comp3_31 (
    .a(i3[31]),
    .b(sum_2[31]),
    .c(cout_3[30]),
    .cout(cout_3[31]),
    .sum(sum_3[31]));
  AL_FADD comp3_32 (
    .a(i3[32]),
    .b(sum_2[32]),
    .c(cout_3[31]),
    .cout(cout_3[32]),
    .sum(sum_3[32]));
  AL_FADD comp3_33 (
    .a(i3[33]),
    .b(sum_2[33]),
    .c(cout_3[32]),
    .cout(cout_3[33]),
    .sum(sum_3[33]));
  AL_FADD comp3_34 (
    .a(i3[34]),
    .b(sum_2[34]),
    .c(cout_3[33]),
    .cout(cout_3[34]),
    .sum(sum_3[34]));
  AL_FADD comp3_35 (
    .a(i3[35]),
    .b(sum_2[35]),
    .c(cout_3[34]),
    .cout(cout_3[35]),
    .sum(sum_3[35]));
  AL_FADD comp3_36 (
    .a(i3[36]),
    .b(sum_2[36]),
    .c(cout_3[35]),
    .cout(cout_3[36]),
    .sum(sum_3[36]));
  AL_FADD comp3_37 (
    .a(i3[37]),
    .b(sum_2[37]),
    .c(cout_3[36]),
    .cout(cout_3[37]),
    .sum(sum_3[37]));
  AL_FADD comp3_38 (
    .a(i3[38]),
    .b(sum_2[38]),
    .c(cout_3[37]),
    .cout(cout_3[38]),
    .sum(sum_3[38]));
  AL_FADD comp3_39 (
    .a(i3[39]),
    .b(sum_2[39]),
    .c(cout_3[38]),
    .cout(cout_3[39]),
    .sum(sum_3[39]));
  AL_FADD comp3_4 (
    .a(i3[4]),
    .b(sum_2[4]),
    .c(cout_3[3]),
    .cout(cout_3[4]),
    .sum(sum_3[4]));
  AL_FADD comp3_40 (
    .a(i3[40]),
    .b(sum_2[40]),
    .c(cout_3[39]),
    .cout(cout_3[40]),
    .sum(sum_3[40]));
  AL_FADD comp3_41 (
    .a(i3[41]),
    .b(sum_2[41]),
    .c(cout_3[40]),
    .cout(cout_3[41]),
    .sum(sum_3[41]));
  AL_FADD comp3_42 (
    .a(i3[42]),
    .b(sum_2[42]),
    .c(cout_3[41]),
    .cout(cout_3[42]),
    .sum(sum_3[42]));
  AL_FADD comp3_43 (
    .a(i3[43]),
    .b(sum_2[43]),
    .c(cout_3[42]),
    .cout(cout_3[43]),
    .sum(sum_3[43]));
  AL_FADD comp3_44 (
    .a(1'b0),
    .b(sum_2[44]),
    .c(cout_3[43]),
    .cout(cout_3[44]),
    .sum(sum_3[44]));
  AL_FADD comp3_45 (
    .a(1'b0),
    .b(sum_2[45]),
    .c(cout_3[44]),
    .cout(cout_3[45]),
    .sum(sum_3[45]));
  AL_FADD comp3_46 (
    .a(1'b0),
    .b(sum_2[46]),
    .c(cout_3[45]),
    .cout(cout_3[46]),
    .sum(sum_3[46]));
  AL_FADD comp3_47 (
    .a(1'b0),
    .b(sum_2[47]),
    .c(cout_3[46]),
    .cout(cout_3[47]),
    .sum(sum_3[47]));
  AL_FADD comp3_5 (
    .a(i3[5]),
    .b(sum_2[5]),
    .c(cout_3[4]),
    .cout(cout_3[5]),
    .sum(sum_3[5]));
  AL_FADD comp3_6 (
    .a(i3[6]),
    .b(sum_2[6]),
    .c(cout_3[5]),
    .cout(cout_3[6]),
    .sum(sum_3[6]));
  AL_FADD comp3_7 (
    .a(i3[7]),
    .b(sum_2[7]),
    .c(cout_3[6]),
    .cout(cout_3[7]),
    .sum(sum_3[7]));
  AL_FADD comp3_8 (
    .a(i3[8]),
    .b(sum_2[8]),
    .c(cout_3[7]),
    .cout(cout_3[8]),
    .sum(sum_3[8]));
  AL_FADD comp3_9 (
    .a(i3[9]),
    .b(sum_2[9]),
    .c(cout_3[8]),
    .cout(cout_3[9]),
    .sum(sum_3[9]));
  AL_FADD comp4_0 (
    .a(i4[0]),
    .b(sum_3[0]),
    .c(1'b0),
    .cout(cout_4[0]),
    .sum(sum_4[0]));
  AL_FADD comp4_1 (
    .a(i4[1]),
    .b(sum_3[1]),
    .c(cout_4[0]),
    .cout(cout_4[1]),
    .sum(sum_4[1]));
  AL_FADD comp4_10 (
    .a(i4[10]),
    .b(sum_3[10]),
    .c(cout_4[9]),
    .cout(cout_4[10]),
    .sum(sum_4[10]));
  AL_FADD comp4_11 (
    .a(i4[11]),
    .b(sum_3[11]),
    .c(cout_4[10]),
    .cout(cout_4[11]),
    .sum(sum_4[11]));
  AL_FADD comp4_12 (
    .a(i4[12]),
    .b(sum_3[12]),
    .c(cout_4[11]),
    .cout(cout_4[12]),
    .sum(sum_4[12]));
  AL_FADD comp4_13 (
    .a(i4[13]),
    .b(sum_3[13]),
    .c(cout_4[12]),
    .cout(cout_4[13]),
    .sum(sum_4[13]));
  AL_FADD comp4_14 (
    .a(i4[14]),
    .b(sum_3[14]),
    .c(cout_4[13]),
    .cout(cout_4[14]),
    .sum(sum_4[14]));
  AL_FADD comp4_15 (
    .a(i4[15]),
    .b(sum_3[15]),
    .c(cout_4[14]),
    .cout(cout_4[15]),
    .sum(sum_4[15]));
  AL_FADD comp4_16 (
    .a(i4[16]),
    .b(sum_3[16]),
    .c(cout_4[15]),
    .cout(cout_4[16]),
    .sum(sum_4[16]));
  AL_FADD comp4_17 (
    .a(i4[17]),
    .b(sum_3[17]),
    .c(cout_4[16]),
    .cout(cout_4[17]),
    .sum(sum_4[17]));
  AL_FADD comp4_18 (
    .a(i4[18]),
    .b(sum_3[18]),
    .c(cout_4[17]),
    .cout(cout_4[18]),
    .sum(sum_4[18]));
  AL_FADD comp4_19 (
    .a(i4[19]),
    .b(sum_3[19]),
    .c(cout_4[18]),
    .cout(cout_4[19]),
    .sum(sum_4[19]));
  AL_FADD comp4_2 (
    .a(i4[2]),
    .b(sum_3[2]),
    .c(cout_4[1]),
    .cout(cout_4[2]),
    .sum(sum_4[2]));
  AL_FADD comp4_20 (
    .a(i4[20]),
    .b(sum_3[20]),
    .c(cout_4[19]),
    .cout(cout_4[20]),
    .sum(sum_4[20]));
  AL_FADD comp4_21 (
    .a(i4[21]),
    .b(sum_3[21]),
    .c(cout_4[20]),
    .cout(cout_4[21]),
    .sum(sum_4[21]));
  AL_FADD comp4_22 (
    .a(i4[22]),
    .b(sum_3[22]),
    .c(cout_4[21]),
    .cout(cout_4[22]),
    .sum(sum_4[22]));
  AL_FADD comp4_23 (
    .a(i4[23]),
    .b(sum_3[23]),
    .c(cout_4[22]),
    .cout(cout_4[23]),
    .sum(sum_4[23]));
  AL_FADD comp4_24 (
    .a(i4[24]),
    .b(sum_3[24]),
    .c(cout_4[23]),
    .cout(cout_4[24]),
    .sum(sum_4[24]));
  AL_FADD comp4_25 (
    .a(i4[25]),
    .b(sum_3[25]),
    .c(cout_4[24]),
    .cout(cout_4[25]),
    .sum(sum_4[25]));
  AL_FADD comp4_26 (
    .a(i4[26]),
    .b(sum_3[26]),
    .c(cout_4[25]),
    .cout(cout_4[26]),
    .sum(sum_4[26]));
  AL_FADD comp4_27 (
    .a(i4[27]),
    .b(sum_3[27]),
    .c(cout_4[26]),
    .cout(cout_4[27]),
    .sum(sum_4[27]));
  AL_FADD comp4_28 (
    .a(i4[28]),
    .b(sum_3[28]),
    .c(cout_4[27]),
    .cout(cout_4[28]),
    .sum(sum_4[28]));
  AL_FADD comp4_29 (
    .a(i4[29]),
    .b(sum_3[29]),
    .c(cout_4[28]),
    .cout(cout_4[29]),
    .sum(sum_4[29]));
  AL_FADD comp4_3 (
    .a(i4[3]),
    .b(sum_3[3]),
    .c(cout_4[2]),
    .cout(cout_4[3]),
    .sum(sum_4[3]));
  AL_FADD comp4_30 (
    .a(i4[30]),
    .b(sum_3[30]),
    .c(cout_4[29]),
    .cout(cout_4[30]),
    .sum(sum_4[30]));
  AL_FADD comp4_31 (
    .a(i4[31]),
    .b(sum_3[31]),
    .c(cout_4[30]),
    .cout(cout_4[31]),
    .sum(sum_4[31]));
  AL_FADD comp4_32 (
    .a(i4[32]),
    .b(sum_3[32]),
    .c(cout_4[31]),
    .cout(cout_4[32]),
    .sum(sum_4[32]));
  AL_FADD comp4_33 (
    .a(i4[33]),
    .b(sum_3[33]),
    .c(cout_4[32]),
    .cout(cout_4[33]),
    .sum(sum_4[33]));
  AL_FADD comp4_34 (
    .a(i4[34]),
    .b(sum_3[34]),
    .c(cout_4[33]),
    .cout(cout_4[34]),
    .sum(sum_4[34]));
  AL_FADD comp4_35 (
    .a(i4[35]),
    .b(sum_3[35]),
    .c(cout_4[34]),
    .cout(cout_4[35]),
    .sum(sum_4[35]));
  AL_FADD comp4_36 (
    .a(i4[36]),
    .b(sum_3[36]),
    .c(cout_4[35]),
    .cout(cout_4[36]),
    .sum(sum_4[36]));
  AL_FADD comp4_37 (
    .a(i4[37]),
    .b(sum_3[37]),
    .c(cout_4[36]),
    .cout(cout_4[37]),
    .sum(sum_4[37]));
  AL_FADD comp4_38 (
    .a(i4[38]),
    .b(sum_3[38]),
    .c(cout_4[37]),
    .cout(cout_4[38]),
    .sum(sum_4[38]));
  AL_FADD comp4_39 (
    .a(i4[39]),
    .b(sum_3[39]),
    .c(cout_4[38]),
    .cout(cout_4[39]),
    .sum(sum_4[39]));
  AL_FADD comp4_4 (
    .a(i4[4]),
    .b(sum_3[4]),
    .c(cout_4[3]),
    .cout(cout_4[4]),
    .sum(sum_4[4]));
  AL_FADD comp4_40 (
    .a(i4[40]),
    .b(sum_3[40]),
    .c(cout_4[39]),
    .cout(cout_4[40]),
    .sum(sum_4[40]));
  AL_FADD comp4_41 (
    .a(i4[41]),
    .b(sum_3[41]),
    .c(cout_4[40]),
    .cout(cout_4[41]),
    .sum(sum_4[41]));
  AL_FADD comp4_42 (
    .a(i4[42]),
    .b(sum_3[42]),
    .c(cout_4[41]),
    .cout(cout_4[42]),
    .sum(sum_4[42]));
  AL_FADD comp4_43 (
    .a(1'b0),
    .b(sum_3[43]),
    .c(cout_4[42]),
    .cout(cout_4[43]),
    .sum(sum_4[43]));
  AL_FADD comp4_44 (
    .a(1'b0),
    .b(sum_3[44]),
    .c(cout_4[43]),
    .cout(cout_4[44]),
    .sum(sum_4[44]));
  AL_FADD comp4_45 (
    .a(1'b0),
    .b(sum_3[45]),
    .c(cout_4[44]),
    .cout(cout_4[45]),
    .sum(sum_4[45]));
  AL_FADD comp4_46 (
    .a(1'b0),
    .b(sum_3[46]),
    .c(cout_4[45]),
    .cout(cout_4[46]),
    .sum(sum_4[46]));
  AL_FADD comp4_47 (
    .a(1'b0),
    .b(sum_3[47]),
    .c(cout_4[46]),
    .cout(cout_4[47]),
    .sum(sum_4[47]));
  AL_FADD comp4_5 (
    .a(i4[5]),
    .b(sum_3[5]),
    .c(cout_4[4]),
    .cout(cout_4[5]),
    .sum(sum_4[5]));
  AL_FADD comp4_6 (
    .a(i4[6]),
    .b(sum_3[6]),
    .c(cout_4[5]),
    .cout(cout_4[6]),
    .sum(sum_4[6]));
  AL_FADD comp4_7 (
    .a(i4[7]),
    .b(sum_3[7]),
    .c(cout_4[6]),
    .cout(cout_4[7]),
    .sum(sum_4[7]));
  AL_FADD comp4_8 (
    .a(i4[8]),
    .b(sum_3[8]),
    .c(cout_4[7]),
    .cout(cout_4[8]),
    .sum(sum_4[8]));
  AL_FADD comp4_9 (
    .a(i4[9]),
    .b(sum_3[9]),
    .c(cout_4[8]),
    .cout(cout_4[9]),
    .sum(sum_4[9]));
  AL_FADD comp5_0 (
    .a(i5[0]),
    .b(sum_4[0]),
    .c(1'b0),
    .cout(cout_5[0]),
    .sum(sum_5[0]));
  AL_FADD comp5_1 (
    .a(i5[1]),
    .b(sum_4[1]),
    .c(cout_5[0]),
    .cout(cout_5[1]),
    .sum(sum_5[1]));
  AL_FADD comp5_10 (
    .a(i5[10]),
    .b(sum_4[10]),
    .c(cout_5[9]),
    .cout(cout_5[10]),
    .sum(sum_5[10]));
  AL_FADD comp5_11 (
    .a(i5[11]),
    .b(sum_4[11]),
    .c(cout_5[10]),
    .cout(cout_5[11]),
    .sum(sum_5[11]));
  AL_FADD comp5_12 (
    .a(i5[12]),
    .b(sum_4[12]),
    .c(cout_5[11]),
    .cout(cout_5[12]),
    .sum(sum_5[12]));
  AL_FADD comp5_13 (
    .a(i5[13]),
    .b(sum_4[13]),
    .c(cout_5[12]),
    .cout(cout_5[13]),
    .sum(sum_5[13]));
  AL_FADD comp5_14 (
    .a(i5[14]),
    .b(sum_4[14]),
    .c(cout_5[13]),
    .cout(cout_5[14]),
    .sum(sum_5[14]));
  AL_FADD comp5_15 (
    .a(i5[15]),
    .b(sum_4[15]),
    .c(cout_5[14]),
    .cout(cout_5[15]),
    .sum(sum_5[15]));
  AL_FADD comp5_16 (
    .a(i5[16]),
    .b(sum_4[16]),
    .c(cout_5[15]),
    .cout(cout_5[16]),
    .sum(sum_5[16]));
  AL_FADD comp5_17 (
    .a(i5[17]),
    .b(sum_4[17]),
    .c(cout_5[16]),
    .cout(cout_5[17]),
    .sum(sum_5[17]));
  AL_FADD comp5_18 (
    .a(i5[18]),
    .b(sum_4[18]),
    .c(cout_5[17]),
    .cout(cout_5[18]),
    .sum(sum_5[18]));
  AL_FADD comp5_19 (
    .a(i5[19]),
    .b(sum_4[19]),
    .c(cout_5[18]),
    .cout(cout_5[19]),
    .sum(sum_5[19]));
  AL_FADD comp5_2 (
    .a(i5[2]),
    .b(sum_4[2]),
    .c(cout_5[1]),
    .cout(cout_5[2]),
    .sum(sum_5[2]));
  AL_FADD comp5_20 (
    .a(i5[20]),
    .b(sum_4[20]),
    .c(cout_5[19]),
    .cout(cout_5[20]),
    .sum(sum_5[20]));
  AL_FADD comp5_21 (
    .a(i5[21]),
    .b(sum_4[21]),
    .c(cout_5[20]),
    .cout(cout_5[21]),
    .sum(sum_5[21]));
  AL_FADD comp5_22 (
    .a(i5[22]),
    .b(sum_4[22]),
    .c(cout_5[21]),
    .cout(cout_5[22]),
    .sum(sum_5[22]));
  AL_FADD comp5_23 (
    .a(i5[23]),
    .b(sum_4[23]),
    .c(cout_5[22]),
    .cout(cout_5[23]),
    .sum(sum_5[23]));
  AL_FADD comp5_24 (
    .a(i5[24]),
    .b(sum_4[24]),
    .c(cout_5[23]),
    .cout(cout_5[24]),
    .sum(sum_5[24]));
  AL_FADD comp5_25 (
    .a(i5[25]),
    .b(sum_4[25]),
    .c(cout_5[24]),
    .cout(cout_5[25]),
    .sum(sum_5[25]));
  AL_FADD comp5_26 (
    .a(i5[26]),
    .b(sum_4[26]),
    .c(cout_5[25]),
    .cout(cout_5[26]),
    .sum(sum_5[26]));
  AL_FADD comp5_27 (
    .a(i5[27]),
    .b(sum_4[27]),
    .c(cout_5[26]),
    .cout(cout_5[27]),
    .sum(sum_5[27]));
  AL_FADD comp5_28 (
    .a(i5[28]),
    .b(sum_4[28]),
    .c(cout_5[27]),
    .cout(cout_5[28]),
    .sum(sum_5[28]));
  AL_FADD comp5_29 (
    .a(i5[29]),
    .b(sum_4[29]),
    .c(cout_5[28]),
    .cout(cout_5[29]),
    .sum(sum_5[29]));
  AL_FADD comp5_3 (
    .a(i5[3]),
    .b(sum_4[3]),
    .c(cout_5[2]),
    .cout(cout_5[3]),
    .sum(sum_5[3]));
  AL_FADD comp5_30 (
    .a(i5[30]),
    .b(sum_4[30]),
    .c(cout_5[29]),
    .cout(cout_5[30]),
    .sum(sum_5[30]));
  AL_FADD comp5_31 (
    .a(i5[31]),
    .b(sum_4[31]),
    .c(cout_5[30]),
    .cout(cout_5[31]),
    .sum(sum_5[31]));
  AL_FADD comp5_32 (
    .a(i5[32]),
    .b(sum_4[32]),
    .c(cout_5[31]),
    .cout(cout_5[32]),
    .sum(sum_5[32]));
  AL_FADD comp5_33 (
    .a(i5[33]),
    .b(sum_4[33]),
    .c(cout_5[32]),
    .cout(cout_5[33]),
    .sum(sum_5[33]));
  AL_FADD comp5_34 (
    .a(i5[34]),
    .b(sum_4[34]),
    .c(cout_5[33]),
    .cout(cout_5[34]),
    .sum(sum_5[34]));
  AL_FADD comp5_35 (
    .a(i5[35]),
    .b(sum_4[35]),
    .c(cout_5[34]),
    .cout(cout_5[35]),
    .sum(sum_5[35]));
  AL_FADD comp5_36 (
    .a(i5[36]),
    .b(sum_4[36]),
    .c(cout_5[35]),
    .cout(cout_5[36]),
    .sum(sum_5[36]));
  AL_FADD comp5_37 (
    .a(i5[37]),
    .b(sum_4[37]),
    .c(cout_5[36]),
    .cout(cout_5[37]),
    .sum(sum_5[37]));
  AL_FADD comp5_38 (
    .a(i5[38]),
    .b(sum_4[38]),
    .c(cout_5[37]),
    .cout(cout_5[38]),
    .sum(sum_5[38]));
  AL_FADD comp5_39 (
    .a(i5[39]),
    .b(sum_4[39]),
    .c(cout_5[38]),
    .cout(cout_5[39]),
    .sum(sum_5[39]));
  AL_FADD comp5_4 (
    .a(i5[4]),
    .b(sum_4[4]),
    .c(cout_5[3]),
    .cout(cout_5[4]),
    .sum(sum_5[4]));
  AL_FADD comp5_40 (
    .a(i5[40]),
    .b(sum_4[40]),
    .c(cout_5[39]),
    .cout(cout_5[40]),
    .sum(sum_5[40]));
  AL_FADD comp5_41 (
    .a(i5[41]),
    .b(sum_4[41]),
    .c(cout_5[40]),
    .cout(cout_5[41]),
    .sum(sum_5[41]));
  AL_FADD comp5_42 (
    .a(1'b0),
    .b(sum_4[42]),
    .c(cout_5[41]),
    .cout(cout_5[42]),
    .sum(sum_5[42]));
  AL_FADD comp5_43 (
    .a(1'b0),
    .b(sum_4[43]),
    .c(cout_5[42]),
    .cout(cout_5[43]),
    .sum(sum_5[43]));
  AL_FADD comp5_44 (
    .a(1'b0),
    .b(sum_4[44]),
    .c(cout_5[43]),
    .cout(cout_5[44]),
    .sum(sum_5[44]));
  AL_FADD comp5_45 (
    .a(1'b0),
    .b(sum_4[45]),
    .c(cout_5[44]),
    .cout(cout_5[45]),
    .sum(sum_5[45]));
  AL_FADD comp5_46 (
    .a(1'b0),
    .b(sum_4[46]),
    .c(cout_5[45]),
    .cout(cout_5[46]),
    .sum(sum_5[46]));
  AL_FADD comp5_47 (
    .a(1'b0),
    .b(sum_4[47]),
    .c(cout_5[46]),
    .cout(cout_5[47]),
    .sum(sum_5[47]));
  AL_FADD comp5_5 (
    .a(i5[5]),
    .b(sum_4[5]),
    .c(cout_5[4]),
    .cout(cout_5[5]),
    .sum(sum_5[5]));
  AL_FADD comp5_6 (
    .a(i5[6]),
    .b(sum_4[6]),
    .c(cout_5[5]),
    .cout(cout_5[6]),
    .sum(sum_5[6]));
  AL_FADD comp5_7 (
    .a(i5[7]),
    .b(sum_4[7]),
    .c(cout_5[6]),
    .cout(cout_5[7]),
    .sum(sum_5[7]));
  AL_FADD comp5_8 (
    .a(i5[8]),
    .b(sum_4[8]),
    .c(cout_5[7]),
    .cout(cout_5[8]),
    .sum(sum_5[8]));
  AL_FADD comp5_9 (
    .a(i5[9]),
    .b(sum_4[9]),
    .c(cout_5[8]),
    .cout(cout_5[9]),
    .sum(sum_5[9]));
  AL_FADD comp6_0 (
    .a(i6[0]),
    .b(sum_5[0]),
    .c(1'b0),
    .cout(cout_6[0]),
    .sum(sum_6[0]));
  AL_FADD comp6_1 (
    .a(i6[1]),
    .b(sum_5[1]),
    .c(cout_6[0]),
    .cout(cout_6[1]),
    .sum(sum_6[1]));
  AL_FADD comp6_10 (
    .a(i6[10]),
    .b(sum_5[10]),
    .c(cout_6[9]),
    .cout(cout_6[10]),
    .sum(sum_6[10]));
  AL_FADD comp6_11 (
    .a(i6[11]),
    .b(sum_5[11]),
    .c(cout_6[10]),
    .cout(cout_6[11]),
    .sum(sum_6[11]));
  AL_FADD comp6_12 (
    .a(i6[12]),
    .b(sum_5[12]),
    .c(cout_6[11]),
    .cout(cout_6[12]),
    .sum(sum_6[12]));
  AL_FADD comp6_13 (
    .a(i6[13]),
    .b(sum_5[13]),
    .c(cout_6[12]),
    .cout(cout_6[13]),
    .sum(sum_6[13]));
  AL_FADD comp6_14 (
    .a(i6[14]),
    .b(sum_5[14]),
    .c(cout_6[13]),
    .cout(cout_6[14]),
    .sum(sum_6[14]));
  AL_FADD comp6_15 (
    .a(i6[15]),
    .b(sum_5[15]),
    .c(cout_6[14]),
    .cout(cout_6[15]),
    .sum(sum_6[15]));
  AL_FADD comp6_16 (
    .a(i6[16]),
    .b(sum_5[16]),
    .c(cout_6[15]),
    .cout(cout_6[16]),
    .sum(sum_6[16]));
  AL_FADD comp6_17 (
    .a(i6[17]),
    .b(sum_5[17]),
    .c(cout_6[16]),
    .cout(cout_6[17]),
    .sum(sum_6[17]));
  AL_FADD comp6_18 (
    .a(i6[18]),
    .b(sum_5[18]),
    .c(cout_6[17]),
    .cout(cout_6[18]),
    .sum(sum_6[18]));
  AL_FADD comp6_19 (
    .a(i6[19]),
    .b(sum_5[19]),
    .c(cout_6[18]),
    .cout(cout_6[19]),
    .sum(sum_6[19]));
  AL_FADD comp6_2 (
    .a(i6[2]),
    .b(sum_5[2]),
    .c(cout_6[1]),
    .cout(cout_6[2]),
    .sum(sum_6[2]));
  AL_FADD comp6_20 (
    .a(i6[20]),
    .b(sum_5[20]),
    .c(cout_6[19]),
    .cout(cout_6[20]),
    .sum(sum_6[20]));
  AL_FADD comp6_21 (
    .a(i6[21]),
    .b(sum_5[21]),
    .c(cout_6[20]),
    .cout(cout_6[21]),
    .sum(sum_6[21]));
  AL_FADD comp6_22 (
    .a(i6[22]),
    .b(sum_5[22]),
    .c(cout_6[21]),
    .cout(cout_6[22]),
    .sum(sum_6[22]));
  AL_FADD comp6_23 (
    .a(i6[23]),
    .b(sum_5[23]),
    .c(cout_6[22]),
    .cout(cout_6[23]),
    .sum(sum_6[23]));
  AL_FADD comp6_24 (
    .a(i6[24]),
    .b(sum_5[24]),
    .c(cout_6[23]),
    .cout(cout_6[24]),
    .sum(sum_6[24]));
  AL_FADD comp6_25 (
    .a(i6[25]),
    .b(sum_5[25]),
    .c(cout_6[24]),
    .cout(cout_6[25]),
    .sum(sum_6[25]));
  AL_FADD comp6_26 (
    .a(i6[26]),
    .b(sum_5[26]),
    .c(cout_6[25]),
    .cout(cout_6[26]),
    .sum(sum_6[26]));
  AL_FADD comp6_27 (
    .a(i6[27]),
    .b(sum_5[27]),
    .c(cout_6[26]),
    .cout(cout_6[27]),
    .sum(sum_6[27]));
  AL_FADD comp6_28 (
    .a(i6[28]),
    .b(sum_5[28]),
    .c(cout_6[27]),
    .cout(cout_6[28]),
    .sum(sum_6[28]));
  AL_FADD comp6_29 (
    .a(i6[29]),
    .b(sum_5[29]),
    .c(cout_6[28]),
    .cout(cout_6[29]),
    .sum(sum_6[29]));
  AL_FADD comp6_3 (
    .a(i6[3]),
    .b(sum_5[3]),
    .c(cout_6[2]),
    .cout(cout_6[3]),
    .sum(sum_6[3]));
  AL_FADD comp6_30 (
    .a(i6[30]),
    .b(sum_5[30]),
    .c(cout_6[29]),
    .cout(cout_6[30]),
    .sum(sum_6[30]));
  AL_FADD comp6_31 (
    .a(i6[31]),
    .b(sum_5[31]),
    .c(cout_6[30]),
    .cout(cout_6[31]),
    .sum(sum_6[31]));
  AL_FADD comp6_32 (
    .a(i6[32]),
    .b(sum_5[32]),
    .c(cout_6[31]),
    .cout(cout_6[32]),
    .sum(sum_6[32]));
  AL_FADD comp6_33 (
    .a(i6[33]),
    .b(sum_5[33]),
    .c(cout_6[32]),
    .cout(cout_6[33]),
    .sum(sum_6[33]));
  AL_FADD comp6_34 (
    .a(i6[34]),
    .b(sum_5[34]),
    .c(cout_6[33]),
    .cout(cout_6[34]),
    .sum(sum_6[34]));
  AL_FADD comp6_35 (
    .a(i6[35]),
    .b(sum_5[35]),
    .c(cout_6[34]),
    .cout(cout_6[35]),
    .sum(sum_6[35]));
  AL_FADD comp6_36 (
    .a(i6[36]),
    .b(sum_5[36]),
    .c(cout_6[35]),
    .cout(cout_6[36]),
    .sum(sum_6[36]));
  AL_FADD comp6_37 (
    .a(i6[37]),
    .b(sum_5[37]),
    .c(cout_6[36]),
    .cout(cout_6[37]),
    .sum(sum_6[37]));
  AL_FADD comp6_38 (
    .a(i6[38]),
    .b(sum_5[38]),
    .c(cout_6[37]),
    .cout(cout_6[38]),
    .sum(sum_6[38]));
  AL_FADD comp6_39 (
    .a(i6[39]),
    .b(sum_5[39]),
    .c(cout_6[38]),
    .cout(cout_6[39]),
    .sum(sum_6[39]));
  AL_FADD comp6_4 (
    .a(i6[4]),
    .b(sum_5[4]),
    .c(cout_6[3]),
    .cout(cout_6[4]),
    .sum(sum_6[4]));
  AL_FADD comp6_40 (
    .a(i6[40]),
    .b(sum_5[40]),
    .c(cout_6[39]),
    .cout(cout_6[40]),
    .sum(sum_6[40]));
  AL_FADD comp6_41 (
    .a(1'b0),
    .b(sum_5[41]),
    .c(cout_6[40]),
    .cout(cout_6[41]),
    .sum(sum_6[41]));
  AL_FADD comp6_42 (
    .a(1'b0),
    .b(sum_5[42]),
    .c(cout_6[41]),
    .cout(cout_6[42]),
    .sum(sum_6[42]));
  AL_FADD comp6_43 (
    .a(1'b0),
    .b(sum_5[43]),
    .c(cout_6[42]),
    .cout(cout_6[43]),
    .sum(sum_6[43]));
  AL_FADD comp6_44 (
    .a(1'b0),
    .b(sum_5[44]),
    .c(cout_6[43]),
    .cout(cout_6[44]),
    .sum(sum_6[44]));
  AL_FADD comp6_45 (
    .a(1'b0),
    .b(sum_5[45]),
    .c(cout_6[44]),
    .cout(cout_6[45]),
    .sum(sum_6[45]));
  AL_FADD comp6_46 (
    .a(1'b0),
    .b(sum_5[46]),
    .c(cout_6[45]),
    .cout(cout_6[46]),
    .sum(sum_6[46]));
  AL_FADD comp6_47 (
    .a(1'b0),
    .b(sum_5[47]),
    .c(cout_6[46]),
    .cout(cout_6[47]),
    .sum(sum_6[47]));
  AL_FADD comp6_5 (
    .a(i6[5]),
    .b(sum_5[5]),
    .c(cout_6[4]),
    .cout(cout_6[5]),
    .sum(sum_6[5]));
  AL_FADD comp6_6 (
    .a(i6[6]),
    .b(sum_5[6]),
    .c(cout_6[5]),
    .cout(cout_6[6]),
    .sum(sum_6[6]));
  AL_FADD comp6_7 (
    .a(i6[7]),
    .b(sum_5[7]),
    .c(cout_6[6]),
    .cout(cout_6[7]),
    .sum(sum_6[7]));
  AL_FADD comp6_8 (
    .a(i6[8]),
    .b(sum_5[8]),
    .c(cout_6[7]),
    .cout(cout_6[8]),
    .sum(sum_6[8]));
  AL_FADD comp6_9 (
    .a(i6[9]),
    .b(sum_5[9]),
    .c(cout_6[8]),
    .cout(cout_6[9]),
    .sum(sum_6[9]));
  AL_FADD comp7_0 (
    .a(i7[0]),
    .b(sum_6[0]),
    .c(1'b0),
    .cout(cout_7[0]),
    .sum(sum_7[0]));
  AL_FADD comp7_1 (
    .a(i7[1]),
    .b(sum_6[1]),
    .c(cout_7[0]),
    .cout(cout_7[1]),
    .sum(sum_7[1]));
  AL_FADD comp7_10 (
    .a(i7[10]),
    .b(sum_6[10]),
    .c(cout_7[9]),
    .cout(cout_7[10]),
    .sum(sum_7[10]));
  AL_FADD comp7_11 (
    .a(i7[11]),
    .b(sum_6[11]),
    .c(cout_7[10]),
    .cout(cout_7[11]),
    .sum(sum_7[11]));
  AL_FADD comp7_12 (
    .a(i7[12]),
    .b(sum_6[12]),
    .c(cout_7[11]),
    .cout(cout_7[12]),
    .sum(sum_7[12]));
  AL_FADD comp7_13 (
    .a(i7[13]),
    .b(sum_6[13]),
    .c(cout_7[12]),
    .cout(cout_7[13]),
    .sum(sum_7[13]));
  AL_FADD comp7_14 (
    .a(i7[14]),
    .b(sum_6[14]),
    .c(cout_7[13]),
    .cout(cout_7[14]),
    .sum(sum_7[14]));
  AL_FADD comp7_15 (
    .a(i7[15]),
    .b(sum_6[15]),
    .c(cout_7[14]),
    .cout(cout_7[15]),
    .sum(sum_7[15]));
  AL_FADD comp7_16 (
    .a(i7[16]),
    .b(sum_6[16]),
    .c(cout_7[15]),
    .cout(cout_7[16]),
    .sum(sum_7[16]));
  AL_FADD comp7_17 (
    .a(i7[17]),
    .b(sum_6[17]),
    .c(cout_7[16]),
    .cout(cout_7[17]),
    .sum(sum_7[17]));
  AL_FADD comp7_18 (
    .a(i7[18]),
    .b(sum_6[18]),
    .c(cout_7[17]),
    .cout(cout_7[18]),
    .sum(sum_7[18]));
  AL_FADD comp7_19 (
    .a(i7[19]),
    .b(sum_6[19]),
    .c(cout_7[18]),
    .cout(cout_7[19]),
    .sum(sum_7[19]));
  AL_FADD comp7_2 (
    .a(i7[2]),
    .b(sum_6[2]),
    .c(cout_7[1]),
    .cout(cout_7[2]),
    .sum(sum_7[2]));
  AL_FADD comp7_20 (
    .a(i7[20]),
    .b(sum_6[20]),
    .c(cout_7[19]),
    .cout(cout_7[20]),
    .sum(sum_7[20]));
  AL_FADD comp7_21 (
    .a(i7[21]),
    .b(sum_6[21]),
    .c(cout_7[20]),
    .cout(cout_7[21]),
    .sum(sum_7[21]));
  AL_FADD comp7_22 (
    .a(i7[22]),
    .b(sum_6[22]),
    .c(cout_7[21]),
    .cout(cout_7[22]),
    .sum(sum_7[22]));
  AL_FADD comp7_23 (
    .a(i7[23]),
    .b(sum_6[23]),
    .c(cout_7[22]),
    .cout(cout_7[23]),
    .sum(sum_7[23]));
  AL_FADD comp7_24 (
    .a(i7[24]),
    .b(sum_6[24]),
    .c(cout_7[23]),
    .cout(cout_7[24]),
    .sum(sum_7[24]));
  AL_FADD comp7_25 (
    .a(i7[25]),
    .b(sum_6[25]),
    .c(cout_7[24]),
    .cout(cout_7[25]),
    .sum(sum_7[25]));
  AL_FADD comp7_26 (
    .a(i7[26]),
    .b(sum_6[26]),
    .c(cout_7[25]),
    .cout(cout_7[26]),
    .sum(sum_7[26]));
  AL_FADD comp7_27 (
    .a(i7[27]),
    .b(sum_6[27]),
    .c(cout_7[26]),
    .cout(cout_7[27]),
    .sum(sum_7[27]));
  AL_FADD comp7_28 (
    .a(i7[28]),
    .b(sum_6[28]),
    .c(cout_7[27]),
    .cout(cout_7[28]),
    .sum(sum_7[28]));
  AL_FADD comp7_29 (
    .a(i7[29]),
    .b(sum_6[29]),
    .c(cout_7[28]),
    .cout(cout_7[29]),
    .sum(sum_7[29]));
  AL_FADD comp7_3 (
    .a(i7[3]),
    .b(sum_6[3]),
    .c(cout_7[2]),
    .cout(cout_7[3]),
    .sum(sum_7[3]));
  AL_FADD comp7_30 (
    .a(i7[30]),
    .b(sum_6[30]),
    .c(cout_7[29]),
    .cout(cout_7[30]),
    .sum(sum_7[30]));
  AL_FADD comp7_31 (
    .a(i7[31]),
    .b(sum_6[31]),
    .c(cout_7[30]),
    .cout(cout_7[31]),
    .sum(sum_7[31]));
  AL_FADD comp7_32 (
    .a(i7[32]),
    .b(sum_6[32]),
    .c(cout_7[31]),
    .cout(cout_7[32]),
    .sum(sum_7[32]));
  AL_FADD comp7_33 (
    .a(i7[33]),
    .b(sum_6[33]),
    .c(cout_7[32]),
    .cout(cout_7[33]),
    .sum(sum_7[33]));
  AL_FADD comp7_34 (
    .a(i7[34]),
    .b(sum_6[34]),
    .c(cout_7[33]),
    .cout(cout_7[34]),
    .sum(sum_7[34]));
  AL_FADD comp7_35 (
    .a(i7[35]),
    .b(sum_6[35]),
    .c(cout_7[34]),
    .cout(cout_7[35]),
    .sum(sum_7[35]));
  AL_FADD comp7_36 (
    .a(i7[36]),
    .b(sum_6[36]),
    .c(cout_7[35]),
    .cout(cout_7[36]),
    .sum(sum_7[36]));
  AL_FADD comp7_37 (
    .a(i7[37]),
    .b(sum_6[37]),
    .c(cout_7[36]),
    .cout(cout_7[37]),
    .sum(sum_7[37]));
  AL_FADD comp7_38 (
    .a(i7[38]),
    .b(sum_6[38]),
    .c(cout_7[37]),
    .cout(cout_7[38]),
    .sum(sum_7[38]));
  AL_FADD comp7_39 (
    .a(i7[39]),
    .b(sum_6[39]),
    .c(cout_7[38]),
    .cout(cout_7[39]),
    .sum(sum_7[39]));
  AL_FADD comp7_4 (
    .a(i7[4]),
    .b(sum_6[4]),
    .c(cout_7[3]),
    .cout(cout_7[4]),
    .sum(sum_7[4]));
  AL_FADD comp7_40 (
    .a(1'b0),
    .b(sum_6[40]),
    .c(cout_7[39]),
    .cout(cout_7[40]),
    .sum(sum_7[40]));
  AL_FADD comp7_41 (
    .a(1'b0),
    .b(sum_6[41]),
    .c(cout_7[40]),
    .cout(cout_7[41]),
    .sum(sum_7[41]));
  AL_FADD comp7_42 (
    .a(1'b0),
    .b(sum_6[42]),
    .c(cout_7[41]),
    .cout(cout_7[42]),
    .sum(sum_7[42]));
  AL_FADD comp7_43 (
    .a(1'b0),
    .b(sum_6[43]),
    .c(cout_7[42]),
    .cout(cout_7[43]),
    .sum(sum_7[43]));
  AL_FADD comp7_44 (
    .a(1'b0),
    .b(sum_6[44]),
    .c(cout_7[43]),
    .cout(cout_7[44]),
    .sum(sum_7[44]));
  AL_FADD comp7_45 (
    .a(1'b0),
    .b(sum_6[45]),
    .c(cout_7[44]),
    .cout(cout_7[45]),
    .sum(sum_7[45]));
  AL_FADD comp7_46 (
    .a(1'b0),
    .b(sum_6[46]),
    .c(cout_7[45]),
    .cout(cout_7[46]),
    .sum(sum_7[46]));
  AL_FADD comp7_47 (
    .a(1'b0),
    .b(sum_6[47]),
    .c(cout_7[46]),
    .cout(cout_7[47]),
    .sum(sum_7[47]));
  AL_FADD comp7_5 (
    .a(i7[5]),
    .b(sum_6[5]),
    .c(cout_7[4]),
    .cout(cout_7[5]),
    .sum(sum_7[5]));
  AL_FADD comp7_6 (
    .a(i7[6]),
    .b(sum_6[6]),
    .c(cout_7[5]),
    .cout(cout_7[6]),
    .sum(sum_7[6]));
  AL_FADD comp7_7 (
    .a(i7[7]),
    .b(sum_6[7]),
    .c(cout_7[6]),
    .cout(cout_7[7]),
    .sum(sum_7[7]));
  AL_FADD comp7_8 (
    .a(i7[8]),
    .b(sum_6[8]),
    .c(cout_7[7]),
    .cout(cout_7[8]),
    .sum(sum_7[8]));
  AL_FADD comp7_9 (
    .a(i7[9]),
    .b(sum_6[9]),
    .c(cout_7[8]),
    .cout(cout_7[9]),
    .sum(sum_7[9]));
  AL_FADD comp8_0 (
    .a(i8[0]),
    .b(sum_7[0]),
    .c(1'b0),
    .cout(cout_8[0]),
    .sum(sum_8[0]));
  AL_FADD comp8_1 (
    .a(i8[1]),
    .b(sum_7[1]),
    .c(cout_8[0]),
    .cout(cout_8[1]),
    .sum(sum_8[1]));
  AL_FADD comp8_10 (
    .a(i8[10]),
    .b(sum_7[10]),
    .c(cout_8[9]),
    .cout(cout_8[10]),
    .sum(sum_8[10]));
  AL_FADD comp8_11 (
    .a(i8[11]),
    .b(sum_7[11]),
    .c(cout_8[10]),
    .cout(cout_8[11]),
    .sum(sum_8[11]));
  AL_FADD comp8_12 (
    .a(i8[12]),
    .b(sum_7[12]),
    .c(cout_8[11]),
    .cout(cout_8[12]),
    .sum(sum_8[12]));
  AL_FADD comp8_13 (
    .a(i8[13]),
    .b(sum_7[13]),
    .c(cout_8[12]),
    .cout(cout_8[13]),
    .sum(sum_8[13]));
  AL_FADD comp8_14 (
    .a(i8[14]),
    .b(sum_7[14]),
    .c(cout_8[13]),
    .cout(cout_8[14]),
    .sum(sum_8[14]));
  AL_FADD comp8_15 (
    .a(i8[15]),
    .b(sum_7[15]),
    .c(cout_8[14]),
    .cout(cout_8[15]),
    .sum(sum_8[15]));
  AL_FADD comp8_16 (
    .a(i8[16]),
    .b(sum_7[16]),
    .c(cout_8[15]),
    .cout(cout_8[16]),
    .sum(sum_8[16]));
  AL_FADD comp8_17 (
    .a(i8[17]),
    .b(sum_7[17]),
    .c(cout_8[16]),
    .cout(cout_8[17]),
    .sum(sum_8[17]));
  AL_FADD comp8_18 (
    .a(i8[18]),
    .b(sum_7[18]),
    .c(cout_8[17]),
    .cout(cout_8[18]),
    .sum(sum_8[18]));
  AL_FADD comp8_19 (
    .a(i8[19]),
    .b(sum_7[19]),
    .c(cout_8[18]),
    .cout(cout_8[19]),
    .sum(sum_8[19]));
  AL_FADD comp8_2 (
    .a(i8[2]),
    .b(sum_7[2]),
    .c(cout_8[1]),
    .cout(cout_8[2]),
    .sum(sum_8[2]));
  AL_FADD comp8_20 (
    .a(i8[20]),
    .b(sum_7[20]),
    .c(cout_8[19]),
    .cout(cout_8[20]),
    .sum(sum_8[20]));
  AL_FADD comp8_21 (
    .a(i8[21]),
    .b(sum_7[21]),
    .c(cout_8[20]),
    .cout(cout_8[21]),
    .sum(sum_8[21]));
  AL_FADD comp8_22 (
    .a(i8[22]),
    .b(sum_7[22]),
    .c(cout_8[21]),
    .cout(cout_8[22]),
    .sum(sum_8[22]));
  AL_FADD comp8_23 (
    .a(i8[23]),
    .b(sum_7[23]),
    .c(cout_8[22]),
    .cout(cout_8[23]),
    .sum(sum_8[23]));
  AL_FADD comp8_24 (
    .a(i8[24]),
    .b(sum_7[24]),
    .c(cout_8[23]),
    .cout(cout_8[24]),
    .sum(sum_8[24]));
  AL_FADD comp8_25 (
    .a(i8[25]),
    .b(sum_7[25]),
    .c(cout_8[24]),
    .cout(cout_8[25]),
    .sum(sum_8[25]));
  AL_FADD comp8_26 (
    .a(i8[26]),
    .b(sum_7[26]),
    .c(cout_8[25]),
    .cout(cout_8[26]),
    .sum(sum_8[26]));
  AL_FADD comp8_27 (
    .a(i8[27]),
    .b(sum_7[27]),
    .c(cout_8[26]),
    .cout(cout_8[27]),
    .sum(sum_8[27]));
  AL_FADD comp8_28 (
    .a(i8[28]),
    .b(sum_7[28]),
    .c(cout_8[27]),
    .cout(cout_8[28]),
    .sum(sum_8[28]));
  AL_FADD comp8_29 (
    .a(i8[29]),
    .b(sum_7[29]),
    .c(cout_8[28]),
    .cout(cout_8[29]),
    .sum(sum_8[29]));
  AL_FADD comp8_3 (
    .a(i8[3]),
    .b(sum_7[3]),
    .c(cout_8[2]),
    .cout(cout_8[3]),
    .sum(sum_8[3]));
  AL_FADD comp8_30 (
    .a(i8[30]),
    .b(sum_7[30]),
    .c(cout_8[29]),
    .cout(cout_8[30]),
    .sum(sum_8[30]));
  AL_FADD comp8_31 (
    .a(i8[31]),
    .b(sum_7[31]),
    .c(cout_8[30]),
    .cout(cout_8[31]),
    .sum(sum_8[31]));
  AL_FADD comp8_32 (
    .a(i8[32]),
    .b(sum_7[32]),
    .c(cout_8[31]),
    .cout(cout_8[32]),
    .sum(sum_8[32]));
  AL_FADD comp8_33 (
    .a(i8[33]),
    .b(sum_7[33]),
    .c(cout_8[32]),
    .cout(cout_8[33]),
    .sum(sum_8[33]));
  AL_FADD comp8_34 (
    .a(i8[34]),
    .b(sum_7[34]),
    .c(cout_8[33]),
    .cout(cout_8[34]),
    .sum(sum_8[34]));
  AL_FADD comp8_35 (
    .a(i8[35]),
    .b(sum_7[35]),
    .c(cout_8[34]),
    .cout(cout_8[35]),
    .sum(sum_8[35]));
  AL_FADD comp8_36 (
    .a(i8[36]),
    .b(sum_7[36]),
    .c(cout_8[35]),
    .cout(cout_8[36]),
    .sum(sum_8[36]));
  AL_FADD comp8_37 (
    .a(i8[37]),
    .b(sum_7[37]),
    .c(cout_8[36]),
    .cout(cout_8[37]),
    .sum(sum_8[37]));
  AL_FADD comp8_38 (
    .a(i8[38]),
    .b(sum_7[38]),
    .c(cout_8[37]),
    .cout(cout_8[38]),
    .sum(sum_8[38]));
  AL_FADD comp8_39 (
    .a(1'b0),
    .b(sum_7[39]),
    .c(cout_8[38]),
    .cout(cout_8[39]),
    .sum(sum_8[39]));
  AL_FADD comp8_4 (
    .a(i8[4]),
    .b(sum_7[4]),
    .c(cout_8[3]),
    .cout(cout_8[4]),
    .sum(sum_8[4]));
  AL_FADD comp8_40 (
    .a(1'b0),
    .b(sum_7[40]),
    .c(cout_8[39]),
    .cout(cout_8[40]),
    .sum(sum_8[40]));
  AL_FADD comp8_41 (
    .a(1'b0),
    .b(sum_7[41]),
    .c(cout_8[40]),
    .cout(cout_8[41]),
    .sum(sum_8[41]));
  AL_FADD comp8_42 (
    .a(1'b0),
    .b(sum_7[42]),
    .c(cout_8[41]),
    .cout(cout_8[42]),
    .sum(sum_8[42]));
  AL_FADD comp8_43 (
    .a(1'b0),
    .b(sum_7[43]),
    .c(cout_8[42]),
    .cout(cout_8[43]),
    .sum(sum_8[43]));
  AL_FADD comp8_44 (
    .a(1'b0),
    .b(sum_7[44]),
    .c(cout_8[43]),
    .cout(cout_8[44]),
    .sum(sum_8[44]));
  AL_FADD comp8_45 (
    .a(1'b0),
    .b(sum_7[45]),
    .c(cout_8[44]),
    .cout(cout_8[45]),
    .sum(sum_8[45]));
  AL_FADD comp8_46 (
    .a(1'b0),
    .b(sum_7[46]),
    .c(cout_8[45]),
    .cout(cout_8[46]),
    .sum(sum_8[46]));
  AL_FADD comp8_47 (
    .a(1'b0),
    .b(sum_7[47]),
    .c(cout_8[46]),
    .cout(cout_8[47]),
    .sum(sum_8[47]));
  AL_FADD comp8_5 (
    .a(i8[5]),
    .b(sum_7[5]),
    .c(cout_8[4]),
    .cout(cout_8[5]),
    .sum(sum_8[5]));
  AL_FADD comp8_6 (
    .a(i8[6]),
    .b(sum_7[6]),
    .c(cout_8[5]),
    .cout(cout_8[6]),
    .sum(sum_8[6]));
  AL_FADD comp8_7 (
    .a(i8[7]),
    .b(sum_7[7]),
    .c(cout_8[6]),
    .cout(cout_8[7]),
    .sum(sum_8[7]));
  AL_FADD comp8_8 (
    .a(i8[8]),
    .b(sum_7[8]),
    .c(cout_8[7]),
    .cout(cout_8[8]),
    .sum(sum_8[8]));
  AL_FADD comp8_9 (
    .a(i8[9]),
    .b(sum_7[9]),
    .c(cout_8[8]),
    .cout(cout_8[9]),
    .sum(sum_8[9]));
  AL_FADD comp9_0 (
    .a(i9[0]),
    .b(sum_8[0]),
    .c(1'b0),
    .cout(cout_9[0]),
    .sum(sum_9[0]));
  AL_FADD comp9_1 (
    .a(i9[1]),
    .b(sum_8[1]),
    .c(cout_9[0]),
    .cout(cout_9[1]),
    .sum(sum_9[1]));
  AL_FADD comp9_10 (
    .a(i9[10]),
    .b(sum_8[10]),
    .c(cout_9[9]),
    .cout(cout_9[10]),
    .sum(sum_9[10]));
  AL_FADD comp9_11 (
    .a(i9[11]),
    .b(sum_8[11]),
    .c(cout_9[10]),
    .cout(cout_9[11]),
    .sum(sum_9[11]));
  AL_FADD comp9_12 (
    .a(i9[12]),
    .b(sum_8[12]),
    .c(cout_9[11]),
    .cout(cout_9[12]),
    .sum(sum_9[12]));
  AL_FADD comp9_13 (
    .a(i9[13]),
    .b(sum_8[13]),
    .c(cout_9[12]),
    .cout(cout_9[13]),
    .sum(sum_9[13]));
  AL_FADD comp9_14 (
    .a(i9[14]),
    .b(sum_8[14]),
    .c(cout_9[13]),
    .cout(cout_9[14]),
    .sum(sum_9[14]));
  AL_FADD comp9_15 (
    .a(i9[15]),
    .b(sum_8[15]),
    .c(cout_9[14]),
    .cout(cout_9[15]),
    .sum(sum_9[15]));
  AL_FADD comp9_16 (
    .a(i9[16]),
    .b(sum_8[16]),
    .c(cout_9[15]),
    .cout(cout_9[16]),
    .sum(sum_9[16]));
  AL_FADD comp9_17 (
    .a(i9[17]),
    .b(sum_8[17]),
    .c(cout_9[16]),
    .cout(cout_9[17]),
    .sum(sum_9[17]));
  AL_FADD comp9_18 (
    .a(i9[18]),
    .b(sum_8[18]),
    .c(cout_9[17]),
    .cout(cout_9[18]),
    .sum(sum_9[18]));
  AL_FADD comp9_19 (
    .a(i9[19]),
    .b(sum_8[19]),
    .c(cout_9[18]),
    .cout(cout_9[19]),
    .sum(sum_9[19]));
  AL_FADD comp9_2 (
    .a(i9[2]),
    .b(sum_8[2]),
    .c(cout_9[1]),
    .cout(cout_9[2]),
    .sum(sum_9[2]));
  AL_FADD comp9_20 (
    .a(i9[20]),
    .b(sum_8[20]),
    .c(cout_9[19]),
    .cout(cout_9[20]),
    .sum(sum_9[20]));
  AL_FADD comp9_21 (
    .a(i9[21]),
    .b(sum_8[21]),
    .c(cout_9[20]),
    .cout(cout_9[21]),
    .sum(sum_9[21]));
  AL_FADD comp9_22 (
    .a(i9[22]),
    .b(sum_8[22]),
    .c(cout_9[21]),
    .cout(cout_9[22]),
    .sum(sum_9[22]));
  AL_FADD comp9_23 (
    .a(i9[23]),
    .b(sum_8[23]),
    .c(cout_9[22]),
    .cout(cout_9[23]),
    .sum(sum_9[23]));
  AL_FADD comp9_24 (
    .a(i9[24]),
    .b(sum_8[24]),
    .c(cout_9[23]),
    .cout(cout_9[24]),
    .sum(sum_9[24]));
  AL_FADD comp9_25 (
    .a(i9[25]),
    .b(sum_8[25]),
    .c(cout_9[24]),
    .cout(cout_9[25]),
    .sum(sum_9[25]));
  AL_FADD comp9_26 (
    .a(i9[26]),
    .b(sum_8[26]),
    .c(cout_9[25]),
    .cout(cout_9[26]),
    .sum(sum_9[26]));
  AL_FADD comp9_27 (
    .a(i9[27]),
    .b(sum_8[27]),
    .c(cout_9[26]),
    .cout(cout_9[27]),
    .sum(sum_9[27]));
  AL_FADD comp9_28 (
    .a(i9[28]),
    .b(sum_8[28]),
    .c(cout_9[27]),
    .cout(cout_9[28]),
    .sum(sum_9[28]));
  AL_FADD comp9_29 (
    .a(i9[29]),
    .b(sum_8[29]),
    .c(cout_9[28]),
    .cout(cout_9[29]),
    .sum(sum_9[29]));
  AL_FADD comp9_3 (
    .a(i9[3]),
    .b(sum_8[3]),
    .c(cout_9[2]),
    .cout(cout_9[3]),
    .sum(sum_9[3]));
  AL_FADD comp9_30 (
    .a(i9[30]),
    .b(sum_8[30]),
    .c(cout_9[29]),
    .cout(cout_9[30]),
    .sum(sum_9[30]));
  AL_FADD comp9_31 (
    .a(i9[31]),
    .b(sum_8[31]),
    .c(cout_9[30]),
    .cout(cout_9[31]),
    .sum(sum_9[31]));
  AL_FADD comp9_32 (
    .a(i9[32]),
    .b(sum_8[32]),
    .c(cout_9[31]),
    .cout(cout_9[32]),
    .sum(sum_9[32]));
  AL_FADD comp9_33 (
    .a(i9[33]),
    .b(sum_8[33]),
    .c(cout_9[32]),
    .cout(cout_9[33]),
    .sum(sum_9[33]));
  AL_FADD comp9_34 (
    .a(i9[34]),
    .b(sum_8[34]),
    .c(cout_9[33]),
    .cout(cout_9[34]),
    .sum(sum_9[34]));
  AL_FADD comp9_35 (
    .a(i9[35]),
    .b(sum_8[35]),
    .c(cout_9[34]),
    .cout(cout_9[35]),
    .sum(sum_9[35]));
  AL_FADD comp9_36 (
    .a(i9[36]),
    .b(sum_8[36]),
    .c(cout_9[35]),
    .cout(cout_9[36]),
    .sum(sum_9[36]));
  AL_FADD comp9_37 (
    .a(i9[37]),
    .b(sum_8[37]),
    .c(cout_9[36]),
    .cout(cout_9[37]),
    .sum(sum_9[37]));
  AL_FADD comp9_38 (
    .a(1'b0),
    .b(sum_8[38]),
    .c(cout_9[37]),
    .cout(cout_9[38]),
    .sum(sum_9[38]));
  AL_FADD comp9_39 (
    .a(1'b0),
    .b(sum_8[39]),
    .c(cout_9[38]),
    .cout(cout_9[39]),
    .sum(sum_9[39]));
  AL_FADD comp9_4 (
    .a(i9[4]),
    .b(sum_8[4]),
    .c(cout_9[3]),
    .cout(cout_9[4]),
    .sum(sum_9[4]));
  AL_FADD comp9_40 (
    .a(1'b0),
    .b(sum_8[40]),
    .c(cout_9[39]),
    .cout(cout_9[40]),
    .sum(sum_9[40]));
  AL_FADD comp9_41 (
    .a(1'b0),
    .b(sum_8[41]),
    .c(cout_9[40]),
    .cout(cout_9[41]),
    .sum(sum_9[41]));
  AL_FADD comp9_42 (
    .a(1'b0),
    .b(sum_8[42]),
    .c(cout_9[41]),
    .cout(cout_9[42]),
    .sum(sum_9[42]));
  AL_FADD comp9_43 (
    .a(1'b0),
    .b(sum_8[43]),
    .c(cout_9[42]),
    .cout(cout_9[43]),
    .sum(sum_9[43]));
  AL_FADD comp9_44 (
    .a(1'b0),
    .b(sum_8[44]),
    .c(cout_9[43]),
    .cout(cout_9[44]),
    .sum(sum_9[44]));
  AL_FADD comp9_45 (
    .a(1'b0),
    .b(sum_8[45]),
    .c(cout_9[44]),
    .cout(cout_9[45]),
    .sum(sum_9[45]));
  AL_FADD comp9_46 (
    .a(1'b0),
    .b(sum_8[46]),
    .c(cout_9[45]),
    .cout(cout_9[46]),
    .sum(sum_9[46]));
  AL_FADD comp9_47 (
    .a(1'b0),
    .b(sum_8[47]),
    .c(cout_9[46]),
    .cout(cout_9[47]),
    .sum(sum_9[47]));
  AL_FADD comp9_5 (
    .a(i9[5]),
    .b(sum_8[5]),
    .c(cout_9[4]),
    .cout(cout_9[5]),
    .sum(sum_9[5]));
  AL_FADD comp9_6 (
    .a(i9[6]),
    .b(sum_8[6]),
    .c(cout_9[5]),
    .cout(cout_9[6]),
    .sum(sum_9[6]));
  AL_FADD comp9_7 (
    .a(i9[7]),
    .b(sum_8[7]),
    .c(cout_9[6]),
    .cout(cout_9[7]),
    .sum(sum_9[7]));
  AL_FADD comp9_8 (
    .a(i9[8]),
    .b(sum_8[8]),
    .c(cout_9[7]),
    .cout(cout_9[8]),
    .sum(sum_9[8]));
  AL_FADD comp9_9 (
    .a(i9[9]),
    .b(sum_8[9]),
    .c(cout_9[8]),
    .cout(cout_9[9]),
    .sum(sum_9[9]));

endmodule 

module add_pu23_pu23_o23
  (
  i0,
  i1,
  o
  );

  input [22:0] i0;
  input [22:0] i1;
  output [22:0] o;

  wire net_a0;
  wire net_a1;
  wire net_a10;
  wire net_a11;
  wire net_a12;
  wire net_a13;
  wire net_a14;
  wire net_a15;
  wire net_a16;
  wire net_a17;
  wire net_a18;
  wire net_a19;
  wire net_a2;
  wire net_a20;
  wire net_a21;
  wire net_a22;
  wire net_a3;
  wire net_a4;
  wire net_a5;
  wire net_a6;
  wire net_a7;
  wire net_a8;
  wire net_a9;
  wire net_b0;
  wire net_b1;
  wire net_b10;
  wire net_b11;
  wire net_b12;
  wire net_b13;
  wire net_b14;
  wire net_b15;
  wire net_b16;
  wire net_b17;
  wire net_b18;
  wire net_b19;
  wire net_b2;
  wire net_b20;
  wire net_b21;
  wire net_b22;
  wire net_b3;
  wire net_b4;
  wire net_b5;
  wire net_b6;
  wire net_b7;
  wire net_b8;
  wire net_b9;
  wire net_cout0;
  wire net_cout1;
  wire net_cout10;
  wire net_cout11;
  wire net_cout12;
  wire net_cout13;
  wire net_cout14;
  wire net_cout15;
  wire net_cout16;
  wire net_cout17;
  wire net_cout18;
  wire net_cout19;
  wire net_cout2;
  wire net_cout20;
  wire net_cout21;
  wire net_cout22;
  wire net_cout3;
  wire net_cout4;
  wire net_cout5;
  wire net_cout6;
  wire net_cout7;
  wire net_cout8;
  wire net_cout9;
  wire net_sum0;
  wire net_sum1;
  wire net_sum10;
  wire net_sum11;
  wire net_sum12;
  wire net_sum13;
  wire net_sum14;
  wire net_sum15;
  wire net_sum16;
  wire net_sum17;
  wire net_sum18;
  wire net_sum19;
  wire net_sum2;
  wire net_sum20;
  wire net_sum21;
  wire net_sum22;
  wire net_sum3;
  wire net_sum4;
  wire net_sum5;
  wire net_sum6;
  wire net_sum7;
  wire net_sum8;
  wire net_sum9;

  assign net_a22 = i0[22];
  assign net_a21 = i0[21];
  assign net_a20 = i0[20];
  assign net_a19 = i0[19];
  assign net_a18 = i0[18];
  assign net_a17 = i0[17];
  assign net_a16 = i0[16];
  assign net_a15 = i0[15];
  assign net_a14 = i0[14];
  assign net_a13 = i0[13];
  assign net_a12 = i0[12];
  assign net_a11 = i0[11];
  assign net_a10 = i0[10];
  assign net_a9 = i0[9];
  assign net_a8 = i0[8];
  assign net_a7 = i0[7];
  assign net_a6 = i0[6];
  assign net_a5 = i0[5];
  assign net_a4 = i0[4];
  assign net_a3 = i0[3];
  assign net_a2 = i0[2];
  assign net_a1 = i0[1];
  assign net_a0 = i0[0];
  assign net_b22 = i1[22];
  assign net_b21 = i1[21];
  assign net_b20 = i1[20];
  assign net_b19 = i1[19];
  assign net_b18 = i1[18];
  assign net_b17 = i1[17];
  assign net_b16 = i1[16];
  assign net_b15 = i1[15];
  assign net_b14 = i1[14];
  assign net_b13 = i1[13];
  assign net_b12 = i1[12];
  assign net_b11 = i1[11];
  assign net_b10 = i1[10];
  assign net_b9 = i1[9];
  assign net_b8 = i1[8];
  assign net_b7 = i1[7];
  assign net_b6 = i1[6];
  assign net_b5 = i1[5];
  assign net_b4 = i1[4];
  assign net_b3 = i1[3];
  assign net_b2 = i1[2];
  assign net_b1 = i1[1];
  assign net_b0 = i1[0];
  assign o[22] = net_sum22;
  assign o[21] = net_sum21;
  assign o[20] = net_sum20;
  assign o[19] = net_sum19;
  assign o[18] = net_sum18;
  assign o[17] = net_sum17;
  assign o[16] = net_sum16;
  assign o[15] = net_sum15;
  assign o[14] = net_sum14;
  assign o[13] = net_sum13;
  assign o[12] = net_sum12;
  assign o[11] = net_sum11;
  assign o[10] = net_sum10;
  assign o[9] = net_sum9;
  assign o[8] = net_sum8;
  assign o[7] = net_sum7;
  assign o[6] = net_sum6;
  assign o[5] = net_sum5;
  assign o[4] = net_sum4;
  assign o[3] = net_sum3;
  assign o[2] = net_sum2;
  assign o[1] = net_sum1;
  assign o[0] = net_sum0;
  AL_FADD comp_0 (
    .a(net_a0),
    .b(net_b0),
    .c(1'b0),
    .cout(net_cout0),
    .sum(net_sum0));
  AL_FADD comp_1 (
    .a(net_a1),
    .b(net_b1),
    .c(net_cout0),
    .cout(net_cout1),
    .sum(net_sum1));
  AL_FADD comp_10 (
    .a(net_a10),
    .b(net_b10),
    .c(net_cout9),
    .cout(net_cout10),
    .sum(net_sum10));
  AL_FADD comp_11 (
    .a(net_a11),
    .b(net_b11),
    .c(net_cout10),
    .cout(net_cout11),
    .sum(net_sum11));
  AL_FADD comp_12 (
    .a(net_a12),
    .b(net_b12),
    .c(net_cout11),
    .cout(net_cout12),
    .sum(net_sum12));
  AL_FADD comp_13 (
    .a(net_a13),
    .b(net_b13),
    .c(net_cout12),
    .cout(net_cout13),
    .sum(net_sum13));
  AL_FADD comp_14 (
    .a(net_a14),
    .b(net_b14),
    .c(net_cout13),
    .cout(net_cout14),
    .sum(net_sum14));
  AL_FADD comp_15 (
    .a(net_a15),
    .b(net_b15),
    .c(net_cout14),
    .cout(net_cout15),
    .sum(net_sum15));
  AL_FADD comp_16 (
    .a(net_a16),
    .b(net_b16),
    .c(net_cout15),
    .cout(net_cout16),
    .sum(net_sum16));
  AL_FADD comp_17 (
    .a(net_a17),
    .b(net_b17),
    .c(net_cout16),
    .cout(net_cout17),
    .sum(net_sum17));
  AL_FADD comp_18 (
    .a(net_a18),
    .b(net_b18),
    .c(net_cout17),
    .cout(net_cout18),
    .sum(net_sum18));
  AL_FADD comp_19 (
    .a(net_a19),
    .b(net_b19),
    .c(net_cout18),
    .cout(net_cout19),
    .sum(net_sum19));
  AL_FADD comp_2 (
    .a(net_a2),
    .b(net_b2),
    .c(net_cout1),
    .cout(net_cout2),
    .sum(net_sum2));
  AL_FADD comp_20 (
    .a(net_a20),
    .b(net_b20),
    .c(net_cout19),
    .cout(net_cout20),
    .sum(net_sum20));
  AL_FADD comp_21 (
    .a(net_a21),
    .b(net_b21),
    .c(net_cout20),
    .cout(net_cout21),
    .sum(net_sum21));
  AL_FADD comp_22 (
    .a(net_a22),
    .b(net_b22),
    .c(net_cout21),
    .cout(net_cout22),
    .sum(net_sum22));
  AL_FADD comp_3 (
    .a(net_a3),
    .b(net_b3),
    .c(net_cout2),
    .cout(net_cout3),
    .sum(net_sum3));
  AL_FADD comp_4 (
    .a(net_a4),
    .b(net_b4),
    .c(net_cout3),
    .cout(net_cout4),
    .sum(net_sum4));
  AL_FADD comp_5 (
    .a(net_a5),
    .b(net_b5),
    .c(net_cout4),
    .cout(net_cout5),
    .sum(net_sum5));
  AL_FADD comp_6 (
    .a(net_a6),
    .b(net_b6),
    .c(net_cout5),
    .cout(net_cout6),
    .sum(net_sum6));
  AL_FADD comp_7 (
    .a(net_a7),
    .b(net_b7),
    .c(net_cout6),
    .cout(net_cout7),
    .sum(net_sum7));
  AL_FADD comp_8 (
    .a(net_a8),
    .b(net_b8),
    .c(net_cout7),
    .cout(net_cout8),
    .sum(net_sum8));
  AL_FADD comp_9 (
    .a(net_a9),
    .b(net_b9),
    .c(net_cout8),
    .cout(net_cout9),
    .sum(net_sum9));

endmodule 

module eq_w24
  (
  i0,
  i1,
  o
  );

  input [23:0] i0;
  input [23:0] i1;
  output o;

  wire \or_or_or_or_xor_i0[0_o ;
  wire \or_or_or_xor_i0[0]_i_o ;
  wire \or_or_or_xor_i0[12]__o ;
  wire \or_or_xor_i0[0]_i1[0_o ;
  wire \or_or_xor_i0[12]_i1[_o ;
  wire \or_or_xor_i0[18]_i1[_o ;
  wire \or_or_xor_i0[6]_i1[6_o ;
  wire \or_xor_i0[0]_i1[0]_o_o ;
  wire \or_xor_i0[10]_i1[10]_o ;
  wire \or_xor_i0[12]_i1[12]_o ;
  wire \or_xor_i0[13]_i1[13]_o ;
  wire \or_xor_i0[15]_i1[15]_o ;
  wire \or_xor_i0[16]_i1[16]_o ;
  wire \or_xor_i0[18]_i1[18]_o ;
  wire \or_xor_i0[19]_i1[19]_o ;
  wire \or_xor_i0[1]_i1[1]_o_o ;
  wire \or_xor_i0[21]_i1[21]_o ;
  wire \or_xor_i0[22]_i1[22]_o ;
  wire \or_xor_i0[3]_i1[3]_o_o ;
  wire \or_xor_i0[4]_i1[4]_o_o ;
  wire \or_xor_i0[6]_i1[6]_o_o ;
  wire \or_xor_i0[7]_i1[7]_o_o ;
  wire \or_xor_i0[9]_i1[9]_o_o ;
  wire \xor_i0[0]_i1[0]_o ;
  wire \xor_i0[10]_i1[10]_o ;
  wire \xor_i0[11]_i1[11]_o ;
  wire \xor_i0[12]_i1[12]_o ;
  wire \xor_i0[13]_i1[13]_o ;
  wire \xor_i0[14]_i1[14]_o ;
  wire \xor_i0[15]_i1[15]_o ;
  wire \xor_i0[16]_i1[16]_o ;
  wire \xor_i0[17]_i1[17]_o ;
  wire \xor_i0[18]_i1[18]_o ;
  wire \xor_i0[19]_i1[19]_o ;
  wire \xor_i0[1]_i1[1]_o ;
  wire \xor_i0[20]_i1[20]_o ;
  wire \xor_i0[21]_i1[21]_o ;
  wire \xor_i0[22]_i1[22]_o ;
  wire \xor_i0[23]_i1[23]_o ;
  wire \xor_i0[2]_i1[2]_o ;
  wire \xor_i0[3]_i1[3]_o ;
  wire \xor_i0[4]_i1[4]_o ;
  wire \xor_i0[5]_i1[5]_o ;
  wire \xor_i0[6]_i1[6]_o ;
  wire \xor_i0[7]_i1[7]_o ;
  wire \xor_i0[8]_i1[8]_o ;
  wire \xor_i0[9]_i1[9]_o ;

  not none_diff (o, \or_or_or_or_xor_i0[0_o );
  or \or_or_or_or_xor_i0[0  (\or_or_or_or_xor_i0[0_o , \or_or_or_xor_i0[0]_i_o , \or_or_or_xor_i0[12]__o );
  or \or_or_or_xor_i0[0]_i  (\or_or_or_xor_i0[0]_i_o , \or_or_xor_i0[0]_i1[0_o , \or_or_xor_i0[6]_i1[6_o );
  or \or_or_or_xor_i0[12]_  (\or_or_or_xor_i0[12]__o , \or_or_xor_i0[12]_i1[_o , \or_or_xor_i0[18]_i1[_o );
  or \or_or_xor_i0[0]_i1[0  (\or_or_xor_i0[0]_i1[0_o , \or_xor_i0[0]_i1[0]_o_o , \or_xor_i0[3]_i1[3]_o_o );
  or \or_or_xor_i0[12]_i1[  (\or_or_xor_i0[12]_i1[_o , \or_xor_i0[12]_i1[12]_o , \or_xor_i0[15]_i1[15]_o );
  or \or_or_xor_i0[18]_i1[  (\or_or_xor_i0[18]_i1[_o , \or_xor_i0[18]_i1[18]_o , \or_xor_i0[21]_i1[21]_o );
  or \or_or_xor_i0[6]_i1[6  (\or_or_xor_i0[6]_i1[6_o , \or_xor_i0[6]_i1[6]_o_o , \or_xor_i0[9]_i1[9]_o_o );
  or \or_xor_i0[0]_i1[0]_o  (\or_xor_i0[0]_i1[0]_o_o , \xor_i0[0]_i1[0]_o , \or_xor_i0[1]_i1[1]_o_o );
  or \or_xor_i0[10]_i1[10]  (\or_xor_i0[10]_i1[10]_o , \xor_i0[10]_i1[10]_o , \xor_i0[11]_i1[11]_o );
  or \or_xor_i0[12]_i1[12]  (\or_xor_i0[12]_i1[12]_o , \xor_i0[12]_i1[12]_o , \or_xor_i0[13]_i1[13]_o );
  or \or_xor_i0[13]_i1[13]  (\or_xor_i0[13]_i1[13]_o , \xor_i0[13]_i1[13]_o , \xor_i0[14]_i1[14]_o );
  or \or_xor_i0[15]_i1[15]  (\or_xor_i0[15]_i1[15]_o , \xor_i0[15]_i1[15]_o , \or_xor_i0[16]_i1[16]_o );
  or \or_xor_i0[16]_i1[16]  (\or_xor_i0[16]_i1[16]_o , \xor_i0[16]_i1[16]_o , \xor_i0[17]_i1[17]_o );
  or \or_xor_i0[18]_i1[18]  (\or_xor_i0[18]_i1[18]_o , \xor_i0[18]_i1[18]_o , \or_xor_i0[19]_i1[19]_o );
  or \or_xor_i0[19]_i1[19]  (\or_xor_i0[19]_i1[19]_o , \xor_i0[19]_i1[19]_o , \xor_i0[20]_i1[20]_o );
  or \or_xor_i0[1]_i1[1]_o  (\or_xor_i0[1]_i1[1]_o_o , \xor_i0[1]_i1[1]_o , \xor_i0[2]_i1[2]_o );
  or \or_xor_i0[21]_i1[21]  (\or_xor_i0[21]_i1[21]_o , \xor_i0[21]_i1[21]_o , \or_xor_i0[22]_i1[22]_o );
  or \or_xor_i0[22]_i1[22]  (\or_xor_i0[22]_i1[22]_o , \xor_i0[22]_i1[22]_o , \xor_i0[23]_i1[23]_o );
  or \or_xor_i0[3]_i1[3]_o  (\or_xor_i0[3]_i1[3]_o_o , \xor_i0[3]_i1[3]_o , \or_xor_i0[4]_i1[4]_o_o );
  or \or_xor_i0[4]_i1[4]_o  (\or_xor_i0[4]_i1[4]_o_o , \xor_i0[4]_i1[4]_o , \xor_i0[5]_i1[5]_o );
  or \or_xor_i0[6]_i1[6]_o  (\or_xor_i0[6]_i1[6]_o_o , \xor_i0[6]_i1[6]_o , \or_xor_i0[7]_i1[7]_o_o );
  or \or_xor_i0[7]_i1[7]_o  (\or_xor_i0[7]_i1[7]_o_o , \xor_i0[7]_i1[7]_o , \xor_i0[8]_i1[8]_o );
  or \or_xor_i0[9]_i1[9]_o  (\or_xor_i0[9]_i1[9]_o_o , \xor_i0[9]_i1[9]_o , \or_xor_i0[10]_i1[10]_o );
  xor \xor_i0[0]_i1[0]  (\xor_i0[0]_i1[0]_o , i0[0], i1[0]);
  xor \xor_i0[10]_i1[10]  (\xor_i0[10]_i1[10]_o , i0[10], i1[10]);
  xor \xor_i0[11]_i1[11]  (\xor_i0[11]_i1[11]_o , i0[11], i1[11]);
  xor \xor_i0[12]_i1[12]  (\xor_i0[12]_i1[12]_o , i0[12], i1[12]);
  xor \xor_i0[13]_i1[13]  (\xor_i0[13]_i1[13]_o , i0[13], i1[13]);
  xor \xor_i0[14]_i1[14]  (\xor_i0[14]_i1[14]_o , i0[14], i1[14]);
  xor \xor_i0[15]_i1[15]  (\xor_i0[15]_i1[15]_o , i0[15], i1[15]);
  xor \xor_i0[16]_i1[16]  (\xor_i0[16]_i1[16]_o , i0[16], i1[16]);
  xor \xor_i0[17]_i1[17]  (\xor_i0[17]_i1[17]_o , i0[17], i1[17]);
  xor \xor_i0[18]_i1[18]  (\xor_i0[18]_i1[18]_o , i0[18], i1[18]);
  xor \xor_i0[19]_i1[19]  (\xor_i0[19]_i1[19]_o , i0[19], i1[19]);
  xor \xor_i0[1]_i1[1]  (\xor_i0[1]_i1[1]_o , i0[1], i1[1]);
  xor \xor_i0[20]_i1[20]  (\xor_i0[20]_i1[20]_o , i0[20], i1[20]);
  xor \xor_i0[21]_i1[21]  (\xor_i0[21]_i1[21]_o , i0[21], i1[21]);
  xor \xor_i0[22]_i1[22]  (\xor_i0[22]_i1[22]_o , i0[22], i1[22]);
  xor \xor_i0[23]_i1[23]  (\xor_i0[23]_i1[23]_o , i0[23], i1[23]);
  xor \xor_i0[2]_i1[2]  (\xor_i0[2]_i1[2]_o , i0[2], i1[2]);
  xor \xor_i0[3]_i1[3]  (\xor_i0[3]_i1[3]_o , i0[3], i1[3]);
  xor \xor_i0[4]_i1[4]  (\xor_i0[4]_i1[4]_o , i0[4], i1[4]);
  xor \xor_i0[5]_i1[5]  (\xor_i0[5]_i1[5]_o , i0[5], i1[5]);
  xor \xor_i0[6]_i1[6]  (\xor_i0[6]_i1[6]_o , i0[6], i1[6]);
  xor \xor_i0[7]_i1[7]  (\xor_i0[7]_i1[7]_o , i0[7], i1[7]);
  xor \xor_i0[8]_i1[8]  (\xor_i0[8]_i1[8]_o , i0[8], i1[8]);
  xor \xor_i0[9]_i1[9]  (\xor_i0[9]_i1[9]_o , i0[9], i1[9]);

endmodule 

module add_pu63_pu60_pu59_pu58_pu57_pu56_pu55_pu54_pu53_pu52_pu51_pu50_pu49_pu48_pu47_pu46_pu45_pu44_pu43_pu42_pu41_pu40_pu39_pu38_pu37_pu36_pu35_pu34_pu33_pu32_pu31_mu62_mu62_o64
  (
  i0,
  i1,
  i10,
  i11,
  i12,
  i13,
  i14,
  i15,
  i16,
  i17,
  i18,
  i19,
  i2,
  i20,
  i21,
  i22,
  i23,
  i24,
  i25,
  i26,
  i27,
  i28,
  i29,
  i3,
  i30,
  i31,
  i32,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  o
  );

  input [62:0] i0;
  input [59:0] i1;
  input [50:0] i10;
  input [49:0] i11;
  input [48:0] i12;
  input [47:0] i13;
  input [46:0] i14;
  input [45:0] i15;
  input [44:0] i16;
  input [43:0] i17;
  input [42:0] i18;
  input [41:0] i19;
  input [58:0] i2;
  input [40:0] i20;
  input [39:0] i21;
  input [38:0] i22;
  input [37:0] i23;
  input [36:0] i24;
  input [35:0] i25;
  input [34:0] i26;
  input [33:0] i27;
  input [32:0] i28;
  input [31:0] i29;
  input [57:0] i3;
  input [30:0] i30;
  input [61:0] i31;
  input [61:0] i32;
  input [56:0] i4;
  input [55:0] i5;
  input [54:0] i6;
  input [53:0] i7;
  input [52:0] i8;
  input [51:0] i9;
  output [63:0] o;

  wire [62:0] cout_1;
  wire [63:0] cout_10;
  wire [63:0] cout_11;
  wire [63:0] cout_12;
  wire [63:0] cout_13;
  wire [63:0] cout_14;
  wire [63:0] cout_15;
  wire [63:0] cout_16;
  wire [63:0] cout_17;
  wire [63:0] cout_18;
  wire [63:0] cout_19;
  wire [63:0] cout_2;
  wire [63:0] cout_20;
  wire [63:0] cout_21;
  wire [63:0] cout_22;
  wire [63:0] cout_23;
  wire [63:0] cout_24;
  wire [63:0] cout_25;
  wire [63:0] cout_26;
  wire [63:0] cout_27;
  wire [63:0] cout_28;
  wire [63:0] cout_29;
  wire [63:0] cout_3;
  wire [63:0] cout_30;
  wire [63:0] cout_31;
  wire [63:0] cout_32;
  wire [63:0] cout_4;
  wire [63:0] cout_5;
  wire [63:0] cout_6;
  wire [63:0] cout_7;
  wire [63:0] cout_8;
  wire [63:0] cout_9;
  wire [62:0] sum_1;
  wire [63:0] sum_10;
  wire [63:0] sum_11;
  wire [63:0] sum_12;
  wire [63:0] sum_13;
  wire [63:0] sum_14;
  wire [63:0] sum_15;
  wire [63:0] sum_16;
  wire [63:0] sum_17;
  wire [63:0] sum_18;
  wire [63:0] sum_19;
  wire [63:0] sum_2;
  wire [63:0] sum_20;
  wire [63:0] sum_21;
  wire [63:0] sum_22;
  wire [63:0] sum_23;
  wire [63:0] sum_24;
  wire [63:0] sum_25;
  wire [63:0] sum_26;
  wire [63:0] sum_27;
  wire [63:0] sum_28;
  wire [63:0] sum_29;
  wire [63:0] sum_3;
  wire [63:0] sum_30;
  wire [63:0] sum_31;
  wire [63:0] sum_32;
  wire [63:0] sum_4;
  wire [63:0] sum_5;
  wire [63:0] sum_6;
  wire [63:0] sum_7;
  wire [63:0] sum_8;
  wire [63:0] sum_9;
  wire net_nb31_0;
  wire net_nb31_1;
  wire net_nb31_10;
  wire net_nb31_11;
  wire net_nb31_12;
  wire net_nb31_13;
  wire net_nb31_14;
  wire net_nb31_15;
  wire net_nb31_16;
  wire net_nb31_17;
  wire net_nb31_18;
  wire net_nb31_19;
  wire net_nb31_2;
  wire net_nb31_20;
  wire net_nb31_21;
  wire net_nb31_22;
  wire net_nb31_23;
  wire net_nb31_24;
  wire net_nb31_25;
  wire net_nb31_26;
  wire net_nb31_27;
  wire net_nb31_28;
  wire net_nb31_29;
  wire net_nb31_3;
  wire net_nb31_30;
  wire net_nb31_31;
  wire net_nb31_32;
  wire net_nb31_33;
  wire net_nb31_34;
  wire net_nb31_35;
  wire net_nb31_36;
  wire net_nb31_37;
  wire net_nb31_38;
  wire net_nb31_39;
  wire net_nb31_4;
  wire net_nb31_40;
  wire net_nb31_41;
  wire net_nb31_42;
  wire net_nb31_43;
  wire net_nb31_44;
  wire net_nb31_45;
  wire net_nb31_46;
  wire net_nb31_47;
  wire net_nb31_48;
  wire net_nb31_49;
  wire net_nb31_5;
  wire net_nb31_50;
  wire net_nb31_51;
  wire net_nb31_52;
  wire net_nb31_53;
  wire net_nb31_54;
  wire net_nb31_55;
  wire net_nb31_56;
  wire net_nb31_57;
  wire net_nb31_58;
  wire net_nb31_59;
  wire net_nb31_6;
  wire net_nb31_60;
  wire net_nb31_61;
  wire net_nb31_62;
  wire net_nb31_63;
  wire net_nb31_7;
  wire net_nb31_8;
  wire net_nb31_9;
  wire net_nb32_0;
  wire net_nb32_1;
  wire net_nb32_10;
  wire net_nb32_11;
  wire net_nb32_12;
  wire net_nb32_13;
  wire net_nb32_14;
  wire net_nb32_15;
  wire net_nb32_16;
  wire net_nb32_17;
  wire net_nb32_18;
  wire net_nb32_19;
  wire net_nb32_2;
  wire net_nb32_20;
  wire net_nb32_21;
  wire net_nb32_22;
  wire net_nb32_23;
  wire net_nb32_24;
  wire net_nb32_25;
  wire net_nb32_26;
  wire net_nb32_27;
  wire net_nb32_28;
  wire net_nb32_29;
  wire net_nb32_3;
  wire net_nb32_30;
  wire net_nb32_31;
  wire net_nb32_32;
  wire net_nb32_33;
  wire net_nb32_34;
  wire net_nb32_35;
  wire net_nb32_36;
  wire net_nb32_37;
  wire net_nb32_38;
  wire net_nb32_39;
  wire net_nb32_4;
  wire net_nb32_40;
  wire net_nb32_41;
  wire net_nb32_42;
  wire net_nb32_43;
  wire net_nb32_44;
  wire net_nb32_45;
  wire net_nb32_46;
  wire net_nb32_47;
  wire net_nb32_48;
  wire net_nb32_49;
  wire net_nb32_5;
  wire net_nb32_50;
  wire net_nb32_51;
  wire net_nb32_52;
  wire net_nb32_53;
  wire net_nb32_54;
  wire net_nb32_55;
  wire net_nb32_56;
  wire net_nb32_57;
  wire net_nb32_58;
  wire net_nb32_59;
  wire net_nb32_6;
  wire net_nb32_60;
  wire net_nb32_61;
  wire net_nb32_62;
  wire net_nb32_63;
  wire net_nb32_7;
  wire net_nb32_8;
  wire net_nb32_9;
  wire net_ncout31_63;
  wire net_ncout32_63;

  assign o[63] = sum_32[63];
  assign o[62] = sum_32[62];
  assign o[61] = sum_32[61];
  assign o[60] = sum_32[60];
  assign o[59] = sum_32[59];
  assign o[58] = sum_32[58];
  assign o[57] = sum_32[57];
  assign o[56] = sum_32[56];
  assign o[55] = sum_32[55];
  assign o[54] = sum_32[54];
  assign o[53] = sum_32[53];
  assign o[52] = sum_32[52];
  assign o[51] = sum_32[51];
  assign o[50] = sum_32[50];
  assign o[49] = sum_32[49];
  assign o[48] = sum_32[48];
  assign o[47] = sum_32[47];
  assign o[46] = sum_32[46];
  assign o[45] = sum_32[45];
  assign o[44] = sum_32[44];
  assign o[43] = sum_32[43];
  assign o[42] = sum_32[42];
  assign o[41] = sum_32[41];
  assign o[40] = sum_32[40];
  assign o[39] = sum_32[39];
  assign o[38] = sum_32[38];
  assign o[37] = sum_32[37];
  assign o[36] = sum_32[36];
  assign o[35] = sum_32[35];
  assign o[34] = sum_32[34];
  assign o[33] = sum_32[33];
  assign o[32] = sum_32[32];
  assign o[31] = sum_32[31];
  assign o[30] = sum_32[30];
  assign o[29] = sum_32[29];
  assign o[28] = sum_32[28];
  assign o[27] = sum_32[27];
  assign o[26] = sum_32[26];
  assign o[25] = sum_32[25];
  assign o[24] = sum_32[24];
  assign o[23] = sum_32[23];
  assign o[22] = sum_32[22];
  assign o[21] = sum_32[21];
  assign o[20] = sum_32[20];
  assign o[19] = sum_32[19];
  assign o[18] = sum_32[18];
  assign o[17] = sum_32[17];
  assign o[16] = sum_32[16];
  assign o[15] = sum_32[15];
  assign o[14] = sum_32[14];
  assign o[13] = sum_32[13];
  assign o[12] = sum_32[12];
  assign o[11] = sum_32[11];
  assign o[10] = sum_32[10];
  assign o[9] = sum_32[9];
  assign o[8] = sum_32[8];
  assign o[7] = sum_32[7];
  assign o[6] = sum_32[6];
  assign o[5] = sum_32[5];
  assign o[4] = sum_32[4];
  assign o[3] = sum_32[3];
  assign o[2] = sum_32[2];
  assign o[1] = sum_32[1];
  assign o[0] = sum_32[0];
  AL_FADD comp10_0 (
    .a(i10[0]),
    .b(sum_9[0]),
    .c(1'b0),
    .cout(cout_10[0]),
    .sum(sum_10[0]));
  AL_FADD comp10_1 (
    .a(i10[1]),
    .b(sum_9[1]),
    .c(cout_10[0]),
    .cout(cout_10[1]),
    .sum(sum_10[1]));
  AL_FADD comp10_10 (
    .a(i10[10]),
    .b(sum_9[10]),
    .c(cout_10[9]),
    .cout(cout_10[10]),
    .sum(sum_10[10]));
  AL_FADD comp10_11 (
    .a(i10[11]),
    .b(sum_9[11]),
    .c(cout_10[10]),
    .cout(cout_10[11]),
    .sum(sum_10[11]));
  AL_FADD comp10_12 (
    .a(i10[12]),
    .b(sum_9[12]),
    .c(cout_10[11]),
    .cout(cout_10[12]),
    .sum(sum_10[12]));
  AL_FADD comp10_13 (
    .a(i10[13]),
    .b(sum_9[13]),
    .c(cout_10[12]),
    .cout(cout_10[13]),
    .sum(sum_10[13]));
  AL_FADD comp10_14 (
    .a(i10[14]),
    .b(sum_9[14]),
    .c(cout_10[13]),
    .cout(cout_10[14]),
    .sum(sum_10[14]));
  AL_FADD comp10_15 (
    .a(i10[15]),
    .b(sum_9[15]),
    .c(cout_10[14]),
    .cout(cout_10[15]),
    .sum(sum_10[15]));
  AL_FADD comp10_16 (
    .a(i10[16]),
    .b(sum_9[16]),
    .c(cout_10[15]),
    .cout(cout_10[16]),
    .sum(sum_10[16]));
  AL_FADD comp10_17 (
    .a(i10[17]),
    .b(sum_9[17]),
    .c(cout_10[16]),
    .cout(cout_10[17]),
    .sum(sum_10[17]));
  AL_FADD comp10_18 (
    .a(i10[18]),
    .b(sum_9[18]),
    .c(cout_10[17]),
    .cout(cout_10[18]),
    .sum(sum_10[18]));
  AL_FADD comp10_19 (
    .a(i10[19]),
    .b(sum_9[19]),
    .c(cout_10[18]),
    .cout(cout_10[19]),
    .sum(sum_10[19]));
  AL_FADD comp10_2 (
    .a(i10[2]),
    .b(sum_9[2]),
    .c(cout_10[1]),
    .cout(cout_10[2]),
    .sum(sum_10[2]));
  AL_FADD comp10_20 (
    .a(i10[20]),
    .b(sum_9[20]),
    .c(cout_10[19]),
    .cout(cout_10[20]),
    .sum(sum_10[20]));
  AL_FADD comp10_21 (
    .a(i10[21]),
    .b(sum_9[21]),
    .c(cout_10[20]),
    .cout(cout_10[21]),
    .sum(sum_10[21]));
  AL_FADD comp10_22 (
    .a(i10[22]),
    .b(sum_9[22]),
    .c(cout_10[21]),
    .cout(cout_10[22]),
    .sum(sum_10[22]));
  AL_FADD comp10_23 (
    .a(i10[23]),
    .b(sum_9[23]),
    .c(cout_10[22]),
    .cout(cout_10[23]),
    .sum(sum_10[23]));
  AL_FADD comp10_24 (
    .a(i10[24]),
    .b(sum_9[24]),
    .c(cout_10[23]),
    .cout(cout_10[24]),
    .sum(sum_10[24]));
  AL_FADD comp10_25 (
    .a(i10[25]),
    .b(sum_9[25]),
    .c(cout_10[24]),
    .cout(cout_10[25]),
    .sum(sum_10[25]));
  AL_FADD comp10_26 (
    .a(i10[26]),
    .b(sum_9[26]),
    .c(cout_10[25]),
    .cout(cout_10[26]),
    .sum(sum_10[26]));
  AL_FADD comp10_27 (
    .a(i10[27]),
    .b(sum_9[27]),
    .c(cout_10[26]),
    .cout(cout_10[27]),
    .sum(sum_10[27]));
  AL_FADD comp10_28 (
    .a(i10[28]),
    .b(sum_9[28]),
    .c(cout_10[27]),
    .cout(cout_10[28]),
    .sum(sum_10[28]));
  AL_FADD comp10_29 (
    .a(i10[29]),
    .b(sum_9[29]),
    .c(cout_10[28]),
    .cout(cout_10[29]),
    .sum(sum_10[29]));
  AL_FADD comp10_3 (
    .a(i10[3]),
    .b(sum_9[3]),
    .c(cout_10[2]),
    .cout(cout_10[3]),
    .sum(sum_10[3]));
  AL_FADD comp10_30 (
    .a(i10[30]),
    .b(sum_9[30]),
    .c(cout_10[29]),
    .cout(cout_10[30]),
    .sum(sum_10[30]));
  AL_FADD comp10_31 (
    .a(i10[31]),
    .b(sum_9[31]),
    .c(cout_10[30]),
    .cout(cout_10[31]),
    .sum(sum_10[31]));
  AL_FADD comp10_32 (
    .a(i10[32]),
    .b(sum_9[32]),
    .c(cout_10[31]),
    .cout(cout_10[32]),
    .sum(sum_10[32]));
  AL_FADD comp10_33 (
    .a(i10[33]),
    .b(sum_9[33]),
    .c(cout_10[32]),
    .cout(cout_10[33]),
    .sum(sum_10[33]));
  AL_FADD comp10_34 (
    .a(i10[34]),
    .b(sum_9[34]),
    .c(cout_10[33]),
    .cout(cout_10[34]),
    .sum(sum_10[34]));
  AL_FADD comp10_35 (
    .a(i10[35]),
    .b(sum_9[35]),
    .c(cout_10[34]),
    .cout(cout_10[35]),
    .sum(sum_10[35]));
  AL_FADD comp10_36 (
    .a(i10[36]),
    .b(sum_9[36]),
    .c(cout_10[35]),
    .cout(cout_10[36]),
    .sum(sum_10[36]));
  AL_FADD comp10_37 (
    .a(i10[37]),
    .b(sum_9[37]),
    .c(cout_10[36]),
    .cout(cout_10[37]),
    .sum(sum_10[37]));
  AL_FADD comp10_38 (
    .a(i10[38]),
    .b(sum_9[38]),
    .c(cout_10[37]),
    .cout(cout_10[38]),
    .sum(sum_10[38]));
  AL_FADD comp10_39 (
    .a(i10[39]),
    .b(sum_9[39]),
    .c(cout_10[38]),
    .cout(cout_10[39]),
    .sum(sum_10[39]));
  AL_FADD comp10_4 (
    .a(i10[4]),
    .b(sum_9[4]),
    .c(cout_10[3]),
    .cout(cout_10[4]),
    .sum(sum_10[4]));
  AL_FADD comp10_40 (
    .a(i10[40]),
    .b(sum_9[40]),
    .c(cout_10[39]),
    .cout(cout_10[40]),
    .sum(sum_10[40]));
  AL_FADD comp10_41 (
    .a(i10[41]),
    .b(sum_9[41]),
    .c(cout_10[40]),
    .cout(cout_10[41]),
    .sum(sum_10[41]));
  AL_FADD comp10_42 (
    .a(i10[42]),
    .b(sum_9[42]),
    .c(cout_10[41]),
    .cout(cout_10[42]),
    .sum(sum_10[42]));
  AL_FADD comp10_43 (
    .a(i10[43]),
    .b(sum_9[43]),
    .c(cout_10[42]),
    .cout(cout_10[43]),
    .sum(sum_10[43]));
  AL_FADD comp10_44 (
    .a(i10[44]),
    .b(sum_9[44]),
    .c(cout_10[43]),
    .cout(cout_10[44]),
    .sum(sum_10[44]));
  AL_FADD comp10_45 (
    .a(i10[45]),
    .b(sum_9[45]),
    .c(cout_10[44]),
    .cout(cout_10[45]),
    .sum(sum_10[45]));
  AL_FADD comp10_46 (
    .a(i10[46]),
    .b(sum_9[46]),
    .c(cout_10[45]),
    .cout(cout_10[46]),
    .sum(sum_10[46]));
  AL_FADD comp10_47 (
    .a(i10[47]),
    .b(sum_9[47]),
    .c(cout_10[46]),
    .cout(cout_10[47]),
    .sum(sum_10[47]));
  AL_FADD comp10_48 (
    .a(i10[48]),
    .b(sum_9[48]),
    .c(cout_10[47]),
    .cout(cout_10[48]),
    .sum(sum_10[48]));
  AL_FADD comp10_49 (
    .a(i10[49]),
    .b(sum_9[49]),
    .c(cout_10[48]),
    .cout(cout_10[49]),
    .sum(sum_10[49]));
  AL_FADD comp10_5 (
    .a(i10[5]),
    .b(sum_9[5]),
    .c(cout_10[4]),
    .cout(cout_10[5]),
    .sum(sum_10[5]));
  AL_FADD comp10_50 (
    .a(i10[50]),
    .b(sum_9[50]),
    .c(cout_10[49]),
    .cout(cout_10[50]),
    .sum(sum_10[50]));
  AL_FADD comp10_51 (
    .a(1'b0),
    .b(sum_9[51]),
    .c(cout_10[50]),
    .cout(cout_10[51]),
    .sum(sum_10[51]));
  AL_FADD comp10_52 (
    .a(1'b0),
    .b(sum_9[52]),
    .c(cout_10[51]),
    .cout(cout_10[52]),
    .sum(sum_10[52]));
  AL_FADD comp10_53 (
    .a(1'b0),
    .b(sum_9[53]),
    .c(cout_10[52]),
    .cout(cout_10[53]),
    .sum(sum_10[53]));
  AL_FADD comp10_54 (
    .a(1'b0),
    .b(sum_9[54]),
    .c(cout_10[53]),
    .cout(cout_10[54]),
    .sum(sum_10[54]));
  AL_FADD comp10_55 (
    .a(1'b0),
    .b(sum_9[55]),
    .c(cout_10[54]),
    .cout(cout_10[55]),
    .sum(sum_10[55]));
  AL_FADD comp10_56 (
    .a(1'b0),
    .b(sum_9[56]),
    .c(cout_10[55]),
    .cout(cout_10[56]),
    .sum(sum_10[56]));
  AL_FADD comp10_57 (
    .a(1'b0),
    .b(sum_9[57]),
    .c(cout_10[56]),
    .cout(cout_10[57]),
    .sum(sum_10[57]));
  AL_FADD comp10_58 (
    .a(1'b0),
    .b(sum_9[58]),
    .c(cout_10[57]),
    .cout(cout_10[58]),
    .sum(sum_10[58]));
  AL_FADD comp10_59 (
    .a(1'b0),
    .b(sum_9[59]),
    .c(cout_10[58]),
    .cout(cout_10[59]),
    .sum(sum_10[59]));
  AL_FADD comp10_6 (
    .a(i10[6]),
    .b(sum_9[6]),
    .c(cout_10[5]),
    .cout(cout_10[6]),
    .sum(sum_10[6]));
  AL_FADD comp10_60 (
    .a(1'b0),
    .b(sum_9[60]),
    .c(cout_10[59]),
    .cout(cout_10[60]),
    .sum(sum_10[60]));
  AL_FADD comp10_61 (
    .a(1'b0),
    .b(sum_9[61]),
    .c(cout_10[60]),
    .cout(cout_10[61]),
    .sum(sum_10[61]));
  AL_FADD comp10_62 (
    .a(1'b0),
    .b(sum_9[62]),
    .c(cout_10[61]),
    .cout(cout_10[62]),
    .sum(sum_10[62]));
  AL_FADD comp10_63 (
    .a(1'b0),
    .b(sum_9[63]),
    .c(cout_10[62]),
    .cout(cout_10[63]),
    .sum(sum_10[63]));
  AL_FADD comp10_7 (
    .a(i10[7]),
    .b(sum_9[7]),
    .c(cout_10[6]),
    .cout(cout_10[7]),
    .sum(sum_10[7]));
  AL_FADD comp10_8 (
    .a(i10[8]),
    .b(sum_9[8]),
    .c(cout_10[7]),
    .cout(cout_10[8]),
    .sum(sum_10[8]));
  AL_FADD comp10_9 (
    .a(i10[9]),
    .b(sum_9[9]),
    .c(cout_10[8]),
    .cout(cout_10[9]),
    .sum(sum_10[9]));
  AL_FADD comp11_0 (
    .a(i11[0]),
    .b(sum_10[0]),
    .c(1'b0),
    .cout(cout_11[0]),
    .sum(sum_11[0]));
  AL_FADD comp11_1 (
    .a(i11[1]),
    .b(sum_10[1]),
    .c(cout_11[0]),
    .cout(cout_11[1]),
    .sum(sum_11[1]));
  AL_FADD comp11_10 (
    .a(i11[10]),
    .b(sum_10[10]),
    .c(cout_11[9]),
    .cout(cout_11[10]),
    .sum(sum_11[10]));
  AL_FADD comp11_11 (
    .a(i11[11]),
    .b(sum_10[11]),
    .c(cout_11[10]),
    .cout(cout_11[11]),
    .sum(sum_11[11]));
  AL_FADD comp11_12 (
    .a(i11[12]),
    .b(sum_10[12]),
    .c(cout_11[11]),
    .cout(cout_11[12]),
    .sum(sum_11[12]));
  AL_FADD comp11_13 (
    .a(i11[13]),
    .b(sum_10[13]),
    .c(cout_11[12]),
    .cout(cout_11[13]),
    .sum(sum_11[13]));
  AL_FADD comp11_14 (
    .a(i11[14]),
    .b(sum_10[14]),
    .c(cout_11[13]),
    .cout(cout_11[14]),
    .sum(sum_11[14]));
  AL_FADD comp11_15 (
    .a(i11[15]),
    .b(sum_10[15]),
    .c(cout_11[14]),
    .cout(cout_11[15]),
    .sum(sum_11[15]));
  AL_FADD comp11_16 (
    .a(i11[16]),
    .b(sum_10[16]),
    .c(cout_11[15]),
    .cout(cout_11[16]),
    .sum(sum_11[16]));
  AL_FADD comp11_17 (
    .a(i11[17]),
    .b(sum_10[17]),
    .c(cout_11[16]),
    .cout(cout_11[17]),
    .sum(sum_11[17]));
  AL_FADD comp11_18 (
    .a(i11[18]),
    .b(sum_10[18]),
    .c(cout_11[17]),
    .cout(cout_11[18]),
    .sum(sum_11[18]));
  AL_FADD comp11_19 (
    .a(i11[19]),
    .b(sum_10[19]),
    .c(cout_11[18]),
    .cout(cout_11[19]),
    .sum(sum_11[19]));
  AL_FADD comp11_2 (
    .a(i11[2]),
    .b(sum_10[2]),
    .c(cout_11[1]),
    .cout(cout_11[2]),
    .sum(sum_11[2]));
  AL_FADD comp11_20 (
    .a(i11[20]),
    .b(sum_10[20]),
    .c(cout_11[19]),
    .cout(cout_11[20]),
    .sum(sum_11[20]));
  AL_FADD comp11_21 (
    .a(i11[21]),
    .b(sum_10[21]),
    .c(cout_11[20]),
    .cout(cout_11[21]),
    .sum(sum_11[21]));
  AL_FADD comp11_22 (
    .a(i11[22]),
    .b(sum_10[22]),
    .c(cout_11[21]),
    .cout(cout_11[22]),
    .sum(sum_11[22]));
  AL_FADD comp11_23 (
    .a(i11[23]),
    .b(sum_10[23]),
    .c(cout_11[22]),
    .cout(cout_11[23]),
    .sum(sum_11[23]));
  AL_FADD comp11_24 (
    .a(i11[24]),
    .b(sum_10[24]),
    .c(cout_11[23]),
    .cout(cout_11[24]),
    .sum(sum_11[24]));
  AL_FADD comp11_25 (
    .a(i11[25]),
    .b(sum_10[25]),
    .c(cout_11[24]),
    .cout(cout_11[25]),
    .sum(sum_11[25]));
  AL_FADD comp11_26 (
    .a(i11[26]),
    .b(sum_10[26]),
    .c(cout_11[25]),
    .cout(cout_11[26]),
    .sum(sum_11[26]));
  AL_FADD comp11_27 (
    .a(i11[27]),
    .b(sum_10[27]),
    .c(cout_11[26]),
    .cout(cout_11[27]),
    .sum(sum_11[27]));
  AL_FADD comp11_28 (
    .a(i11[28]),
    .b(sum_10[28]),
    .c(cout_11[27]),
    .cout(cout_11[28]),
    .sum(sum_11[28]));
  AL_FADD comp11_29 (
    .a(i11[29]),
    .b(sum_10[29]),
    .c(cout_11[28]),
    .cout(cout_11[29]),
    .sum(sum_11[29]));
  AL_FADD comp11_3 (
    .a(i11[3]),
    .b(sum_10[3]),
    .c(cout_11[2]),
    .cout(cout_11[3]),
    .sum(sum_11[3]));
  AL_FADD comp11_30 (
    .a(i11[30]),
    .b(sum_10[30]),
    .c(cout_11[29]),
    .cout(cout_11[30]),
    .sum(sum_11[30]));
  AL_FADD comp11_31 (
    .a(i11[31]),
    .b(sum_10[31]),
    .c(cout_11[30]),
    .cout(cout_11[31]),
    .sum(sum_11[31]));
  AL_FADD comp11_32 (
    .a(i11[32]),
    .b(sum_10[32]),
    .c(cout_11[31]),
    .cout(cout_11[32]),
    .sum(sum_11[32]));
  AL_FADD comp11_33 (
    .a(i11[33]),
    .b(sum_10[33]),
    .c(cout_11[32]),
    .cout(cout_11[33]),
    .sum(sum_11[33]));
  AL_FADD comp11_34 (
    .a(i11[34]),
    .b(sum_10[34]),
    .c(cout_11[33]),
    .cout(cout_11[34]),
    .sum(sum_11[34]));
  AL_FADD comp11_35 (
    .a(i11[35]),
    .b(sum_10[35]),
    .c(cout_11[34]),
    .cout(cout_11[35]),
    .sum(sum_11[35]));
  AL_FADD comp11_36 (
    .a(i11[36]),
    .b(sum_10[36]),
    .c(cout_11[35]),
    .cout(cout_11[36]),
    .sum(sum_11[36]));
  AL_FADD comp11_37 (
    .a(i11[37]),
    .b(sum_10[37]),
    .c(cout_11[36]),
    .cout(cout_11[37]),
    .sum(sum_11[37]));
  AL_FADD comp11_38 (
    .a(i11[38]),
    .b(sum_10[38]),
    .c(cout_11[37]),
    .cout(cout_11[38]),
    .sum(sum_11[38]));
  AL_FADD comp11_39 (
    .a(i11[39]),
    .b(sum_10[39]),
    .c(cout_11[38]),
    .cout(cout_11[39]),
    .sum(sum_11[39]));
  AL_FADD comp11_4 (
    .a(i11[4]),
    .b(sum_10[4]),
    .c(cout_11[3]),
    .cout(cout_11[4]),
    .sum(sum_11[4]));
  AL_FADD comp11_40 (
    .a(i11[40]),
    .b(sum_10[40]),
    .c(cout_11[39]),
    .cout(cout_11[40]),
    .sum(sum_11[40]));
  AL_FADD comp11_41 (
    .a(i11[41]),
    .b(sum_10[41]),
    .c(cout_11[40]),
    .cout(cout_11[41]),
    .sum(sum_11[41]));
  AL_FADD comp11_42 (
    .a(i11[42]),
    .b(sum_10[42]),
    .c(cout_11[41]),
    .cout(cout_11[42]),
    .sum(sum_11[42]));
  AL_FADD comp11_43 (
    .a(i11[43]),
    .b(sum_10[43]),
    .c(cout_11[42]),
    .cout(cout_11[43]),
    .sum(sum_11[43]));
  AL_FADD comp11_44 (
    .a(i11[44]),
    .b(sum_10[44]),
    .c(cout_11[43]),
    .cout(cout_11[44]),
    .sum(sum_11[44]));
  AL_FADD comp11_45 (
    .a(i11[45]),
    .b(sum_10[45]),
    .c(cout_11[44]),
    .cout(cout_11[45]),
    .sum(sum_11[45]));
  AL_FADD comp11_46 (
    .a(i11[46]),
    .b(sum_10[46]),
    .c(cout_11[45]),
    .cout(cout_11[46]),
    .sum(sum_11[46]));
  AL_FADD comp11_47 (
    .a(i11[47]),
    .b(sum_10[47]),
    .c(cout_11[46]),
    .cout(cout_11[47]),
    .sum(sum_11[47]));
  AL_FADD comp11_48 (
    .a(i11[48]),
    .b(sum_10[48]),
    .c(cout_11[47]),
    .cout(cout_11[48]),
    .sum(sum_11[48]));
  AL_FADD comp11_49 (
    .a(i11[49]),
    .b(sum_10[49]),
    .c(cout_11[48]),
    .cout(cout_11[49]),
    .sum(sum_11[49]));
  AL_FADD comp11_5 (
    .a(i11[5]),
    .b(sum_10[5]),
    .c(cout_11[4]),
    .cout(cout_11[5]),
    .sum(sum_11[5]));
  AL_FADD comp11_50 (
    .a(1'b0),
    .b(sum_10[50]),
    .c(cout_11[49]),
    .cout(cout_11[50]),
    .sum(sum_11[50]));
  AL_FADD comp11_51 (
    .a(1'b0),
    .b(sum_10[51]),
    .c(cout_11[50]),
    .cout(cout_11[51]),
    .sum(sum_11[51]));
  AL_FADD comp11_52 (
    .a(1'b0),
    .b(sum_10[52]),
    .c(cout_11[51]),
    .cout(cout_11[52]),
    .sum(sum_11[52]));
  AL_FADD comp11_53 (
    .a(1'b0),
    .b(sum_10[53]),
    .c(cout_11[52]),
    .cout(cout_11[53]),
    .sum(sum_11[53]));
  AL_FADD comp11_54 (
    .a(1'b0),
    .b(sum_10[54]),
    .c(cout_11[53]),
    .cout(cout_11[54]),
    .sum(sum_11[54]));
  AL_FADD comp11_55 (
    .a(1'b0),
    .b(sum_10[55]),
    .c(cout_11[54]),
    .cout(cout_11[55]),
    .sum(sum_11[55]));
  AL_FADD comp11_56 (
    .a(1'b0),
    .b(sum_10[56]),
    .c(cout_11[55]),
    .cout(cout_11[56]),
    .sum(sum_11[56]));
  AL_FADD comp11_57 (
    .a(1'b0),
    .b(sum_10[57]),
    .c(cout_11[56]),
    .cout(cout_11[57]),
    .sum(sum_11[57]));
  AL_FADD comp11_58 (
    .a(1'b0),
    .b(sum_10[58]),
    .c(cout_11[57]),
    .cout(cout_11[58]),
    .sum(sum_11[58]));
  AL_FADD comp11_59 (
    .a(1'b0),
    .b(sum_10[59]),
    .c(cout_11[58]),
    .cout(cout_11[59]),
    .sum(sum_11[59]));
  AL_FADD comp11_6 (
    .a(i11[6]),
    .b(sum_10[6]),
    .c(cout_11[5]),
    .cout(cout_11[6]),
    .sum(sum_11[6]));
  AL_FADD comp11_60 (
    .a(1'b0),
    .b(sum_10[60]),
    .c(cout_11[59]),
    .cout(cout_11[60]),
    .sum(sum_11[60]));
  AL_FADD comp11_61 (
    .a(1'b0),
    .b(sum_10[61]),
    .c(cout_11[60]),
    .cout(cout_11[61]),
    .sum(sum_11[61]));
  AL_FADD comp11_62 (
    .a(1'b0),
    .b(sum_10[62]),
    .c(cout_11[61]),
    .cout(cout_11[62]),
    .sum(sum_11[62]));
  AL_FADD comp11_63 (
    .a(1'b0),
    .b(sum_10[63]),
    .c(cout_11[62]),
    .cout(cout_11[63]),
    .sum(sum_11[63]));
  AL_FADD comp11_7 (
    .a(i11[7]),
    .b(sum_10[7]),
    .c(cout_11[6]),
    .cout(cout_11[7]),
    .sum(sum_11[7]));
  AL_FADD comp11_8 (
    .a(i11[8]),
    .b(sum_10[8]),
    .c(cout_11[7]),
    .cout(cout_11[8]),
    .sum(sum_11[8]));
  AL_FADD comp11_9 (
    .a(i11[9]),
    .b(sum_10[9]),
    .c(cout_11[8]),
    .cout(cout_11[9]),
    .sum(sum_11[9]));
  AL_FADD comp12_0 (
    .a(i12[0]),
    .b(sum_11[0]),
    .c(1'b0),
    .cout(cout_12[0]),
    .sum(sum_12[0]));
  AL_FADD comp12_1 (
    .a(i12[1]),
    .b(sum_11[1]),
    .c(cout_12[0]),
    .cout(cout_12[1]),
    .sum(sum_12[1]));
  AL_FADD comp12_10 (
    .a(i12[10]),
    .b(sum_11[10]),
    .c(cout_12[9]),
    .cout(cout_12[10]),
    .sum(sum_12[10]));
  AL_FADD comp12_11 (
    .a(i12[11]),
    .b(sum_11[11]),
    .c(cout_12[10]),
    .cout(cout_12[11]),
    .sum(sum_12[11]));
  AL_FADD comp12_12 (
    .a(i12[12]),
    .b(sum_11[12]),
    .c(cout_12[11]),
    .cout(cout_12[12]),
    .sum(sum_12[12]));
  AL_FADD comp12_13 (
    .a(i12[13]),
    .b(sum_11[13]),
    .c(cout_12[12]),
    .cout(cout_12[13]),
    .sum(sum_12[13]));
  AL_FADD comp12_14 (
    .a(i12[14]),
    .b(sum_11[14]),
    .c(cout_12[13]),
    .cout(cout_12[14]),
    .sum(sum_12[14]));
  AL_FADD comp12_15 (
    .a(i12[15]),
    .b(sum_11[15]),
    .c(cout_12[14]),
    .cout(cout_12[15]),
    .sum(sum_12[15]));
  AL_FADD comp12_16 (
    .a(i12[16]),
    .b(sum_11[16]),
    .c(cout_12[15]),
    .cout(cout_12[16]),
    .sum(sum_12[16]));
  AL_FADD comp12_17 (
    .a(i12[17]),
    .b(sum_11[17]),
    .c(cout_12[16]),
    .cout(cout_12[17]),
    .sum(sum_12[17]));
  AL_FADD comp12_18 (
    .a(i12[18]),
    .b(sum_11[18]),
    .c(cout_12[17]),
    .cout(cout_12[18]),
    .sum(sum_12[18]));
  AL_FADD comp12_19 (
    .a(i12[19]),
    .b(sum_11[19]),
    .c(cout_12[18]),
    .cout(cout_12[19]),
    .sum(sum_12[19]));
  AL_FADD comp12_2 (
    .a(i12[2]),
    .b(sum_11[2]),
    .c(cout_12[1]),
    .cout(cout_12[2]),
    .sum(sum_12[2]));
  AL_FADD comp12_20 (
    .a(i12[20]),
    .b(sum_11[20]),
    .c(cout_12[19]),
    .cout(cout_12[20]),
    .sum(sum_12[20]));
  AL_FADD comp12_21 (
    .a(i12[21]),
    .b(sum_11[21]),
    .c(cout_12[20]),
    .cout(cout_12[21]),
    .sum(sum_12[21]));
  AL_FADD comp12_22 (
    .a(i12[22]),
    .b(sum_11[22]),
    .c(cout_12[21]),
    .cout(cout_12[22]),
    .sum(sum_12[22]));
  AL_FADD comp12_23 (
    .a(i12[23]),
    .b(sum_11[23]),
    .c(cout_12[22]),
    .cout(cout_12[23]),
    .sum(sum_12[23]));
  AL_FADD comp12_24 (
    .a(i12[24]),
    .b(sum_11[24]),
    .c(cout_12[23]),
    .cout(cout_12[24]),
    .sum(sum_12[24]));
  AL_FADD comp12_25 (
    .a(i12[25]),
    .b(sum_11[25]),
    .c(cout_12[24]),
    .cout(cout_12[25]),
    .sum(sum_12[25]));
  AL_FADD comp12_26 (
    .a(i12[26]),
    .b(sum_11[26]),
    .c(cout_12[25]),
    .cout(cout_12[26]),
    .sum(sum_12[26]));
  AL_FADD comp12_27 (
    .a(i12[27]),
    .b(sum_11[27]),
    .c(cout_12[26]),
    .cout(cout_12[27]),
    .sum(sum_12[27]));
  AL_FADD comp12_28 (
    .a(i12[28]),
    .b(sum_11[28]),
    .c(cout_12[27]),
    .cout(cout_12[28]),
    .sum(sum_12[28]));
  AL_FADD comp12_29 (
    .a(i12[29]),
    .b(sum_11[29]),
    .c(cout_12[28]),
    .cout(cout_12[29]),
    .sum(sum_12[29]));
  AL_FADD comp12_3 (
    .a(i12[3]),
    .b(sum_11[3]),
    .c(cout_12[2]),
    .cout(cout_12[3]),
    .sum(sum_12[3]));
  AL_FADD comp12_30 (
    .a(i12[30]),
    .b(sum_11[30]),
    .c(cout_12[29]),
    .cout(cout_12[30]),
    .sum(sum_12[30]));
  AL_FADD comp12_31 (
    .a(i12[31]),
    .b(sum_11[31]),
    .c(cout_12[30]),
    .cout(cout_12[31]),
    .sum(sum_12[31]));
  AL_FADD comp12_32 (
    .a(i12[32]),
    .b(sum_11[32]),
    .c(cout_12[31]),
    .cout(cout_12[32]),
    .sum(sum_12[32]));
  AL_FADD comp12_33 (
    .a(i12[33]),
    .b(sum_11[33]),
    .c(cout_12[32]),
    .cout(cout_12[33]),
    .sum(sum_12[33]));
  AL_FADD comp12_34 (
    .a(i12[34]),
    .b(sum_11[34]),
    .c(cout_12[33]),
    .cout(cout_12[34]),
    .sum(sum_12[34]));
  AL_FADD comp12_35 (
    .a(i12[35]),
    .b(sum_11[35]),
    .c(cout_12[34]),
    .cout(cout_12[35]),
    .sum(sum_12[35]));
  AL_FADD comp12_36 (
    .a(i12[36]),
    .b(sum_11[36]),
    .c(cout_12[35]),
    .cout(cout_12[36]),
    .sum(sum_12[36]));
  AL_FADD comp12_37 (
    .a(i12[37]),
    .b(sum_11[37]),
    .c(cout_12[36]),
    .cout(cout_12[37]),
    .sum(sum_12[37]));
  AL_FADD comp12_38 (
    .a(i12[38]),
    .b(sum_11[38]),
    .c(cout_12[37]),
    .cout(cout_12[38]),
    .sum(sum_12[38]));
  AL_FADD comp12_39 (
    .a(i12[39]),
    .b(sum_11[39]),
    .c(cout_12[38]),
    .cout(cout_12[39]),
    .sum(sum_12[39]));
  AL_FADD comp12_4 (
    .a(i12[4]),
    .b(sum_11[4]),
    .c(cout_12[3]),
    .cout(cout_12[4]),
    .sum(sum_12[4]));
  AL_FADD comp12_40 (
    .a(i12[40]),
    .b(sum_11[40]),
    .c(cout_12[39]),
    .cout(cout_12[40]),
    .sum(sum_12[40]));
  AL_FADD comp12_41 (
    .a(i12[41]),
    .b(sum_11[41]),
    .c(cout_12[40]),
    .cout(cout_12[41]),
    .sum(sum_12[41]));
  AL_FADD comp12_42 (
    .a(i12[42]),
    .b(sum_11[42]),
    .c(cout_12[41]),
    .cout(cout_12[42]),
    .sum(sum_12[42]));
  AL_FADD comp12_43 (
    .a(i12[43]),
    .b(sum_11[43]),
    .c(cout_12[42]),
    .cout(cout_12[43]),
    .sum(sum_12[43]));
  AL_FADD comp12_44 (
    .a(i12[44]),
    .b(sum_11[44]),
    .c(cout_12[43]),
    .cout(cout_12[44]),
    .sum(sum_12[44]));
  AL_FADD comp12_45 (
    .a(i12[45]),
    .b(sum_11[45]),
    .c(cout_12[44]),
    .cout(cout_12[45]),
    .sum(sum_12[45]));
  AL_FADD comp12_46 (
    .a(i12[46]),
    .b(sum_11[46]),
    .c(cout_12[45]),
    .cout(cout_12[46]),
    .sum(sum_12[46]));
  AL_FADD comp12_47 (
    .a(i12[47]),
    .b(sum_11[47]),
    .c(cout_12[46]),
    .cout(cout_12[47]),
    .sum(sum_12[47]));
  AL_FADD comp12_48 (
    .a(i12[48]),
    .b(sum_11[48]),
    .c(cout_12[47]),
    .cout(cout_12[48]),
    .sum(sum_12[48]));
  AL_FADD comp12_49 (
    .a(1'b0),
    .b(sum_11[49]),
    .c(cout_12[48]),
    .cout(cout_12[49]),
    .sum(sum_12[49]));
  AL_FADD comp12_5 (
    .a(i12[5]),
    .b(sum_11[5]),
    .c(cout_12[4]),
    .cout(cout_12[5]),
    .sum(sum_12[5]));
  AL_FADD comp12_50 (
    .a(1'b0),
    .b(sum_11[50]),
    .c(cout_12[49]),
    .cout(cout_12[50]),
    .sum(sum_12[50]));
  AL_FADD comp12_51 (
    .a(1'b0),
    .b(sum_11[51]),
    .c(cout_12[50]),
    .cout(cout_12[51]),
    .sum(sum_12[51]));
  AL_FADD comp12_52 (
    .a(1'b0),
    .b(sum_11[52]),
    .c(cout_12[51]),
    .cout(cout_12[52]),
    .sum(sum_12[52]));
  AL_FADD comp12_53 (
    .a(1'b0),
    .b(sum_11[53]),
    .c(cout_12[52]),
    .cout(cout_12[53]),
    .sum(sum_12[53]));
  AL_FADD comp12_54 (
    .a(1'b0),
    .b(sum_11[54]),
    .c(cout_12[53]),
    .cout(cout_12[54]),
    .sum(sum_12[54]));
  AL_FADD comp12_55 (
    .a(1'b0),
    .b(sum_11[55]),
    .c(cout_12[54]),
    .cout(cout_12[55]),
    .sum(sum_12[55]));
  AL_FADD comp12_56 (
    .a(1'b0),
    .b(sum_11[56]),
    .c(cout_12[55]),
    .cout(cout_12[56]),
    .sum(sum_12[56]));
  AL_FADD comp12_57 (
    .a(1'b0),
    .b(sum_11[57]),
    .c(cout_12[56]),
    .cout(cout_12[57]),
    .sum(sum_12[57]));
  AL_FADD comp12_58 (
    .a(1'b0),
    .b(sum_11[58]),
    .c(cout_12[57]),
    .cout(cout_12[58]),
    .sum(sum_12[58]));
  AL_FADD comp12_59 (
    .a(1'b0),
    .b(sum_11[59]),
    .c(cout_12[58]),
    .cout(cout_12[59]),
    .sum(sum_12[59]));
  AL_FADD comp12_6 (
    .a(i12[6]),
    .b(sum_11[6]),
    .c(cout_12[5]),
    .cout(cout_12[6]),
    .sum(sum_12[6]));
  AL_FADD comp12_60 (
    .a(1'b0),
    .b(sum_11[60]),
    .c(cout_12[59]),
    .cout(cout_12[60]),
    .sum(sum_12[60]));
  AL_FADD comp12_61 (
    .a(1'b0),
    .b(sum_11[61]),
    .c(cout_12[60]),
    .cout(cout_12[61]),
    .sum(sum_12[61]));
  AL_FADD comp12_62 (
    .a(1'b0),
    .b(sum_11[62]),
    .c(cout_12[61]),
    .cout(cout_12[62]),
    .sum(sum_12[62]));
  AL_FADD comp12_63 (
    .a(1'b0),
    .b(sum_11[63]),
    .c(cout_12[62]),
    .cout(cout_12[63]),
    .sum(sum_12[63]));
  AL_FADD comp12_7 (
    .a(i12[7]),
    .b(sum_11[7]),
    .c(cout_12[6]),
    .cout(cout_12[7]),
    .sum(sum_12[7]));
  AL_FADD comp12_8 (
    .a(i12[8]),
    .b(sum_11[8]),
    .c(cout_12[7]),
    .cout(cout_12[8]),
    .sum(sum_12[8]));
  AL_FADD comp12_9 (
    .a(i12[9]),
    .b(sum_11[9]),
    .c(cout_12[8]),
    .cout(cout_12[9]),
    .sum(sum_12[9]));
  AL_FADD comp13_0 (
    .a(i13[0]),
    .b(sum_12[0]),
    .c(1'b0),
    .cout(cout_13[0]),
    .sum(sum_13[0]));
  AL_FADD comp13_1 (
    .a(i13[1]),
    .b(sum_12[1]),
    .c(cout_13[0]),
    .cout(cout_13[1]),
    .sum(sum_13[1]));
  AL_FADD comp13_10 (
    .a(i13[10]),
    .b(sum_12[10]),
    .c(cout_13[9]),
    .cout(cout_13[10]),
    .sum(sum_13[10]));
  AL_FADD comp13_11 (
    .a(i13[11]),
    .b(sum_12[11]),
    .c(cout_13[10]),
    .cout(cout_13[11]),
    .sum(sum_13[11]));
  AL_FADD comp13_12 (
    .a(i13[12]),
    .b(sum_12[12]),
    .c(cout_13[11]),
    .cout(cout_13[12]),
    .sum(sum_13[12]));
  AL_FADD comp13_13 (
    .a(i13[13]),
    .b(sum_12[13]),
    .c(cout_13[12]),
    .cout(cout_13[13]),
    .sum(sum_13[13]));
  AL_FADD comp13_14 (
    .a(i13[14]),
    .b(sum_12[14]),
    .c(cout_13[13]),
    .cout(cout_13[14]),
    .sum(sum_13[14]));
  AL_FADD comp13_15 (
    .a(i13[15]),
    .b(sum_12[15]),
    .c(cout_13[14]),
    .cout(cout_13[15]),
    .sum(sum_13[15]));
  AL_FADD comp13_16 (
    .a(i13[16]),
    .b(sum_12[16]),
    .c(cout_13[15]),
    .cout(cout_13[16]),
    .sum(sum_13[16]));
  AL_FADD comp13_17 (
    .a(i13[17]),
    .b(sum_12[17]),
    .c(cout_13[16]),
    .cout(cout_13[17]),
    .sum(sum_13[17]));
  AL_FADD comp13_18 (
    .a(i13[18]),
    .b(sum_12[18]),
    .c(cout_13[17]),
    .cout(cout_13[18]),
    .sum(sum_13[18]));
  AL_FADD comp13_19 (
    .a(i13[19]),
    .b(sum_12[19]),
    .c(cout_13[18]),
    .cout(cout_13[19]),
    .sum(sum_13[19]));
  AL_FADD comp13_2 (
    .a(i13[2]),
    .b(sum_12[2]),
    .c(cout_13[1]),
    .cout(cout_13[2]),
    .sum(sum_13[2]));
  AL_FADD comp13_20 (
    .a(i13[20]),
    .b(sum_12[20]),
    .c(cout_13[19]),
    .cout(cout_13[20]),
    .sum(sum_13[20]));
  AL_FADD comp13_21 (
    .a(i13[21]),
    .b(sum_12[21]),
    .c(cout_13[20]),
    .cout(cout_13[21]),
    .sum(sum_13[21]));
  AL_FADD comp13_22 (
    .a(i13[22]),
    .b(sum_12[22]),
    .c(cout_13[21]),
    .cout(cout_13[22]),
    .sum(sum_13[22]));
  AL_FADD comp13_23 (
    .a(i13[23]),
    .b(sum_12[23]),
    .c(cout_13[22]),
    .cout(cout_13[23]),
    .sum(sum_13[23]));
  AL_FADD comp13_24 (
    .a(i13[24]),
    .b(sum_12[24]),
    .c(cout_13[23]),
    .cout(cout_13[24]),
    .sum(sum_13[24]));
  AL_FADD comp13_25 (
    .a(i13[25]),
    .b(sum_12[25]),
    .c(cout_13[24]),
    .cout(cout_13[25]),
    .sum(sum_13[25]));
  AL_FADD comp13_26 (
    .a(i13[26]),
    .b(sum_12[26]),
    .c(cout_13[25]),
    .cout(cout_13[26]),
    .sum(sum_13[26]));
  AL_FADD comp13_27 (
    .a(i13[27]),
    .b(sum_12[27]),
    .c(cout_13[26]),
    .cout(cout_13[27]),
    .sum(sum_13[27]));
  AL_FADD comp13_28 (
    .a(i13[28]),
    .b(sum_12[28]),
    .c(cout_13[27]),
    .cout(cout_13[28]),
    .sum(sum_13[28]));
  AL_FADD comp13_29 (
    .a(i13[29]),
    .b(sum_12[29]),
    .c(cout_13[28]),
    .cout(cout_13[29]),
    .sum(sum_13[29]));
  AL_FADD comp13_3 (
    .a(i13[3]),
    .b(sum_12[3]),
    .c(cout_13[2]),
    .cout(cout_13[3]),
    .sum(sum_13[3]));
  AL_FADD comp13_30 (
    .a(i13[30]),
    .b(sum_12[30]),
    .c(cout_13[29]),
    .cout(cout_13[30]),
    .sum(sum_13[30]));
  AL_FADD comp13_31 (
    .a(i13[31]),
    .b(sum_12[31]),
    .c(cout_13[30]),
    .cout(cout_13[31]),
    .sum(sum_13[31]));
  AL_FADD comp13_32 (
    .a(i13[32]),
    .b(sum_12[32]),
    .c(cout_13[31]),
    .cout(cout_13[32]),
    .sum(sum_13[32]));
  AL_FADD comp13_33 (
    .a(i13[33]),
    .b(sum_12[33]),
    .c(cout_13[32]),
    .cout(cout_13[33]),
    .sum(sum_13[33]));
  AL_FADD comp13_34 (
    .a(i13[34]),
    .b(sum_12[34]),
    .c(cout_13[33]),
    .cout(cout_13[34]),
    .sum(sum_13[34]));
  AL_FADD comp13_35 (
    .a(i13[35]),
    .b(sum_12[35]),
    .c(cout_13[34]),
    .cout(cout_13[35]),
    .sum(sum_13[35]));
  AL_FADD comp13_36 (
    .a(i13[36]),
    .b(sum_12[36]),
    .c(cout_13[35]),
    .cout(cout_13[36]),
    .sum(sum_13[36]));
  AL_FADD comp13_37 (
    .a(i13[37]),
    .b(sum_12[37]),
    .c(cout_13[36]),
    .cout(cout_13[37]),
    .sum(sum_13[37]));
  AL_FADD comp13_38 (
    .a(i13[38]),
    .b(sum_12[38]),
    .c(cout_13[37]),
    .cout(cout_13[38]),
    .sum(sum_13[38]));
  AL_FADD comp13_39 (
    .a(i13[39]),
    .b(sum_12[39]),
    .c(cout_13[38]),
    .cout(cout_13[39]),
    .sum(sum_13[39]));
  AL_FADD comp13_4 (
    .a(i13[4]),
    .b(sum_12[4]),
    .c(cout_13[3]),
    .cout(cout_13[4]),
    .sum(sum_13[4]));
  AL_FADD comp13_40 (
    .a(i13[40]),
    .b(sum_12[40]),
    .c(cout_13[39]),
    .cout(cout_13[40]),
    .sum(sum_13[40]));
  AL_FADD comp13_41 (
    .a(i13[41]),
    .b(sum_12[41]),
    .c(cout_13[40]),
    .cout(cout_13[41]),
    .sum(sum_13[41]));
  AL_FADD comp13_42 (
    .a(i13[42]),
    .b(sum_12[42]),
    .c(cout_13[41]),
    .cout(cout_13[42]),
    .sum(sum_13[42]));
  AL_FADD comp13_43 (
    .a(i13[43]),
    .b(sum_12[43]),
    .c(cout_13[42]),
    .cout(cout_13[43]),
    .sum(sum_13[43]));
  AL_FADD comp13_44 (
    .a(i13[44]),
    .b(sum_12[44]),
    .c(cout_13[43]),
    .cout(cout_13[44]),
    .sum(sum_13[44]));
  AL_FADD comp13_45 (
    .a(i13[45]),
    .b(sum_12[45]),
    .c(cout_13[44]),
    .cout(cout_13[45]),
    .sum(sum_13[45]));
  AL_FADD comp13_46 (
    .a(i13[46]),
    .b(sum_12[46]),
    .c(cout_13[45]),
    .cout(cout_13[46]),
    .sum(sum_13[46]));
  AL_FADD comp13_47 (
    .a(i13[47]),
    .b(sum_12[47]),
    .c(cout_13[46]),
    .cout(cout_13[47]),
    .sum(sum_13[47]));
  AL_FADD comp13_48 (
    .a(1'b0),
    .b(sum_12[48]),
    .c(cout_13[47]),
    .cout(cout_13[48]),
    .sum(sum_13[48]));
  AL_FADD comp13_49 (
    .a(1'b0),
    .b(sum_12[49]),
    .c(cout_13[48]),
    .cout(cout_13[49]),
    .sum(sum_13[49]));
  AL_FADD comp13_5 (
    .a(i13[5]),
    .b(sum_12[5]),
    .c(cout_13[4]),
    .cout(cout_13[5]),
    .sum(sum_13[5]));
  AL_FADD comp13_50 (
    .a(1'b0),
    .b(sum_12[50]),
    .c(cout_13[49]),
    .cout(cout_13[50]),
    .sum(sum_13[50]));
  AL_FADD comp13_51 (
    .a(1'b0),
    .b(sum_12[51]),
    .c(cout_13[50]),
    .cout(cout_13[51]),
    .sum(sum_13[51]));
  AL_FADD comp13_52 (
    .a(1'b0),
    .b(sum_12[52]),
    .c(cout_13[51]),
    .cout(cout_13[52]),
    .sum(sum_13[52]));
  AL_FADD comp13_53 (
    .a(1'b0),
    .b(sum_12[53]),
    .c(cout_13[52]),
    .cout(cout_13[53]),
    .sum(sum_13[53]));
  AL_FADD comp13_54 (
    .a(1'b0),
    .b(sum_12[54]),
    .c(cout_13[53]),
    .cout(cout_13[54]),
    .sum(sum_13[54]));
  AL_FADD comp13_55 (
    .a(1'b0),
    .b(sum_12[55]),
    .c(cout_13[54]),
    .cout(cout_13[55]),
    .sum(sum_13[55]));
  AL_FADD comp13_56 (
    .a(1'b0),
    .b(sum_12[56]),
    .c(cout_13[55]),
    .cout(cout_13[56]),
    .sum(sum_13[56]));
  AL_FADD comp13_57 (
    .a(1'b0),
    .b(sum_12[57]),
    .c(cout_13[56]),
    .cout(cout_13[57]),
    .sum(sum_13[57]));
  AL_FADD comp13_58 (
    .a(1'b0),
    .b(sum_12[58]),
    .c(cout_13[57]),
    .cout(cout_13[58]),
    .sum(sum_13[58]));
  AL_FADD comp13_59 (
    .a(1'b0),
    .b(sum_12[59]),
    .c(cout_13[58]),
    .cout(cout_13[59]),
    .sum(sum_13[59]));
  AL_FADD comp13_6 (
    .a(i13[6]),
    .b(sum_12[6]),
    .c(cout_13[5]),
    .cout(cout_13[6]),
    .sum(sum_13[6]));
  AL_FADD comp13_60 (
    .a(1'b0),
    .b(sum_12[60]),
    .c(cout_13[59]),
    .cout(cout_13[60]),
    .sum(sum_13[60]));
  AL_FADD comp13_61 (
    .a(1'b0),
    .b(sum_12[61]),
    .c(cout_13[60]),
    .cout(cout_13[61]),
    .sum(sum_13[61]));
  AL_FADD comp13_62 (
    .a(1'b0),
    .b(sum_12[62]),
    .c(cout_13[61]),
    .cout(cout_13[62]),
    .sum(sum_13[62]));
  AL_FADD comp13_63 (
    .a(1'b0),
    .b(sum_12[63]),
    .c(cout_13[62]),
    .cout(cout_13[63]),
    .sum(sum_13[63]));
  AL_FADD comp13_7 (
    .a(i13[7]),
    .b(sum_12[7]),
    .c(cout_13[6]),
    .cout(cout_13[7]),
    .sum(sum_13[7]));
  AL_FADD comp13_8 (
    .a(i13[8]),
    .b(sum_12[8]),
    .c(cout_13[7]),
    .cout(cout_13[8]),
    .sum(sum_13[8]));
  AL_FADD comp13_9 (
    .a(i13[9]),
    .b(sum_12[9]),
    .c(cout_13[8]),
    .cout(cout_13[9]),
    .sum(sum_13[9]));
  AL_FADD comp14_0 (
    .a(i14[0]),
    .b(sum_13[0]),
    .c(1'b0),
    .cout(cout_14[0]),
    .sum(sum_14[0]));
  AL_FADD comp14_1 (
    .a(i14[1]),
    .b(sum_13[1]),
    .c(cout_14[0]),
    .cout(cout_14[1]),
    .sum(sum_14[1]));
  AL_FADD comp14_10 (
    .a(i14[10]),
    .b(sum_13[10]),
    .c(cout_14[9]),
    .cout(cout_14[10]),
    .sum(sum_14[10]));
  AL_FADD comp14_11 (
    .a(i14[11]),
    .b(sum_13[11]),
    .c(cout_14[10]),
    .cout(cout_14[11]),
    .sum(sum_14[11]));
  AL_FADD comp14_12 (
    .a(i14[12]),
    .b(sum_13[12]),
    .c(cout_14[11]),
    .cout(cout_14[12]),
    .sum(sum_14[12]));
  AL_FADD comp14_13 (
    .a(i14[13]),
    .b(sum_13[13]),
    .c(cout_14[12]),
    .cout(cout_14[13]),
    .sum(sum_14[13]));
  AL_FADD comp14_14 (
    .a(i14[14]),
    .b(sum_13[14]),
    .c(cout_14[13]),
    .cout(cout_14[14]),
    .sum(sum_14[14]));
  AL_FADD comp14_15 (
    .a(i14[15]),
    .b(sum_13[15]),
    .c(cout_14[14]),
    .cout(cout_14[15]),
    .sum(sum_14[15]));
  AL_FADD comp14_16 (
    .a(i14[16]),
    .b(sum_13[16]),
    .c(cout_14[15]),
    .cout(cout_14[16]),
    .sum(sum_14[16]));
  AL_FADD comp14_17 (
    .a(i14[17]),
    .b(sum_13[17]),
    .c(cout_14[16]),
    .cout(cout_14[17]),
    .sum(sum_14[17]));
  AL_FADD comp14_18 (
    .a(i14[18]),
    .b(sum_13[18]),
    .c(cout_14[17]),
    .cout(cout_14[18]),
    .sum(sum_14[18]));
  AL_FADD comp14_19 (
    .a(i14[19]),
    .b(sum_13[19]),
    .c(cout_14[18]),
    .cout(cout_14[19]),
    .sum(sum_14[19]));
  AL_FADD comp14_2 (
    .a(i14[2]),
    .b(sum_13[2]),
    .c(cout_14[1]),
    .cout(cout_14[2]),
    .sum(sum_14[2]));
  AL_FADD comp14_20 (
    .a(i14[20]),
    .b(sum_13[20]),
    .c(cout_14[19]),
    .cout(cout_14[20]),
    .sum(sum_14[20]));
  AL_FADD comp14_21 (
    .a(i14[21]),
    .b(sum_13[21]),
    .c(cout_14[20]),
    .cout(cout_14[21]),
    .sum(sum_14[21]));
  AL_FADD comp14_22 (
    .a(i14[22]),
    .b(sum_13[22]),
    .c(cout_14[21]),
    .cout(cout_14[22]),
    .sum(sum_14[22]));
  AL_FADD comp14_23 (
    .a(i14[23]),
    .b(sum_13[23]),
    .c(cout_14[22]),
    .cout(cout_14[23]),
    .sum(sum_14[23]));
  AL_FADD comp14_24 (
    .a(i14[24]),
    .b(sum_13[24]),
    .c(cout_14[23]),
    .cout(cout_14[24]),
    .sum(sum_14[24]));
  AL_FADD comp14_25 (
    .a(i14[25]),
    .b(sum_13[25]),
    .c(cout_14[24]),
    .cout(cout_14[25]),
    .sum(sum_14[25]));
  AL_FADD comp14_26 (
    .a(i14[26]),
    .b(sum_13[26]),
    .c(cout_14[25]),
    .cout(cout_14[26]),
    .sum(sum_14[26]));
  AL_FADD comp14_27 (
    .a(i14[27]),
    .b(sum_13[27]),
    .c(cout_14[26]),
    .cout(cout_14[27]),
    .sum(sum_14[27]));
  AL_FADD comp14_28 (
    .a(i14[28]),
    .b(sum_13[28]),
    .c(cout_14[27]),
    .cout(cout_14[28]),
    .sum(sum_14[28]));
  AL_FADD comp14_29 (
    .a(i14[29]),
    .b(sum_13[29]),
    .c(cout_14[28]),
    .cout(cout_14[29]),
    .sum(sum_14[29]));
  AL_FADD comp14_3 (
    .a(i14[3]),
    .b(sum_13[3]),
    .c(cout_14[2]),
    .cout(cout_14[3]),
    .sum(sum_14[3]));
  AL_FADD comp14_30 (
    .a(i14[30]),
    .b(sum_13[30]),
    .c(cout_14[29]),
    .cout(cout_14[30]),
    .sum(sum_14[30]));
  AL_FADD comp14_31 (
    .a(i14[31]),
    .b(sum_13[31]),
    .c(cout_14[30]),
    .cout(cout_14[31]),
    .sum(sum_14[31]));
  AL_FADD comp14_32 (
    .a(i14[32]),
    .b(sum_13[32]),
    .c(cout_14[31]),
    .cout(cout_14[32]),
    .sum(sum_14[32]));
  AL_FADD comp14_33 (
    .a(i14[33]),
    .b(sum_13[33]),
    .c(cout_14[32]),
    .cout(cout_14[33]),
    .sum(sum_14[33]));
  AL_FADD comp14_34 (
    .a(i14[34]),
    .b(sum_13[34]),
    .c(cout_14[33]),
    .cout(cout_14[34]),
    .sum(sum_14[34]));
  AL_FADD comp14_35 (
    .a(i14[35]),
    .b(sum_13[35]),
    .c(cout_14[34]),
    .cout(cout_14[35]),
    .sum(sum_14[35]));
  AL_FADD comp14_36 (
    .a(i14[36]),
    .b(sum_13[36]),
    .c(cout_14[35]),
    .cout(cout_14[36]),
    .sum(sum_14[36]));
  AL_FADD comp14_37 (
    .a(i14[37]),
    .b(sum_13[37]),
    .c(cout_14[36]),
    .cout(cout_14[37]),
    .sum(sum_14[37]));
  AL_FADD comp14_38 (
    .a(i14[38]),
    .b(sum_13[38]),
    .c(cout_14[37]),
    .cout(cout_14[38]),
    .sum(sum_14[38]));
  AL_FADD comp14_39 (
    .a(i14[39]),
    .b(sum_13[39]),
    .c(cout_14[38]),
    .cout(cout_14[39]),
    .sum(sum_14[39]));
  AL_FADD comp14_4 (
    .a(i14[4]),
    .b(sum_13[4]),
    .c(cout_14[3]),
    .cout(cout_14[4]),
    .sum(sum_14[4]));
  AL_FADD comp14_40 (
    .a(i14[40]),
    .b(sum_13[40]),
    .c(cout_14[39]),
    .cout(cout_14[40]),
    .sum(sum_14[40]));
  AL_FADD comp14_41 (
    .a(i14[41]),
    .b(sum_13[41]),
    .c(cout_14[40]),
    .cout(cout_14[41]),
    .sum(sum_14[41]));
  AL_FADD comp14_42 (
    .a(i14[42]),
    .b(sum_13[42]),
    .c(cout_14[41]),
    .cout(cout_14[42]),
    .sum(sum_14[42]));
  AL_FADD comp14_43 (
    .a(i14[43]),
    .b(sum_13[43]),
    .c(cout_14[42]),
    .cout(cout_14[43]),
    .sum(sum_14[43]));
  AL_FADD comp14_44 (
    .a(i14[44]),
    .b(sum_13[44]),
    .c(cout_14[43]),
    .cout(cout_14[44]),
    .sum(sum_14[44]));
  AL_FADD comp14_45 (
    .a(i14[45]),
    .b(sum_13[45]),
    .c(cout_14[44]),
    .cout(cout_14[45]),
    .sum(sum_14[45]));
  AL_FADD comp14_46 (
    .a(i14[46]),
    .b(sum_13[46]),
    .c(cout_14[45]),
    .cout(cout_14[46]),
    .sum(sum_14[46]));
  AL_FADD comp14_47 (
    .a(1'b0),
    .b(sum_13[47]),
    .c(cout_14[46]),
    .cout(cout_14[47]),
    .sum(sum_14[47]));
  AL_FADD comp14_48 (
    .a(1'b0),
    .b(sum_13[48]),
    .c(cout_14[47]),
    .cout(cout_14[48]),
    .sum(sum_14[48]));
  AL_FADD comp14_49 (
    .a(1'b0),
    .b(sum_13[49]),
    .c(cout_14[48]),
    .cout(cout_14[49]),
    .sum(sum_14[49]));
  AL_FADD comp14_5 (
    .a(i14[5]),
    .b(sum_13[5]),
    .c(cout_14[4]),
    .cout(cout_14[5]),
    .sum(sum_14[5]));
  AL_FADD comp14_50 (
    .a(1'b0),
    .b(sum_13[50]),
    .c(cout_14[49]),
    .cout(cout_14[50]),
    .sum(sum_14[50]));
  AL_FADD comp14_51 (
    .a(1'b0),
    .b(sum_13[51]),
    .c(cout_14[50]),
    .cout(cout_14[51]),
    .sum(sum_14[51]));
  AL_FADD comp14_52 (
    .a(1'b0),
    .b(sum_13[52]),
    .c(cout_14[51]),
    .cout(cout_14[52]),
    .sum(sum_14[52]));
  AL_FADD comp14_53 (
    .a(1'b0),
    .b(sum_13[53]),
    .c(cout_14[52]),
    .cout(cout_14[53]),
    .sum(sum_14[53]));
  AL_FADD comp14_54 (
    .a(1'b0),
    .b(sum_13[54]),
    .c(cout_14[53]),
    .cout(cout_14[54]),
    .sum(sum_14[54]));
  AL_FADD comp14_55 (
    .a(1'b0),
    .b(sum_13[55]),
    .c(cout_14[54]),
    .cout(cout_14[55]),
    .sum(sum_14[55]));
  AL_FADD comp14_56 (
    .a(1'b0),
    .b(sum_13[56]),
    .c(cout_14[55]),
    .cout(cout_14[56]),
    .sum(sum_14[56]));
  AL_FADD comp14_57 (
    .a(1'b0),
    .b(sum_13[57]),
    .c(cout_14[56]),
    .cout(cout_14[57]),
    .sum(sum_14[57]));
  AL_FADD comp14_58 (
    .a(1'b0),
    .b(sum_13[58]),
    .c(cout_14[57]),
    .cout(cout_14[58]),
    .sum(sum_14[58]));
  AL_FADD comp14_59 (
    .a(1'b0),
    .b(sum_13[59]),
    .c(cout_14[58]),
    .cout(cout_14[59]),
    .sum(sum_14[59]));
  AL_FADD comp14_6 (
    .a(i14[6]),
    .b(sum_13[6]),
    .c(cout_14[5]),
    .cout(cout_14[6]),
    .sum(sum_14[6]));
  AL_FADD comp14_60 (
    .a(1'b0),
    .b(sum_13[60]),
    .c(cout_14[59]),
    .cout(cout_14[60]),
    .sum(sum_14[60]));
  AL_FADD comp14_61 (
    .a(1'b0),
    .b(sum_13[61]),
    .c(cout_14[60]),
    .cout(cout_14[61]),
    .sum(sum_14[61]));
  AL_FADD comp14_62 (
    .a(1'b0),
    .b(sum_13[62]),
    .c(cout_14[61]),
    .cout(cout_14[62]),
    .sum(sum_14[62]));
  AL_FADD comp14_63 (
    .a(1'b0),
    .b(sum_13[63]),
    .c(cout_14[62]),
    .cout(cout_14[63]),
    .sum(sum_14[63]));
  AL_FADD comp14_7 (
    .a(i14[7]),
    .b(sum_13[7]),
    .c(cout_14[6]),
    .cout(cout_14[7]),
    .sum(sum_14[7]));
  AL_FADD comp14_8 (
    .a(i14[8]),
    .b(sum_13[8]),
    .c(cout_14[7]),
    .cout(cout_14[8]),
    .sum(sum_14[8]));
  AL_FADD comp14_9 (
    .a(i14[9]),
    .b(sum_13[9]),
    .c(cout_14[8]),
    .cout(cout_14[9]),
    .sum(sum_14[9]));
  AL_FADD comp15_0 (
    .a(i15[0]),
    .b(sum_14[0]),
    .c(1'b0),
    .cout(cout_15[0]),
    .sum(sum_15[0]));
  AL_FADD comp15_1 (
    .a(i15[1]),
    .b(sum_14[1]),
    .c(cout_15[0]),
    .cout(cout_15[1]),
    .sum(sum_15[1]));
  AL_FADD comp15_10 (
    .a(i15[10]),
    .b(sum_14[10]),
    .c(cout_15[9]),
    .cout(cout_15[10]),
    .sum(sum_15[10]));
  AL_FADD comp15_11 (
    .a(i15[11]),
    .b(sum_14[11]),
    .c(cout_15[10]),
    .cout(cout_15[11]),
    .sum(sum_15[11]));
  AL_FADD comp15_12 (
    .a(i15[12]),
    .b(sum_14[12]),
    .c(cout_15[11]),
    .cout(cout_15[12]),
    .sum(sum_15[12]));
  AL_FADD comp15_13 (
    .a(i15[13]),
    .b(sum_14[13]),
    .c(cout_15[12]),
    .cout(cout_15[13]),
    .sum(sum_15[13]));
  AL_FADD comp15_14 (
    .a(i15[14]),
    .b(sum_14[14]),
    .c(cout_15[13]),
    .cout(cout_15[14]),
    .sum(sum_15[14]));
  AL_FADD comp15_15 (
    .a(i15[15]),
    .b(sum_14[15]),
    .c(cout_15[14]),
    .cout(cout_15[15]),
    .sum(sum_15[15]));
  AL_FADD comp15_16 (
    .a(i15[16]),
    .b(sum_14[16]),
    .c(cout_15[15]),
    .cout(cout_15[16]),
    .sum(sum_15[16]));
  AL_FADD comp15_17 (
    .a(i15[17]),
    .b(sum_14[17]),
    .c(cout_15[16]),
    .cout(cout_15[17]),
    .sum(sum_15[17]));
  AL_FADD comp15_18 (
    .a(i15[18]),
    .b(sum_14[18]),
    .c(cout_15[17]),
    .cout(cout_15[18]),
    .sum(sum_15[18]));
  AL_FADD comp15_19 (
    .a(i15[19]),
    .b(sum_14[19]),
    .c(cout_15[18]),
    .cout(cout_15[19]),
    .sum(sum_15[19]));
  AL_FADD comp15_2 (
    .a(i15[2]),
    .b(sum_14[2]),
    .c(cout_15[1]),
    .cout(cout_15[2]),
    .sum(sum_15[2]));
  AL_FADD comp15_20 (
    .a(i15[20]),
    .b(sum_14[20]),
    .c(cout_15[19]),
    .cout(cout_15[20]),
    .sum(sum_15[20]));
  AL_FADD comp15_21 (
    .a(i15[21]),
    .b(sum_14[21]),
    .c(cout_15[20]),
    .cout(cout_15[21]),
    .sum(sum_15[21]));
  AL_FADD comp15_22 (
    .a(i15[22]),
    .b(sum_14[22]),
    .c(cout_15[21]),
    .cout(cout_15[22]),
    .sum(sum_15[22]));
  AL_FADD comp15_23 (
    .a(i15[23]),
    .b(sum_14[23]),
    .c(cout_15[22]),
    .cout(cout_15[23]),
    .sum(sum_15[23]));
  AL_FADD comp15_24 (
    .a(i15[24]),
    .b(sum_14[24]),
    .c(cout_15[23]),
    .cout(cout_15[24]),
    .sum(sum_15[24]));
  AL_FADD comp15_25 (
    .a(i15[25]),
    .b(sum_14[25]),
    .c(cout_15[24]),
    .cout(cout_15[25]),
    .sum(sum_15[25]));
  AL_FADD comp15_26 (
    .a(i15[26]),
    .b(sum_14[26]),
    .c(cout_15[25]),
    .cout(cout_15[26]),
    .sum(sum_15[26]));
  AL_FADD comp15_27 (
    .a(i15[27]),
    .b(sum_14[27]),
    .c(cout_15[26]),
    .cout(cout_15[27]),
    .sum(sum_15[27]));
  AL_FADD comp15_28 (
    .a(i15[28]),
    .b(sum_14[28]),
    .c(cout_15[27]),
    .cout(cout_15[28]),
    .sum(sum_15[28]));
  AL_FADD comp15_29 (
    .a(i15[29]),
    .b(sum_14[29]),
    .c(cout_15[28]),
    .cout(cout_15[29]),
    .sum(sum_15[29]));
  AL_FADD comp15_3 (
    .a(i15[3]),
    .b(sum_14[3]),
    .c(cout_15[2]),
    .cout(cout_15[3]),
    .sum(sum_15[3]));
  AL_FADD comp15_30 (
    .a(i15[30]),
    .b(sum_14[30]),
    .c(cout_15[29]),
    .cout(cout_15[30]),
    .sum(sum_15[30]));
  AL_FADD comp15_31 (
    .a(i15[31]),
    .b(sum_14[31]),
    .c(cout_15[30]),
    .cout(cout_15[31]),
    .sum(sum_15[31]));
  AL_FADD comp15_32 (
    .a(i15[32]),
    .b(sum_14[32]),
    .c(cout_15[31]),
    .cout(cout_15[32]),
    .sum(sum_15[32]));
  AL_FADD comp15_33 (
    .a(i15[33]),
    .b(sum_14[33]),
    .c(cout_15[32]),
    .cout(cout_15[33]),
    .sum(sum_15[33]));
  AL_FADD comp15_34 (
    .a(i15[34]),
    .b(sum_14[34]),
    .c(cout_15[33]),
    .cout(cout_15[34]),
    .sum(sum_15[34]));
  AL_FADD comp15_35 (
    .a(i15[35]),
    .b(sum_14[35]),
    .c(cout_15[34]),
    .cout(cout_15[35]),
    .sum(sum_15[35]));
  AL_FADD comp15_36 (
    .a(i15[36]),
    .b(sum_14[36]),
    .c(cout_15[35]),
    .cout(cout_15[36]),
    .sum(sum_15[36]));
  AL_FADD comp15_37 (
    .a(i15[37]),
    .b(sum_14[37]),
    .c(cout_15[36]),
    .cout(cout_15[37]),
    .sum(sum_15[37]));
  AL_FADD comp15_38 (
    .a(i15[38]),
    .b(sum_14[38]),
    .c(cout_15[37]),
    .cout(cout_15[38]),
    .sum(sum_15[38]));
  AL_FADD comp15_39 (
    .a(i15[39]),
    .b(sum_14[39]),
    .c(cout_15[38]),
    .cout(cout_15[39]),
    .sum(sum_15[39]));
  AL_FADD comp15_4 (
    .a(i15[4]),
    .b(sum_14[4]),
    .c(cout_15[3]),
    .cout(cout_15[4]),
    .sum(sum_15[4]));
  AL_FADD comp15_40 (
    .a(i15[40]),
    .b(sum_14[40]),
    .c(cout_15[39]),
    .cout(cout_15[40]),
    .sum(sum_15[40]));
  AL_FADD comp15_41 (
    .a(i15[41]),
    .b(sum_14[41]),
    .c(cout_15[40]),
    .cout(cout_15[41]),
    .sum(sum_15[41]));
  AL_FADD comp15_42 (
    .a(i15[42]),
    .b(sum_14[42]),
    .c(cout_15[41]),
    .cout(cout_15[42]),
    .sum(sum_15[42]));
  AL_FADD comp15_43 (
    .a(i15[43]),
    .b(sum_14[43]),
    .c(cout_15[42]),
    .cout(cout_15[43]),
    .sum(sum_15[43]));
  AL_FADD comp15_44 (
    .a(i15[44]),
    .b(sum_14[44]),
    .c(cout_15[43]),
    .cout(cout_15[44]),
    .sum(sum_15[44]));
  AL_FADD comp15_45 (
    .a(i15[45]),
    .b(sum_14[45]),
    .c(cout_15[44]),
    .cout(cout_15[45]),
    .sum(sum_15[45]));
  AL_FADD comp15_46 (
    .a(1'b0),
    .b(sum_14[46]),
    .c(cout_15[45]),
    .cout(cout_15[46]),
    .sum(sum_15[46]));
  AL_FADD comp15_47 (
    .a(1'b0),
    .b(sum_14[47]),
    .c(cout_15[46]),
    .cout(cout_15[47]),
    .sum(sum_15[47]));
  AL_FADD comp15_48 (
    .a(1'b0),
    .b(sum_14[48]),
    .c(cout_15[47]),
    .cout(cout_15[48]),
    .sum(sum_15[48]));
  AL_FADD comp15_49 (
    .a(1'b0),
    .b(sum_14[49]),
    .c(cout_15[48]),
    .cout(cout_15[49]),
    .sum(sum_15[49]));
  AL_FADD comp15_5 (
    .a(i15[5]),
    .b(sum_14[5]),
    .c(cout_15[4]),
    .cout(cout_15[5]),
    .sum(sum_15[5]));
  AL_FADD comp15_50 (
    .a(1'b0),
    .b(sum_14[50]),
    .c(cout_15[49]),
    .cout(cout_15[50]),
    .sum(sum_15[50]));
  AL_FADD comp15_51 (
    .a(1'b0),
    .b(sum_14[51]),
    .c(cout_15[50]),
    .cout(cout_15[51]),
    .sum(sum_15[51]));
  AL_FADD comp15_52 (
    .a(1'b0),
    .b(sum_14[52]),
    .c(cout_15[51]),
    .cout(cout_15[52]),
    .sum(sum_15[52]));
  AL_FADD comp15_53 (
    .a(1'b0),
    .b(sum_14[53]),
    .c(cout_15[52]),
    .cout(cout_15[53]),
    .sum(sum_15[53]));
  AL_FADD comp15_54 (
    .a(1'b0),
    .b(sum_14[54]),
    .c(cout_15[53]),
    .cout(cout_15[54]),
    .sum(sum_15[54]));
  AL_FADD comp15_55 (
    .a(1'b0),
    .b(sum_14[55]),
    .c(cout_15[54]),
    .cout(cout_15[55]),
    .sum(sum_15[55]));
  AL_FADD comp15_56 (
    .a(1'b0),
    .b(sum_14[56]),
    .c(cout_15[55]),
    .cout(cout_15[56]),
    .sum(sum_15[56]));
  AL_FADD comp15_57 (
    .a(1'b0),
    .b(sum_14[57]),
    .c(cout_15[56]),
    .cout(cout_15[57]),
    .sum(sum_15[57]));
  AL_FADD comp15_58 (
    .a(1'b0),
    .b(sum_14[58]),
    .c(cout_15[57]),
    .cout(cout_15[58]),
    .sum(sum_15[58]));
  AL_FADD comp15_59 (
    .a(1'b0),
    .b(sum_14[59]),
    .c(cout_15[58]),
    .cout(cout_15[59]),
    .sum(sum_15[59]));
  AL_FADD comp15_6 (
    .a(i15[6]),
    .b(sum_14[6]),
    .c(cout_15[5]),
    .cout(cout_15[6]),
    .sum(sum_15[6]));
  AL_FADD comp15_60 (
    .a(1'b0),
    .b(sum_14[60]),
    .c(cout_15[59]),
    .cout(cout_15[60]),
    .sum(sum_15[60]));
  AL_FADD comp15_61 (
    .a(1'b0),
    .b(sum_14[61]),
    .c(cout_15[60]),
    .cout(cout_15[61]),
    .sum(sum_15[61]));
  AL_FADD comp15_62 (
    .a(1'b0),
    .b(sum_14[62]),
    .c(cout_15[61]),
    .cout(cout_15[62]),
    .sum(sum_15[62]));
  AL_FADD comp15_63 (
    .a(1'b0),
    .b(sum_14[63]),
    .c(cout_15[62]),
    .cout(cout_15[63]),
    .sum(sum_15[63]));
  AL_FADD comp15_7 (
    .a(i15[7]),
    .b(sum_14[7]),
    .c(cout_15[6]),
    .cout(cout_15[7]),
    .sum(sum_15[7]));
  AL_FADD comp15_8 (
    .a(i15[8]),
    .b(sum_14[8]),
    .c(cout_15[7]),
    .cout(cout_15[8]),
    .sum(sum_15[8]));
  AL_FADD comp15_9 (
    .a(i15[9]),
    .b(sum_14[9]),
    .c(cout_15[8]),
    .cout(cout_15[9]),
    .sum(sum_15[9]));
  AL_FADD comp16_0 (
    .a(i16[0]),
    .b(sum_15[0]),
    .c(1'b0),
    .cout(cout_16[0]),
    .sum(sum_16[0]));
  AL_FADD comp16_1 (
    .a(i16[1]),
    .b(sum_15[1]),
    .c(cout_16[0]),
    .cout(cout_16[1]),
    .sum(sum_16[1]));
  AL_FADD comp16_10 (
    .a(i16[10]),
    .b(sum_15[10]),
    .c(cout_16[9]),
    .cout(cout_16[10]),
    .sum(sum_16[10]));
  AL_FADD comp16_11 (
    .a(i16[11]),
    .b(sum_15[11]),
    .c(cout_16[10]),
    .cout(cout_16[11]),
    .sum(sum_16[11]));
  AL_FADD comp16_12 (
    .a(i16[12]),
    .b(sum_15[12]),
    .c(cout_16[11]),
    .cout(cout_16[12]),
    .sum(sum_16[12]));
  AL_FADD comp16_13 (
    .a(i16[13]),
    .b(sum_15[13]),
    .c(cout_16[12]),
    .cout(cout_16[13]),
    .sum(sum_16[13]));
  AL_FADD comp16_14 (
    .a(i16[14]),
    .b(sum_15[14]),
    .c(cout_16[13]),
    .cout(cout_16[14]),
    .sum(sum_16[14]));
  AL_FADD comp16_15 (
    .a(i16[15]),
    .b(sum_15[15]),
    .c(cout_16[14]),
    .cout(cout_16[15]),
    .sum(sum_16[15]));
  AL_FADD comp16_16 (
    .a(i16[16]),
    .b(sum_15[16]),
    .c(cout_16[15]),
    .cout(cout_16[16]),
    .sum(sum_16[16]));
  AL_FADD comp16_17 (
    .a(i16[17]),
    .b(sum_15[17]),
    .c(cout_16[16]),
    .cout(cout_16[17]),
    .sum(sum_16[17]));
  AL_FADD comp16_18 (
    .a(i16[18]),
    .b(sum_15[18]),
    .c(cout_16[17]),
    .cout(cout_16[18]),
    .sum(sum_16[18]));
  AL_FADD comp16_19 (
    .a(i16[19]),
    .b(sum_15[19]),
    .c(cout_16[18]),
    .cout(cout_16[19]),
    .sum(sum_16[19]));
  AL_FADD comp16_2 (
    .a(i16[2]),
    .b(sum_15[2]),
    .c(cout_16[1]),
    .cout(cout_16[2]),
    .sum(sum_16[2]));
  AL_FADD comp16_20 (
    .a(i16[20]),
    .b(sum_15[20]),
    .c(cout_16[19]),
    .cout(cout_16[20]),
    .sum(sum_16[20]));
  AL_FADD comp16_21 (
    .a(i16[21]),
    .b(sum_15[21]),
    .c(cout_16[20]),
    .cout(cout_16[21]),
    .sum(sum_16[21]));
  AL_FADD comp16_22 (
    .a(i16[22]),
    .b(sum_15[22]),
    .c(cout_16[21]),
    .cout(cout_16[22]),
    .sum(sum_16[22]));
  AL_FADD comp16_23 (
    .a(i16[23]),
    .b(sum_15[23]),
    .c(cout_16[22]),
    .cout(cout_16[23]),
    .sum(sum_16[23]));
  AL_FADD comp16_24 (
    .a(i16[24]),
    .b(sum_15[24]),
    .c(cout_16[23]),
    .cout(cout_16[24]),
    .sum(sum_16[24]));
  AL_FADD comp16_25 (
    .a(i16[25]),
    .b(sum_15[25]),
    .c(cout_16[24]),
    .cout(cout_16[25]),
    .sum(sum_16[25]));
  AL_FADD comp16_26 (
    .a(i16[26]),
    .b(sum_15[26]),
    .c(cout_16[25]),
    .cout(cout_16[26]),
    .sum(sum_16[26]));
  AL_FADD comp16_27 (
    .a(i16[27]),
    .b(sum_15[27]),
    .c(cout_16[26]),
    .cout(cout_16[27]),
    .sum(sum_16[27]));
  AL_FADD comp16_28 (
    .a(i16[28]),
    .b(sum_15[28]),
    .c(cout_16[27]),
    .cout(cout_16[28]),
    .sum(sum_16[28]));
  AL_FADD comp16_29 (
    .a(i16[29]),
    .b(sum_15[29]),
    .c(cout_16[28]),
    .cout(cout_16[29]),
    .sum(sum_16[29]));
  AL_FADD comp16_3 (
    .a(i16[3]),
    .b(sum_15[3]),
    .c(cout_16[2]),
    .cout(cout_16[3]),
    .sum(sum_16[3]));
  AL_FADD comp16_30 (
    .a(i16[30]),
    .b(sum_15[30]),
    .c(cout_16[29]),
    .cout(cout_16[30]),
    .sum(sum_16[30]));
  AL_FADD comp16_31 (
    .a(i16[31]),
    .b(sum_15[31]),
    .c(cout_16[30]),
    .cout(cout_16[31]),
    .sum(sum_16[31]));
  AL_FADD comp16_32 (
    .a(i16[32]),
    .b(sum_15[32]),
    .c(cout_16[31]),
    .cout(cout_16[32]),
    .sum(sum_16[32]));
  AL_FADD comp16_33 (
    .a(i16[33]),
    .b(sum_15[33]),
    .c(cout_16[32]),
    .cout(cout_16[33]),
    .sum(sum_16[33]));
  AL_FADD comp16_34 (
    .a(i16[34]),
    .b(sum_15[34]),
    .c(cout_16[33]),
    .cout(cout_16[34]),
    .sum(sum_16[34]));
  AL_FADD comp16_35 (
    .a(i16[35]),
    .b(sum_15[35]),
    .c(cout_16[34]),
    .cout(cout_16[35]),
    .sum(sum_16[35]));
  AL_FADD comp16_36 (
    .a(i16[36]),
    .b(sum_15[36]),
    .c(cout_16[35]),
    .cout(cout_16[36]),
    .sum(sum_16[36]));
  AL_FADD comp16_37 (
    .a(i16[37]),
    .b(sum_15[37]),
    .c(cout_16[36]),
    .cout(cout_16[37]),
    .sum(sum_16[37]));
  AL_FADD comp16_38 (
    .a(i16[38]),
    .b(sum_15[38]),
    .c(cout_16[37]),
    .cout(cout_16[38]),
    .sum(sum_16[38]));
  AL_FADD comp16_39 (
    .a(i16[39]),
    .b(sum_15[39]),
    .c(cout_16[38]),
    .cout(cout_16[39]),
    .sum(sum_16[39]));
  AL_FADD comp16_4 (
    .a(i16[4]),
    .b(sum_15[4]),
    .c(cout_16[3]),
    .cout(cout_16[4]),
    .sum(sum_16[4]));
  AL_FADD comp16_40 (
    .a(i16[40]),
    .b(sum_15[40]),
    .c(cout_16[39]),
    .cout(cout_16[40]),
    .sum(sum_16[40]));
  AL_FADD comp16_41 (
    .a(i16[41]),
    .b(sum_15[41]),
    .c(cout_16[40]),
    .cout(cout_16[41]),
    .sum(sum_16[41]));
  AL_FADD comp16_42 (
    .a(i16[42]),
    .b(sum_15[42]),
    .c(cout_16[41]),
    .cout(cout_16[42]),
    .sum(sum_16[42]));
  AL_FADD comp16_43 (
    .a(i16[43]),
    .b(sum_15[43]),
    .c(cout_16[42]),
    .cout(cout_16[43]),
    .sum(sum_16[43]));
  AL_FADD comp16_44 (
    .a(i16[44]),
    .b(sum_15[44]),
    .c(cout_16[43]),
    .cout(cout_16[44]),
    .sum(sum_16[44]));
  AL_FADD comp16_45 (
    .a(1'b0),
    .b(sum_15[45]),
    .c(cout_16[44]),
    .cout(cout_16[45]),
    .sum(sum_16[45]));
  AL_FADD comp16_46 (
    .a(1'b0),
    .b(sum_15[46]),
    .c(cout_16[45]),
    .cout(cout_16[46]),
    .sum(sum_16[46]));
  AL_FADD comp16_47 (
    .a(1'b0),
    .b(sum_15[47]),
    .c(cout_16[46]),
    .cout(cout_16[47]),
    .sum(sum_16[47]));
  AL_FADD comp16_48 (
    .a(1'b0),
    .b(sum_15[48]),
    .c(cout_16[47]),
    .cout(cout_16[48]),
    .sum(sum_16[48]));
  AL_FADD comp16_49 (
    .a(1'b0),
    .b(sum_15[49]),
    .c(cout_16[48]),
    .cout(cout_16[49]),
    .sum(sum_16[49]));
  AL_FADD comp16_5 (
    .a(i16[5]),
    .b(sum_15[5]),
    .c(cout_16[4]),
    .cout(cout_16[5]),
    .sum(sum_16[5]));
  AL_FADD comp16_50 (
    .a(1'b0),
    .b(sum_15[50]),
    .c(cout_16[49]),
    .cout(cout_16[50]),
    .sum(sum_16[50]));
  AL_FADD comp16_51 (
    .a(1'b0),
    .b(sum_15[51]),
    .c(cout_16[50]),
    .cout(cout_16[51]),
    .sum(sum_16[51]));
  AL_FADD comp16_52 (
    .a(1'b0),
    .b(sum_15[52]),
    .c(cout_16[51]),
    .cout(cout_16[52]),
    .sum(sum_16[52]));
  AL_FADD comp16_53 (
    .a(1'b0),
    .b(sum_15[53]),
    .c(cout_16[52]),
    .cout(cout_16[53]),
    .sum(sum_16[53]));
  AL_FADD comp16_54 (
    .a(1'b0),
    .b(sum_15[54]),
    .c(cout_16[53]),
    .cout(cout_16[54]),
    .sum(sum_16[54]));
  AL_FADD comp16_55 (
    .a(1'b0),
    .b(sum_15[55]),
    .c(cout_16[54]),
    .cout(cout_16[55]),
    .sum(sum_16[55]));
  AL_FADD comp16_56 (
    .a(1'b0),
    .b(sum_15[56]),
    .c(cout_16[55]),
    .cout(cout_16[56]),
    .sum(sum_16[56]));
  AL_FADD comp16_57 (
    .a(1'b0),
    .b(sum_15[57]),
    .c(cout_16[56]),
    .cout(cout_16[57]),
    .sum(sum_16[57]));
  AL_FADD comp16_58 (
    .a(1'b0),
    .b(sum_15[58]),
    .c(cout_16[57]),
    .cout(cout_16[58]),
    .sum(sum_16[58]));
  AL_FADD comp16_59 (
    .a(1'b0),
    .b(sum_15[59]),
    .c(cout_16[58]),
    .cout(cout_16[59]),
    .sum(sum_16[59]));
  AL_FADD comp16_6 (
    .a(i16[6]),
    .b(sum_15[6]),
    .c(cout_16[5]),
    .cout(cout_16[6]),
    .sum(sum_16[6]));
  AL_FADD comp16_60 (
    .a(1'b0),
    .b(sum_15[60]),
    .c(cout_16[59]),
    .cout(cout_16[60]),
    .sum(sum_16[60]));
  AL_FADD comp16_61 (
    .a(1'b0),
    .b(sum_15[61]),
    .c(cout_16[60]),
    .cout(cout_16[61]),
    .sum(sum_16[61]));
  AL_FADD comp16_62 (
    .a(1'b0),
    .b(sum_15[62]),
    .c(cout_16[61]),
    .cout(cout_16[62]),
    .sum(sum_16[62]));
  AL_FADD comp16_63 (
    .a(1'b0),
    .b(sum_15[63]),
    .c(cout_16[62]),
    .cout(cout_16[63]),
    .sum(sum_16[63]));
  AL_FADD comp16_7 (
    .a(i16[7]),
    .b(sum_15[7]),
    .c(cout_16[6]),
    .cout(cout_16[7]),
    .sum(sum_16[7]));
  AL_FADD comp16_8 (
    .a(i16[8]),
    .b(sum_15[8]),
    .c(cout_16[7]),
    .cout(cout_16[8]),
    .sum(sum_16[8]));
  AL_FADD comp16_9 (
    .a(i16[9]),
    .b(sum_15[9]),
    .c(cout_16[8]),
    .cout(cout_16[9]),
    .sum(sum_16[9]));
  AL_FADD comp17_0 (
    .a(i17[0]),
    .b(sum_16[0]),
    .c(1'b0),
    .cout(cout_17[0]),
    .sum(sum_17[0]));
  AL_FADD comp17_1 (
    .a(i17[1]),
    .b(sum_16[1]),
    .c(cout_17[0]),
    .cout(cout_17[1]),
    .sum(sum_17[1]));
  AL_FADD comp17_10 (
    .a(i17[10]),
    .b(sum_16[10]),
    .c(cout_17[9]),
    .cout(cout_17[10]),
    .sum(sum_17[10]));
  AL_FADD comp17_11 (
    .a(i17[11]),
    .b(sum_16[11]),
    .c(cout_17[10]),
    .cout(cout_17[11]),
    .sum(sum_17[11]));
  AL_FADD comp17_12 (
    .a(i17[12]),
    .b(sum_16[12]),
    .c(cout_17[11]),
    .cout(cout_17[12]),
    .sum(sum_17[12]));
  AL_FADD comp17_13 (
    .a(i17[13]),
    .b(sum_16[13]),
    .c(cout_17[12]),
    .cout(cout_17[13]),
    .sum(sum_17[13]));
  AL_FADD comp17_14 (
    .a(i17[14]),
    .b(sum_16[14]),
    .c(cout_17[13]),
    .cout(cout_17[14]),
    .sum(sum_17[14]));
  AL_FADD comp17_15 (
    .a(i17[15]),
    .b(sum_16[15]),
    .c(cout_17[14]),
    .cout(cout_17[15]),
    .sum(sum_17[15]));
  AL_FADD comp17_16 (
    .a(i17[16]),
    .b(sum_16[16]),
    .c(cout_17[15]),
    .cout(cout_17[16]),
    .sum(sum_17[16]));
  AL_FADD comp17_17 (
    .a(i17[17]),
    .b(sum_16[17]),
    .c(cout_17[16]),
    .cout(cout_17[17]),
    .sum(sum_17[17]));
  AL_FADD comp17_18 (
    .a(i17[18]),
    .b(sum_16[18]),
    .c(cout_17[17]),
    .cout(cout_17[18]),
    .sum(sum_17[18]));
  AL_FADD comp17_19 (
    .a(i17[19]),
    .b(sum_16[19]),
    .c(cout_17[18]),
    .cout(cout_17[19]),
    .sum(sum_17[19]));
  AL_FADD comp17_2 (
    .a(i17[2]),
    .b(sum_16[2]),
    .c(cout_17[1]),
    .cout(cout_17[2]),
    .sum(sum_17[2]));
  AL_FADD comp17_20 (
    .a(i17[20]),
    .b(sum_16[20]),
    .c(cout_17[19]),
    .cout(cout_17[20]),
    .sum(sum_17[20]));
  AL_FADD comp17_21 (
    .a(i17[21]),
    .b(sum_16[21]),
    .c(cout_17[20]),
    .cout(cout_17[21]),
    .sum(sum_17[21]));
  AL_FADD comp17_22 (
    .a(i17[22]),
    .b(sum_16[22]),
    .c(cout_17[21]),
    .cout(cout_17[22]),
    .sum(sum_17[22]));
  AL_FADD comp17_23 (
    .a(i17[23]),
    .b(sum_16[23]),
    .c(cout_17[22]),
    .cout(cout_17[23]),
    .sum(sum_17[23]));
  AL_FADD comp17_24 (
    .a(i17[24]),
    .b(sum_16[24]),
    .c(cout_17[23]),
    .cout(cout_17[24]),
    .sum(sum_17[24]));
  AL_FADD comp17_25 (
    .a(i17[25]),
    .b(sum_16[25]),
    .c(cout_17[24]),
    .cout(cout_17[25]),
    .sum(sum_17[25]));
  AL_FADD comp17_26 (
    .a(i17[26]),
    .b(sum_16[26]),
    .c(cout_17[25]),
    .cout(cout_17[26]),
    .sum(sum_17[26]));
  AL_FADD comp17_27 (
    .a(i17[27]),
    .b(sum_16[27]),
    .c(cout_17[26]),
    .cout(cout_17[27]),
    .sum(sum_17[27]));
  AL_FADD comp17_28 (
    .a(i17[28]),
    .b(sum_16[28]),
    .c(cout_17[27]),
    .cout(cout_17[28]),
    .sum(sum_17[28]));
  AL_FADD comp17_29 (
    .a(i17[29]),
    .b(sum_16[29]),
    .c(cout_17[28]),
    .cout(cout_17[29]),
    .sum(sum_17[29]));
  AL_FADD comp17_3 (
    .a(i17[3]),
    .b(sum_16[3]),
    .c(cout_17[2]),
    .cout(cout_17[3]),
    .sum(sum_17[3]));
  AL_FADD comp17_30 (
    .a(i17[30]),
    .b(sum_16[30]),
    .c(cout_17[29]),
    .cout(cout_17[30]),
    .sum(sum_17[30]));
  AL_FADD comp17_31 (
    .a(i17[31]),
    .b(sum_16[31]),
    .c(cout_17[30]),
    .cout(cout_17[31]),
    .sum(sum_17[31]));
  AL_FADD comp17_32 (
    .a(i17[32]),
    .b(sum_16[32]),
    .c(cout_17[31]),
    .cout(cout_17[32]),
    .sum(sum_17[32]));
  AL_FADD comp17_33 (
    .a(i17[33]),
    .b(sum_16[33]),
    .c(cout_17[32]),
    .cout(cout_17[33]),
    .sum(sum_17[33]));
  AL_FADD comp17_34 (
    .a(i17[34]),
    .b(sum_16[34]),
    .c(cout_17[33]),
    .cout(cout_17[34]),
    .sum(sum_17[34]));
  AL_FADD comp17_35 (
    .a(i17[35]),
    .b(sum_16[35]),
    .c(cout_17[34]),
    .cout(cout_17[35]),
    .sum(sum_17[35]));
  AL_FADD comp17_36 (
    .a(i17[36]),
    .b(sum_16[36]),
    .c(cout_17[35]),
    .cout(cout_17[36]),
    .sum(sum_17[36]));
  AL_FADD comp17_37 (
    .a(i17[37]),
    .b(sum_16[37]),
    .c(cout_17[36]),
    .cout(cout_17[37]),
    .sum(sum_17[37]));
  AL_FADD comp17_38 (
    .a(i17[38]),
    .b(sum_16[38]),
    .c(cout_17[37]),
    .cout(cout_17[38]),
    .sum(sum_17[38]));
  AL_FADD comp17_39 (
    .a(i17[39]),
    .b(sum_16[39]),
    .c(cout_17[38]),
    .cout(cout_17[39]),
    .sum(sum_17[39]));
  AL_FADD comp17_4 (
    .a(i17[4]),
    .b(sum_16[4]),
    .c(cout_17[3]),
    .cout(cout_17[4]),
    .sum(sum_17[4]));
  AL_FADD comp17_40 (
    .a(i17[40]),
    .b(sum_16[40]),
    .c(cout_17[39]),
    .cout(cout_17[40]),
    .sum(sum_17[40]));
  AL_FADD comp17_41 (
    .a(i17[41]),
    .b(sum_16[41]),
    .c(cout_17[40]),
    .cout(cout_17[41]),
    .sum(sum_17[41]));
  AL_FADD comp17_42 (
    .a(i17[42]),
    .b(sum_16[42]),
    .c(cout_17[41]),
    .cout(cout_17[42]),
    .sum(sum_17[42]));
  AL_FADD comp17_43 (
    .a(i17[43]),
    .b(sum_16[43]),
    .c(cout_17[42]),
    .cout(cout_17[43]),
    .sum(sum_17[43]));
  AL_FADD comp17_44 (
    .a(1'b0),
    .b(sum_16[44]),
    .c(cout_17[43]),
    .cout(cout_17[44]),
    .sum(sum_17[44]));
  AL_FADD comp17_45 (
    .a(1'b0),
    .b(sum_16[45]),
    .c(cout_17[44]),
    .cout(cout_17[45]),
    .sum(sum_17[45]));
  AL_FADD comp17_46 (
    .a(1'b0),
    .b(sum_16[46]),
    .c(cout_17[45]),
    .cout(cout_17[46]),
    .sum(sum_17[46]));
  AL_FADD comp17_47 (
    .a(1'b0),
    .b(sum_16[47]),
    .c(cout_17[46]),
    .cout(cout_17[47]),
    .sum(sum_17[47]));
  AL_FADD comp17_48 (
    .a(1'b0),
    .b(sum_16[48]),
    .c(cout_17[47]),
    .cout(cout_17[48]),
    .sum(sum_17[48]));
  AL_FADD comp17_49 (
    .a(1'b0),
    .b(sum_16[49]),
    .c(cout_17[48]),
    .cout(cout_17[49]),
    .sum(sum_17[49]));
  AL_FADD comp17_5 (
    .a(i17[5]),
    .b(sum_16[5]),
    .c(cout_17[4]),
    .cout(cout_17[5]),
    .sum(sum_17[5]));
  AL_FADD comp17_50 (
    .a(1'b0),
    .b(sum_16[50]),
    .c(cout_17[49]),
    .cout(cout_17[50]),
    .sum(sum_17[50]));
  AL_FADD comp17_51 (
    .a(1'b0),
    .b(sum_16[51]),
    .c(cout_17[50]),
    .cout(cout_17[51]),
    .sum(sum_17[51]));
  AL_FADD comp17_52 (
    .a(1'b0),
    .b(sum_16[52]),
    .c(cout_17[51]),
    .cout(cout_17[52]),
    .sum(sum_17[52]));
  AL_FADD comp17_53 (
    .a(1'b0),
    .b(sum_16[53]),
    .c(cout_17[52]),
    .cout(cout_17[53]),
    .sum(sum_17[53]));
  AL_FADD comp17_54 (
    .a(1'b0),
    .b(sum_16[54]),
    .c(cout_17[53]),
    .cout(cout_17[54]),
    .sum(sum_17[54]));
  AL_FADD comp17_55 (
    .a(1'b0),
    .b(sum_16[55]),
    .c(cout_17[54]),
    .cout(cout_17[55]),
    .sum(sum_17[55]));
  AL_FADD comp17_56 (
    .a(1'b0),
    .b(sum_16[56]),
    .c(cout_17[55]),
    .cout(cout_17[56]),
    .sum(sum_17[56]));
  AL_FADD comp17_57 (
    .a(1'b0),
    .b(sum_16[57]),
    .c(cout_17[56]),
    .cout(cout_17[57]),
    .sum(sum_17[57]));
  AL_FADD comp17_58 (
    .a(1'b0),
    .b(sum_16[58]),
    .c(cout_17[57]),
    .cout(cout_17[58]),
    .sum(sum_17[58]));
  AL_FADD comp17_59 (
    .a(1'b0),
    .b(sum_16[59]),
    .c(cout_17[58]),
    .cout(cout_17[59]),
    .sum(sum_17[59]));
  AL_FADD comp17_6 (
    .a(i17[6]),
    .b(sum_16[6]),
    .c(cout_17[5]),
    .cout(cout_17[6]),
    .sum(sum_17[6]));
  AL_FADD comp17_60 (
    .a(1'b0),
    .b(sum_16[60]),
    .c(cout_17[59]),
    .cout(cout_17[60]),
    .sum(sum_17[60]));
  AL_FADD comp17_61 (
    .a(1'b0),
    .b(sum_16[61]),
    .c(cout_17[60]),
    .cout(cout_17[61]),
    .sum(sum_17[61]));
  AL_FADD comp17_62 (
    .a(1'b0),
    .b(sum_16[62]),
    .c(cout_17[61]),
    .cout(cout_17[62]),
    .sum(sum_17[62]));
  AL_FADD comp17_63 (
    .a(1'b0),
    .b(sum_16[63]),
    .c(cout_17[62]),
    .cout(cout_17[63]),
    .sum(sum_17[63]));
  AL_FADD comp17_7 (
    .a(i17[7]),
    .b(sum_16[7]),
    .c(cout_17[6]),
    .cout(cout_17[7]),
    .sum(sum_17[7]));
  AL_FADD comp17_8 (
    .a(i17[8]),
    .b(sum_16[8]),
    .c(cout_17[7]),
    .cout(cout_17[8]),
    .sum(sum_17[8]));
  AL_FADD comp17_9 (
    .a(i17[9]),
    .b(sum_16[9]),
    .c(cout_17[8]),
    .cout(cout_17[9]),
    .sum(sum_17[9]));
  AL_FADD comp18_0 (
    .a(i18[0]),
    .b(sum_17[0]),
    .c(1'b0),
    .cout(cout_18[0]),
    .sum(sum_18[0]));
  AL_FADD comp18_1 (
    .a(i18[1]),
    .b(sum_17[1]),
    .c(cout_18[0]),
    .cout(cout_18[1]),
    .sum(sum_18[1]));
  AL_FADD comp18_10 (
    .a(i18[10]),
    .b(sum_17[10]),
    .c(cout_18[9]),
    .cout(cout_18[10]),
    .sum(sum_18[10]));
  AL_FADD comp18_11 (
    .a(i18[11]),
    .b(sum_17[11]),
    .c(cout_18[10]),
    .cout(cout_18[11]),
    .sum(sum_18[11]));
  AL_FADD comp18_12 (
    .a(i18[12]),
    .b(sum_17[12]),
    .c(cout_18[11]),
    .cout(cout_18[12]),
    .sum(sum_18[12]));
  AL_FADD comp18_13 (
    .a(i18[13]),
    .b(sum_17[13]),
    .c(cout_18[12]),
    .cout(cout_18[13]),
    .sum(sum_18[13]));
  AL_FADD comp18_14 (
    .a(i18[14]),
    .b(sum_17[14]),
    .c(cout_18[13]),
    .cout(cout_18[14]),
    .sum(sum_18[14]));
  AL_FADD comp18_15 (
    .a(i18[15]),
    .b(sum_17[15]),
    .c(cout_18[14]),
    .cout(cout_18[15]),
    .sum(sum_18[15]));
  AL_FADD comp18_16 (
    .a(i18[16]),
    .b(sum_17[16]),
    .c(cout_18[15]),
    .cout(cout_18[16]),
    .sum(sum_18[16]));
  AL_FADD comp18_17 (
    .a(i18[17]),
    .b(sum_17[17]),
    .c(cout_18[16]),
    .cout(cout_18[17]),
    .sum(sum_18[17]));
  AL_FADD comp18_18 (
    .a(i18[18]),
    .b(sum_17[18]),
    .c(cout_18[17]),
    .cout(cout_18[18]),
    .sum(sum_18[18]));
  AL_FADD comp18_19 (
    .a(i18[19]),
    .b(sum_17[19]),
    .c(cout_18[18]),
    .cout(cout_18[19]),
    .sum(sum_18[19]));
  AL_FADD comp18_2 (
    .a(i18[2]),
    .b(sum_17[2]),
    .c(cout_18[1]),
    .cout(cout_18[2]),
    .sum(sum_18[2]));
  AL_FADD comp18_20 (
    .a(i18[20]),
    .b(sum_17[20]),
    .c(cout_18[19]),
    .cout(cout_18[20]),
    .sum(sum_18[20]));
  AL_FADD comp18_21 (
    .a(i18[21]),
    .b(sum_17[21]),
    .c(cout_18[20]),
    .cout(cout_18[21]),
    .sum(sum_18[21]));
  AL_FADD comp18_22 (
    .a(i18[22]),
    .b(sum_17[22]),
    .c(cout_18[21]),
    .cout(cout_18[22]),
    .sum(sum_18[22]));
  AL_FADD comp18_23 (
    .a(i18[23]),
    .b(sum_17[23]),
    .c(cout_18[22]),
    .cout(cout_18[23]),
    .sum(sum_18[23]));
  AL_FADD comp18_24 (
    .a(i18[24]),
    .b(sum_17[24]),
    .c(cout_18[23]),
    .cout(cout_18[24]),
    .sum(sum_18[24]));
  AL_FADD comp18_25 (
    .a(i18[25]),
    .b(sum_17[25]),
    .c(cout_18[24]),
    .cout(cout_18[25]),
    .sum(sum_18[25]));
  AL_FADD comp18_26 (
    .a(i18[26]),
    .b(sum_17[26]),
    .c(cout_18[25]),
    .cout(cout_18[26]),
    .sum(sum_18[26]));
  AL_FADD comp18_27 (
    .a(i18[27]),
    .b(sum_17[27]),
    .c(cout_18[26]),
    .cout(cout_18[27]),
    .sum(sum_18[27]));
  AL_FADD comp18_28 (
    .a(i18[28]),
    .b(sum_17[28]),
    .c(cout_18[27]),
    .cout(cout_18[28]),
    .sum(sum_18[28]));
  AL_FADD comp18_29 (
    .a(i18[29]),
    .b(sum_17[29]),
    .c(cout_18[28]),
    .cout(cout_18[29]),
    .sum(sum_18[29]));
  AL_FADD comp18_3 (
    .a(i18[3]),
    .b(sum_17[3]),
    .c(cout_18[2]),
    .cout(cout_18[3]),
    .sum(sum_18[3]));
  AL_FADD comp18_30 (
    .a(i18[30]),
    .b(sum_17[30]),
    .c(cout_18[29]),
    .cout(cout_18[30]),
    .sum(sum_18[30]));
  AL_FADD comp18_31 (
    .a(i18[31]),
    .b(sum_17[31]),
    .c(cout_18[30]),
    .cout(cout_18[31]),
    .sum(sum_18[31]));
  AL_FADD comp18_32 (
    .a(i18[32]),
    .b(sum_17[32]),
    .c(cout_18[31]),
    .cout(cout_18[32]),
    .sum(sum_18[32]));
  AL_FADD comp18_33 (
    .a(i18[33]),
    .b(sum_17[33]),
    .c(cout_18[32]),
    .cout(cout_18[33]),
    .sum(sum_18[33]));
  AL_FADD comp18_34 (
    .a(i18[34]),
    .b(sum_17[34]),
    .c(cout_18[33]),
    .cout(cout_18[34]),
    .sum(sum_18[34]));
  AL_FADD comp18_35 (
    .a(i18[35]),
    .b(sum_17[35]),
    .c(cout_18[34]),
    .cout(cout_18[35]),
    .sum(sum_18[35]));
  AL_FADD comp18_36 (
    .a(i18[36]),
    .b(sum_17[36]),
    .c(cout_18[35]),
    .cout(cout_18[36]),
    .sum(sum_18[36]));
  AL_FADD comp18_37 (
    .a(i18[37]),
    .b(sum_17[37]),
    .c(cout_18[36]),
    .cout(cout_18[37]),
    .sum(sum_18[37]));
  AL_FADD comp18_38 (
    .a(i18[38]),
    .b(sum_17[38]),
    .c(cout_18[37]),
    .cout(cout_18[38]),
    .sum(sum_18[38]));
  AL_FADD comp18_39 (
    .a(i18[39]),
    .b(sum_17[39]),
    .c(cout_18[38]),
    .cout(cout_18[39]),
    .sum(sum_18[39]));
  AL_FADD comp18_4 (
    .a(i18[4]),
    .b(sum_17[4]),
    .c(cout_18[3]),
    .cout(cout_18[4]),
    .sum(sum_18[4]));
  AL_FADD comp18_40 (
    .a(i18[40]),
    .b(sum_17[40]),
    .c(cout_18[39]),
    .cout(cout_18[40]),
    .sum(sum_18[40]));
  AL_FADD comp18_41 (
    .a(i18[41]),
    .b(sum_17[41]),
    .c(cout_18[40]),
    .cout(cout_18[41]),
    .sum(sum_18[41]));
  AL_FADD comp18_42 (
    .a(i18[42]),
    .b(sum_17[42]),
    .c(cout_18[41]),
    .cout(cout_18[42]),
    .sum(sum_18[42]));
  AL_FADD comp18_43 (
    .a(1'b0),
    .b(sum_17[43]),
    .c(cout_18[42]),
    .cout(cout_18[43]),
    .sum(sum_18[43]));
  AL_FADD comp18_44 (
    .a(1'b0),
    .b(sum_17[44]),
    .c(cout_18[43]),
    .cout(cout_18[44]),
    .sum(sum_18[44]));
  AL_FADD comp18_45 (
    .a(1'b0),
    .b(sum_17[45]),
    .c(cout_18[44]),
    .cout(cout_18[45]),
    .sum(sum_18[45]));
  AL_FADD comp18_46 (
    .a(1'b0),
    .b(sum_17[46]),
    .c(cout_18[45]),
    .cout(cout_18[46]),
    .sum(sum_18[46]));
  AL_FADD comp18_47 (
    .a(1'b0),
    .b(sum_17[47]),
    .c(cout_18[46]),
    .cout(cout_18[47]),
    .sum(sum_18[47]));
  AL_FADD comp18_48 (
    .a(1'b0),
    .b(sum_17[48]),
    .c(cout_18[47]),
    .cout(cout_18[48]),
    .sum(sum_18[48]));
  AL_FADD comp18_49 (
    .a(1'b0),
    .b(sum_17[49]),
    .c(cout_18[48]),
    .cout(cout_18[49]),
    .sum(sum_18[49]));
  AL_FADD comp18_5 (
    .a(i18[5]),
    .b(sum_17[5]),
    .c(cout_18[4]),
    .cout(cout_18[5]),
    .sum(sum_18[5]));
  AL_FADD comp18_50 (
    .a(1'b0),
    .b(sum_17[50]),
    .c(cout_18[49]),
    .cout(cout_18[50]),
    .sum(sum_18[50]));
  AL_FADD comp18_51 (
    .a(1'b0),
    .b(sum_17[51]),
    .c(cout_18[50]),
    .cout(cout_18[51]),
    .sum(sum_18[51]));
  AL_FADD comp18_52 (
    .a(1'b0),
    .b(sum_17[52]),
    .c(cout_18[51]),
    .cout(cout_18[52]),
    .sum(sum_18[52]));
  AL_FADD comp18_53 (
    .a(1'b0),
    .b(sum_17[53]),
    .c(cout_18[52]),
    .cout(cout_18[53]),
    .sum(sum_18[53]));
  AL_FADD comp18_54 (
    .a(1'b0),
    .b(sum_17[54]),
    .c(cout_18[53]),
    .cout(cout_18[54]),
    .sum(sum_18[54]));
  AL_FADD comp18_55 (
    .a(1'b0),
    .b(sum_17[55]),
    .c(cout_18[54]),
    .cout(cout_18[55]),
    .sum(sum_18[55]));
  AL_FADD comp18_56 (
    .a(1'b0),
    .b(sum_17[56]),
    .c(cout_18[55]),
    .cout(cout_18[56]),
    .sum(sum_18[56]));
  AL_FADD comp18_57 (
    .a(1'b0),
    .b(sum_17[57]),
    .c(cout_18[56]),
    .cout(cout_18[57]),
    .sum(sum_18[57]));
  AL_FADD comp18_58 (
    .a(1'b0),
    .b(sum_17[58]),
    .c(cout_18[57]),
    .cout(cout_18[58]),
    .sum(sum_18[58]));
  AL_FADD comp18_59 (
    .a(1'b0),
    .b(sum_17[59]),
    .c(cout_18[58]),
    .cout(cout_18[59]),
    .sum(sum_18[59]));
  AL_FADD comp18_6 (
    .a(i18[6]),
    .b(sum_17[6]),
    .c(cout_18[5]),
    .cout(cout_18[6]),
    .sum(sum_18[6]));
  AL_FADD comp18_60 (
    .a(1'b0),
    .b(sum_17[60]),
    .c(cout_18[59]),
    .cout(cout_18[60]),
    .sum(sum_18[60]));
  AL_FADD comp18_61 (
    .a(1'b0),
    .b(sum_17[61]),
    .c(cout_18[60]),
    .cout(cout_18[61]),
    .sum(sum_18[61]));
  AL_FADD comp18_62 (
    .a(1'b0),
    .b(sum_17[62]),
    .c(cout_18[61]),
    .cout(cout_18[62]),
    .sum(sum_18[62]));
  AL_FADD comp18_63 (
    .a(1'b0),
    .b(sum_17[63]),
    .c(cout_18[62]),
    .cout(cout_18[63]),
    .sum(sum_18[63]));
  AL_FADD comp18_7 (
    .a(i18[7]),
    .b(sum_17[7]),
    .c(cout_18[6]),
    .cout(cout_18[7]),
    .sum(sum_18[7]));
  AL_FADD comp18_8 (
    .a(i18[8]),
    .b(sum_17[8]),
    .c(cout_18[7]),
    .cout(cout_18[8]),
    .sum(sum_18[8]));
  AL_FADD comp18_9 (
    .a(i18[9]),
    .b(sum_17[9]),
    .c(cout_18[8]),
    .cout(cout_18[9]),
    .sum(sum_18[9]));
  AL_FADD comp19_0 (
    .a(i19[0]),
    .b(sum_18[0]),
    .c(1'b0),
    .cout(cout_19[0]),
    .sum(sum_19[0]));
  AL_FADD comp19_1 (
    .a(i19[1]),
    .b(sum_18[1]),
    .c(cout_19[0]),
    .cout(cout_19[1]),
    .sum(sum_19[1]));
  AL_FADD comp19_10 (
    .a(i19[10]),
    .b(sum_18[10]),
    .c(cout_19[9]),
    .cout(cout_19[10]),
    .sum(sum_19[10]));
  AL_FADD comp19_11 (
    .a(i19[11]),
    .b(sum_18[11]),
    .c(cout_19[10]),
    .cout(cout_19[11]),
    .sum(sum_19[11]));
  AL_FADD comp19_12 (
    .a(i19[12]),
    .b(sum_18[12]),
    .c(cout_19[11]),
    .cout(cout_19[12]),
    .sum(sum_19[12]));
  AL_FADD comp19_13 (
    .a(i19[13]),
    .b(sum_18[13]),
    .c(cout_19[12]),
    .cout(cout_19[13]),
    .sum(sum_19[13]));
  AL_FADD comp19_14 (
    .a(i19[14]),
    .b(sum_18[14]),
    .c(cout_19[13]),
    .cout(cout_19[14]),
    .sum(sum_19[14]));
  AL_FADD comp19_15 (
    .a(i19[15]),
    .b(sum_18[15]),
    .c(cout_19[14]),
    .cout(cout_19[15]),
    .sum(sum_19[15]));
  AL_FADD comp19_16 (
    .a(i19[16]),
    .b(sum_18[16]),
    .c(cout_19[15]),
    .cout(cout_19[16]),
    .sum(sum_19[16]));
  AL_FADD comp19_17 (
    .a(i19[17]),
    .b(sum_18[17]),
    .c(cout_19[16]),
    .cout(cout_19[17]),
    .sum(sum_19[17]));
  AL_FADD comp19_18 (
    .a(i19[18]),
    .b(sum_18[18]),
    .c(cout_19[17]),
    .cout(cout_19[18]),
    .sum(sum_19[18]));
  AL_FADD comp19_19 (
    .a(i19[19]),
    .b(sum_18[19]),
    .c(cout_19[18]),
    .cout(cout_19[19]),
    .sum(sum_19[19]));
  AL_FADD comp19_2 (
    .a(i19[2]),
    .b(sum_18[2]),
    .c(cout_19[1]),
    .cout(cout_19[2]),
    .sum(sum_19[2]));
  AL_FADD comp19_20 (
    .a(i19[20]),
    .b(sum_18[20]),
    .c(cout_19[19]),
    .cout(cout_19[20]),
    .sum(sum_19[20]));
  AL_FADD comp19_21 (
    .a(i19[21]),
    .b(sum_18[21]),
    .c(cout_19[20]),
    .cout(cout_19[21]),
    .sum(sum_19[21]));
  AL_FADD comp19_22 (
    .a(i19[22]),
    .b(sum_18[22]),
    .c(cout_19[21]),
    .cout(cout_19[22]),
    .sum(sum_19[22]));
  AL_FADD comp19_23 (
    .a(i19[23]),
    .b(sum_18[23]),
    .c(cout_19[22]),
    .cout(cout_19[23]),
    .sum(sum_19[23]));
  AL_FADD comp19_24 (
    .a(i19[24]),
    .b(sum_18[24]),
    .c(cout_19[23]),
    .cout(cout_19[24]),
    .sum(sum_19[24]));
  AL_FADD comp19_25 (
    .a(i19[25]),
    .b(sum_18[25]),
    .c(cout_19[24]),
    .cout(cout_19[25]),
    .sum(sum_19[25]));
  AL_FADD comp19_26 (
    .a(i19[26]),
    .b(sum_18[26]),
    .c(cout_19[25]),
    .cout(cout_19[26]),
    .sum(sum_19[26]));
  AL_FADD comp19_27 (
    .a(i19[27]),
    .b(sum_18[27]),
    .c(cout_19[26]),
    .cout(cout_19[27]),
    .sum(sum_19[27]));
  AL_FADD comp19_28 (
    .a(i19[28]),
    .b(sum_18[28]),
    .c(cout_19[27]),
    .cout(cout_19[28]),
    .sum(sum_19[28]));
  AL_FADD comp19_29 (
    .a(i19[29]),
    .b(sum_18[29]),
    .c(cout_19[28]),
    .cout(cout_19[29]),
    .sum(sum_19[29]));
  AL_FADD comp19_3 (
    .a(i19[3]),
    .b(sum_18[3]),
    .c(cout_19[2]),
    .cout(cout_19[3]),
    .sum(sum_19[3]));
  AL_FADD comp19_30 (
    .a(i19[30]),
    .b(sum_18[30]),
    .c(cout_19[29]),
    .cout(cout_19[30]),
    .sum(sum_19[30]));
  AL_FADD comp19_31 (
    .a(i19[31]),
    .b(sum_18[31]),
    .c(cout_19[30]),
    .cout(cout_19[31]),
    .sum(sum_19[31]));
  AL_FADD comp19_32 (
    .a(i19[32]),
    .b(sum_18[32]),
    .c(cout_19[31]),
    .cout(cout_19[32]),
    .sum(sum_19[32]));
  AL_FADD comp19_33 (
    .a(i19[33]),
    .b(sum_18[33]),
    .c(cout_19[32]),
    .cout(cout_19[33]),
    .sum(sum_19[33]));
  AL_FADD comp19_34 (
    .a(i19[34]),
    .b(sum_18[34]),
    .c(cout_19[33]),
    .cout(cout_19[34]),
    .sum(sum_19[34]));
  AL_FADD comp19_35 (
    .a(i19[35]),
    .b(sum_18[35]),
    .c(cout_19[34]),
    .cout(cout_19[35]),
    .sum(sum_19[35]));
  AL_FADD comp19_36 (
    .a(i19[36]),
    .b(sum_18[36]),
    .c(cout_19[35]),
    .cout(cout_19[36]),
    .sum(sum_19[36]));
  AL_FADD comp19_37 (
    .a(i19[37]),
    .b(sum_18[37]),
    .c(cout_19[36]),
    .cout(cout_19[37]),
    .sum(sum_19[37]));
  AL_FADD comp19_38 (
    .a(i19[38]),
    .b(sum_18[38]),
    .c(cout_19[37]),
    .cout(cout_19[38]),
    .sum(sum_19[38]));
  AL_FADD comp19_39 (
    .a(i19[39]),
    .b(sum_18[39]),
    .c(cout_19[38]),
    .cout(cout_19[39]),
    .sum(sum_19[39]));
  AL_FADD comp19_4 (
    .a(i19[4]),
    .b(sum_18[4]),
    .c(cout_19[3]),
    .cout(cout_19[4]),
    .sum(sum_19[4]));
  AL_FADD comp19_40 (
    .a(i19[40]),
    .b(sum_18[40]),
    .c(cout_19[39]),
    .cout(cout_19[40]),
    .sum(sum_19[40]));
  AL_FADD comp19_41 (
    .a(i19[41]),
    .b(sum_18[41]),
    .c(cout_19[40]),
    .cout(cout_19[41]),
    .sum(sum_19[41]));
  AL_FADD comp19_42 (
    .a(1'b0),
    .b(sum_18[42]),
    .c(cout_19[41]),
    .cout(cout_19[42]),
    .sum(sum_19[42]));
  AL_FADD comp19_43 (
    .a(1'b0),
    .b(sum_18[43]),
    .c(cout_19[42]),
    .cout(cout_19[43]),
    .sum(sum_19[43]));
  AL_FADD comp19_44 (
    .a(1'b0),
    .b(sum_18[44]),
    .c(cout_19[43]),
    .cout(cout_19[44]),
    .sum(sum_19[44]));
  AL_FADD comp19_45 (
    .a(1'b0),
    .b(sum_18[45]),
    .c(cout_19[44]),
    .cout(cout_19[45]),
    .sum(sum_19[45]));
  AL_FADD comp19_46 (
    .a(1'b0),
    .b(sum_18[46]),
    .c(cout_19[45]),
    .cout(cout_19[46]),
    .sum(sum_19[46]));
  AL_FADD comp19_47 (
    .a(1'b0),
    .b(sum_18[47]),
    .c(cout_19[46]),
    .cout(cout_19[47]),
    .sum(sum_19[47]));
  AL_FADD comp19_48 (
    .a(1'b0),
    .b(sum_18[48]),
    .c(cout_19[47]),
    .cout(cout_19[48]),
    .sum(sum_19[48]));
  AL_FADD comp19_49 (
    .a(1'b0),
    .b(sum_18[49]),
    .c(cout_19[48]),
    .cout(cout_19[49]),
    .sum(sum_19[49]));
  AL_FADD comp19_5 (
    .a(i19[5]),
    .b(sum_18[5]),
    .c(cout_19[4]),
    .cout(cout_19[5]),
    .sum(sum_19[5]));
  AL_FADD comp19_50 (
    .a(1'b0),
    .b(sum_18[50]),
    .c(cout_19[49]),
    .cout(cout_19[50]),
    .sum(sum_19[50]));
  AL_FADD comp19_51 (
    .a(1'b0),
    .b(sum_18[51]),
    .c(cout_19[50]),
    .cout(cout_19[51]),
    .sum(sum_19[51]));
  AL_FADD comp19_52 (
    .a(1'b0),
    .b(sum_18[52]),
    .c(cout_19[51]),
    .cout(cout_19[52]),
    .sum(sum_19[52]));
  AL_FADD comp19_53 (
    .a(1'b0),
    .b(sum_18[53]),
    .c(cout_19[52]),
    .cout(cout_19[53]),
    .sum(sum_19[53]));
  AL_FADD comp19_54 (
    .a(1'b0),
    .b(sum_18[54]),
    .c(cout_19[53]),
    .cout(cout_19[54]),
    .sum(sum_19[54]));
  AL_FADD comp19_55 (
    .a(1'b0),
    .b(sum_18[55]),
    .c(cout_19[54]),
    .cout(cout_19[55]),
    .sum(sum_19[55]));
  AL_FADD comp19_56 (
    .a(1'b0),
    .b(sum_18[56]),
    .c(cout_19[55]),
    .cout(cout_19[56]),
    .sum(sum_19[56]));
  AL_FADD comp19_57 (
    .a(1'b0),
    .b(sum_18[57]),
    .c(cout_19[56]),
    .cout(cout_19[57]),
    .sum(sum_19[57]));
  AL_FADD comp19_58 (
    .a(1'b0),
    .b(sum_18[58]),
    .c(cout_19[57]),
    .cout(cout_19[58]),
    .sum(sum_19[58]));
  AL_FADD comp19_59 (
    .a(1'b0),
    .b(sum_18[59]),
    .c(cout_19[58]),
    .cout(cout_19[59]),
    .sum(sum_19[59]));
  AL_FADD comp19_6 (
    .a(i19[6]),
    .b(sum_18[6]),
    .c(cout_19[5]),
    .cout(cout_19[6]),
    .sum(sum_19[6]));
  AL_FADD comp19_60 (
    .a(1'b0),
    .b(sum_18[60]),
    .c(cout_19[59]),
    .cout(cout_19[60]),
    .sum(sum_19[60]));
  AL_FADD comp19_61 (
    .a(1'b0),
    .b(sum_18[61]),
    .c(cout_19[60]),
    .cout(cout_19[61]),
    .sum(sum_19[61]));
  AL_FADD comp19_62 (
    .a(1'b0),
    .b(sum_18[62]),
    .c(cout_19[61]),
    .cout(cout_19[62]),
    .sum(sum_19[62]));
  AL_FADD comp19_63 (
    .a(1'b0),
    .b(sum_18[63]),
    .c(cout_19[62]),
    .cout(cout_19[63]),
    .sum(sum_19[63]));
  AL_FADD comp19_7 (
    .a(i19[7]),
    .b(sum_18[7]),
    .c(cout_19[6]),
    .cout(cout_19[7]),
    .sum(sum_19[7]));
  AL_FADD comp19_8 (
    .a(i19[8]),
    .b(sum_18[8]),
    .c(cout_19[7]),
    .cout(cout_19[8]),
    .sum(sum_19[8]));
  AL_FADD comp19_9 (
    .a(i19[9]),
    .b(sum_18[9]),
    .c(cout_19[8]),
    .cout(cout_19[9]),
    .sum(sum_19[9]));
  AL_FADD comp1_0 (
    .a(i1[0]),
    .b(i0[0]),
    .c(1'b0),
    .cout(cout_1[0]),
    .sum(sum_1[0]));
  AL_FADD comp1_1 (
    .a(i1[1]),
    .b(i0[1]),
    .c(cout_1[0]),
    .cout(cout_1[1]),
    .sum(sum_1[1]));
  AL_FADD comp1_10 (
    .a(i1[10]),
    .b(i0[10]),
    .c(cout_1[9]),
    .cout(cout_1[10]),
    .sum(sum_1[10]));
  AL_FADD comp1_11 (
    .a(i1[11]),
    .b(i0[11]),
    .c(cout_1[10]),
    .cout(cout_1[11]),
    .sum(sum_1[11]));
  AL_FADD comp1_12 (
    .a(i1[12]),
    .b(i0[12]),
    .c(cout_1[11]),
    .cout(cout_1[12]),
    .sum(sum_1[12]));
  AL_FADD comp1_13 (
    .a(i1[13]),
    .b(i0[13]),
    .c(cout_1[12]),
    .cout(cout_1[13]),
    .sum(sum_1[13]));
  AL_FADD comp1_14 (
    .a(i1[14]),
    .b(i0[14]),
    .c(cout_1[13]),
    .cout(cout_1[14]),
    .sum(sum_1[14]));
  AL_FADD comp1_15 (
    .a(i1[15]),
    .b(i0[15]),
    .c(cout_1[14]),
    .cout(cout_1[15]),
    .sum(sum_1[15]));
  AL_FADD comp1_16 (
    .a(i1[16]),
    .b(i0[16]),
    .c(cout_1[15]),
    .cout(cout_1[16]),
    .sum(sum_1[16]));
  AL_FADD comp1_17 (
    .a(i1[17]),
    .b(i0[17]),
    .c(cout_1[16]),
    .cout(cout_1[17]),
    .sum(sum_1[17]));
  AL_FADD comp1_18 (
    .a(i1[18]),
    .b(i0[18]),
    .c(cout_1[17]),
    .cout(cout_1[18]),
    .sum(sum_1[18]));
  AL_FADD comp1_19 (
    .a(i1[19]),
    .b(i0[19]),
    .c(cout_1[18]),
    .cout(cout_1[19]),
    .sum(sum_1[19]));
  AL_FADD comp1_2 (
    .a(i1[2]),
    .b(i0[2]),
    .c(cout_1[1]),
    .cout(cout_1[2]),
    .sum(sum_1[2]));
  AL_FADD comp1_20 (
    .a(i1[20]),
    .b(i0[20]),
    .c(cout_1[19]),
    .cout(cout_1[20]),
    .sum(sum_1[20]));
  AL_FADD comp1_21 (
    .a(i1[21]),
    .b(i0[21]),
    .c(cout_1[20]),
    .cout(cout_1[21]),
    .sum(sum_1[21]));
  AL_FADD comp1_22 (
    .a(i1[22]),
    .b(i0[22]),
    .c(cout_1[21]),
    .cout(cout_1[22]),
    .sum(sum_1[22]));
  AL_FADD comp1_23 (
    .a(i1[23]),
    .b(i0[23]),
    .c(cout_1[22]),
    .cout(cout_1[23]),
    .sum(sum_1[23]));
  AL_FADD comp1_24 (
    .a(i1[24]),
    .b(i0[24]),
    .c(cout_1[23]),
    .cout(cout_1[24]),
    .sum(sum_1[24]));
  AL_FADD comp1_25 (
    .a(i1[25]),
    .b(i0[25]),
    .c(cout_1[24]),
    .cout(cout_1[25]),
    .sum(sum_1[25]));
  AL_FADD comp1_26 (
    .a(i1[26]),
    .b(i0[26]),
    .c(cout_1[25]),
    .cout(cout_1[26]),
    .sum(sum_1[26]));
  AL_FADD comp1_27 (
    .a(i1[27]),
    .b(i0[27]),
    .c(cout_1[26]),
    .cout(cout_1[27]),
    .sum(sum_1[27]));
  AL_FADD comp1_28 (
    .a(i1[28]),
    .b(i0[28]),
    .c(cout_1[27]),
    .cout(cout_1[28]),
    .sum(sum_1[28]));
  AL_FADD comp1_29 (
    .a(i1[29]),
    .b(i0[29]),
    .c(cout_1[28]),
    .cout(cout_1[29]),
    .sum(sum_1[29]));
  AL_FADD comp1_3 (
    .a(i1[3]),
    .b(i0[3]),
    .c(cout_1[2]),
    .cout(cout_1[3]),
    .sum(sum_1[3]));
  AL_FADD comp1_30 (
    .a(i1[30]),
    .b(i0[30]),
    .c(cout_1[29]),
    .cout(cout_1[30]),
    .sum(sum_1[30]));
  AL_FADD comp1_31 (
    .a(i1[31]),
    .b(i0[31]),
    .c(cout_1[30]),
    .cout(cout_1[31]),
    .sum(sum_1[31]));
  AL_FADD comp1_32 (
    .a(i1[32]),
    .b(i0[32]),
    .c(cout_1[31]),
    .cout(cout_1[32]),
    .sum(sum_1[32]));
  AL_FADD comp1_33 (
    .a(i1[33]),
    .b(i0[33]),
    .c(cout_1[32]),
    .cout(cout_1[33]),
    .sum(sum_1[33]));
  AL_FADD comp1_34 (
    .a(i1[34]),
    .b(i0[34]),
    .c(cout_1[33]),
    .cout(cout_1[34]),
    .sum(sum_1[34]));
  AL_FADD comp1_35 (
    .a(i1[35]),
    .b(i0[35]),
    .c(cout_1[34]),
    .cout(cout_1[35]),
    .sum(sum_1[35]));
  AL_FADD comp1_36 (
    .a(i1[36]),
    .b(i0[36]),
    .c(cout_1[35]),
    .cout(cout_1[36]),
    .sum(sum_1[36]));
  AL_FADD comp1_37 (
    .a(i1[37]),
    .b(i0[37]),
    .c(cout_1[36]),
    .cout(cout_1[37]),
    .sum(sum_1[37]));
  AL_FADD comp1_38 (
    .a(i1[38]),
    .b(i0[38]),
    .c(cout_1[37]),
    .cout(cout_1[38]),
    .sum(sum_1[38]));
  AL_FADD comp1_39 (
    .a(i1[39]),
    .b(i0[39]),
    .c(cout_1[38]),
    .cout(cout_1[39]),
    .sum(sum_1[39]));
  AL_FADD comp1_4 (
    .a(i1[4]),
    .b(i0[4]),
    .c(cout_1[3]),
    .cout(cout_1[4]),
    .sum(sum_1[4]));
  AL_FADD comp1_40 (
    .a(i1[40]),
    .b(i0[40]),
    .c(cout_1[39]),
    .cout(cout_1[40]),
    .sum(sum_1[40]));
  AL_FADD comp1_41 (
    .a(i1[41]),
    .b(i0[41]),
    .c(cout_1[40]),
    .cout(cout_1[41]),
    .sum(sum_1[41]));
  AL_FADD comp1_42 (
    .a(i1[42]),
    .b(i0[42]),
    .c(cout_1[41]),
    .cout(cout_1[42]),
    .sum(sum_1[42]));
  AL_FADD comp1_43 (
    .a(i1[43]),
    .b(i0[43]),
    .c(cout_1[42]),
    .cout(cout_1[43]),
    .sum(sum_1[43]));
  AL_FADD comp1_44 (
    .a(i1[44]),
    .b(i0[44]),
    .c(cout_1[43]),
    .cout(cout_1[44]),
    .sum(sum_1[44]));
  AL_FADD comp1_45 (
    .a(i1[45]),
    .b(i0[45]),
    .c(cout_1[44]),
    .cout(cout_1[45]),
    .sum(sum_1[45]));
  AL_FADD comp1_46 (
    .a(i1[46]),
    .b(i0[46]),
    .c(cout_1[45]),
    .cout(cout_1[46]),
    .sum(sum_1[46]));
  AL_FADD comp1_47 (
    .a(i1[47]),
    .b(i0[47]),
    .c(cout_1[46]),
    .cout(cout_1[47]),
    .sum(sum_1[47]));
  AL_FADD comp1_48 (
    .a(i1[48]),
    .b(i0[48]),
    .c(cout_1[47]),
    .cout(cout_1[48]),
    .sum(sum_1[48]));
  AL_FADD comp1_49 (
    .a(i1[49]),
    .b(i0[49]),
    .c(cout_1[48]),
    .cout(cout_1[49]),
    .sum(sum_1[49]));
  AL_FADD comp1_5 (
    .a(i1[5]),
    .b(i0[5]),
    .c(cout_1[4]),
    .cout(cout_1[5]),
    .sum(sum_1[5]));
  AL_FADD comp1_50 (
    .a(i1[50]),
    .b(i0[50]),
    .c(cout_1[49]),
    .cout(cout_1[50]),
    .sum(sum_1[50]));
  AL_FADD comp1_51 (
    .a(i1[51]),
    .b(i0[51]),
    .c(cout_1[50]),
    .cout(cout_1[51]),
    .sum(sum_1[51]));
  AL_FADD comp1_52 (
    .a(i1[52]),
    .b(i0[52]),
    .c(cout_1[51]),
    .cout(cout_1[52]),
    .sum(sum_1[52]));
  AL_FADD comp1_53 (
    .a(i1[53]),
    .b(i0[53]),
    .c(cout_1[52]),
    .cout(cout_1[53]),
    .sum(sum_1[53]));
  AL_FADD comp1_54 (
    .a(i1[54]),
    .b(i0[54]),
    .c(cout_1[53]),
    .cout(cout_1[54]),
    .sum(sum_1[54]));
  AL_FADD comp1_55 (
    .a(i1[55]),
    .b(i0[55]),
    .c(cout_1[54]),
    .cout(cout_1[55]),
    .sum(sum_1[55]));
  AL_FADD comp1_56 (
    .a(i1[56]),
    .b(i0[56]),
    .c(cout_1[55]),
    .cout(cout_1[56]),
    .sum(sum_1[56]));
  AL_FADD comp1_57 (
    .a(i1[57]),
    .b(i0[57]),
    .c(cout_1[56]),
    .cout(cout_1[57]),
    .sum(sum_1[57]));
  AL_FADD comp1_58 (
    .a(i1[58]),
    .b(i0[58]),
    .c(cout_1[57]),
    .cout(cout_1[58]),
    .sum(sum_1[58]));
  AL_FADD comp1_59 (
    .a(i1[59]),
    .b(i0[59]),
    .c(cout_1[58]),
    .cout(cout_1[59]),
    .sum(sum_1[59]));
  AL_FADD comp1_6 (
    .a(i1[6]),
    .b(i0[6]),
    .c(cout_1[5]),
    .cout(cout_1[6]),
    .sum(sum_1[6]));
  AL_FADD comp1_60 (
    .a(1'b0),
    .b(i0[60]),
    .c(cout_1[59]),
    .cout(cout_1[60]),
    .sum(sum_1[60]));
  AL_FADD comp1_61 (
    .a(1'b0),
    .b(i0[61]),
    .c(cout_1[60]),
    .cout(cout_1[61]),
    .sum(sum_1[61]));
  AL_FADD comp1_62 (
    .a(1'b0),
    .b(i0[62]),
    .c(cout_1[61]),
    .cout(cout_1[62]),
    .sum(sum_1[62]));
  AL_FADD comp1_7 (
    .a(i1[7]),
    .b(i0[7]),
    .c(cout_1[6]),
    .cout(cout_1[7]),
    .sum(sum_1[7]));
  AL_FADD comp1_8 (
    .a(i1[8]),
    .b(i0[8]),
    .c(cout_1[7]),
    .cout(cout_1[8]),
    .sum(sum_1[8]));
  AL_FADD comp1_9 (
    .a(i1[9]),
    .b(i0[9]),
    .c(cout_1[8]),
    .cout(cout_1[9]),
    .sum(sum_1[9]));
  AL_FADD comp20_0 (
    .a(i20[0]),
    .b(sum_19[0]),
    .c(1'b0),
    .cout(cout_20[0]),
    .sum(sum_20[0]));
  AL_FADD comp20_1 (
    .a(i20[1]),
    .b(sum_19[1]),
    .c(cout_20[0]),
    .cout(cout_20[1]),
    .sum(sum_20[1]));
  AL_FADD comp20_10 (
    .a(i20[10]),
    .b(sum_19[10]),
    .c(cout_20[9]),
    .cout(cout_20[10]),
    .sum(sum_20[10]));
  AL_FADD comp20_11 (
    .a(i20[11]),
    .b(sum_19[11]),
    .c(cout_20[10]),
    .cout(cout_20[11]),
    .sum(sum_20[11]));
  AL_FADD comp20_12 (
    .a(i20[12]),
    .b(sum_19[12]),
    .c(cout_20[11]),
    .cout(cout_20[12]),
    .sum(sum_20[12]));
  AL_FADD comp20_13 (
    .a(i20[13]),
    .b(sum_19[13]),
    .c(cout_20[12]),
    .cout(cout_20[13]),
    .sum(sum_20[13]));
  AL_FADD comp20_14 (
    .a(i20[14]),
    .b(sum_19[14]),
    .c(cout_20[13]),
    .cout(cout_20[14]),
    .sum(sum_20[14]));
  AL_FADD comp20_15 (
    .a(i20[15]),
    .b(sum_19[15]),
    .c(cout_20[14]),
    .cout(cout_20[15]),
    .sum(sum_20[15]));
  AL_FADD comp20_16 (
    .a(i20[16]),
    .b(sum_19[16]),
    .c(cout_20[15]),
    .cout(cout_20[16]),
    .sum(sum_20[16]));
  AL_FADD comp20_17 (
    .a(i20[17]),
    .b(sum_19[17]),
    .c(cout_20[16]),
    .cout(cout_20[17]),
    .sum(sum_20[17]));
  AL_FADD comp20_18 (
    .a(i20[18]),
    .b(sum_19[18]),
    .c(cout_20[17]),
    .cout(cout_20[18]),
    .sum(sum_20[18]));
  AL_FADD comp20_19 (
    .a(i20[19]),
    .b(sum_19[19]),
    .c(cout_20[18]),
    .cout(cout_20[19]),
    .sum(sum_20[19]));
  AL_FADD comp20_2 (
    .a(i20[2]),
    .b(sum_19[2]),
    .c(cout_20[1]),
    .cout(cout_20[2]),
    .sum(sum_20[2]));
  AL_FADD comp20_20 (
    .a(i20[20]),
    .b(sum_19[20]),
    .c(cout_20[19]),
    .cout(cout_20[20]),
    .sum(sum_20[20]));
  AL_FADD comp20_21 (
    .a(i20[21]),
    .b(sum_19[21]),
    .c(cout_20[20]),
    .cout(cout_20[21]),
    .sum(sum_20[21]));
  AL_FADD comp20_22 (
    .a(i20[22]),
    .b(sum_19[22]),
    .c(cout_20[21]),
    .cout(cout_20[22]),
    .sum(sum_20[22]));
  AL_FADD comp20_23 (
    .a(i20[23]),
    .b(sum_19[23]),
    .c(cout_20[22]),
    .cout(cout_20[23]),
    .sum(sum_20[23]));
  AL_FADD comp20_24 (
    .a(i20[24]),
    .b(sum_19[24]),
    .c(cout_20[23]),
    .cout(cout_20[24]),
    .sum(sum_20[24]));
  AL_FADD comp20_25 (
    .a(i20[25]),
    .b(sum_19[25]),
    .c(cout_20[24]),
    .cout(cout_20[25]),
    .sum(sum_20[25]));
  AL_FADD comp20_26 (
    .a(i20[26]),
    .b(sum_19[26]),
    .c(cout_20[25]),
    .cout(cout_20[26]),
    .sum(sum_20[26]));
  AL_FADD comp20_27 (
    .a(i20[27]),
    .b(sum_19[27]),
    .c(cout_20[26]),
    .cout(cout_20[27]),
    .sum(sum_20[27]));
  AL_FADD comp20_28 (
    .a(i20[28]),
    .b(sum_19[28]),
    .c(cout_20[27]),
    .cout(cout_20[28]),
    .sum(sum_20[28]));
  AL_FADD comp20_29 (
    .a(i20[29]),
    .b(sum_19[29]),
    .c(cout_20[28]),
    .cout(cout_20[29]),
    .sum(sum_20[29]));
  AL_FADD comp20_3 (
    .a(i20[3]),
    .b(sum_19[3]),
    .c(cout_20[2]),
    .cout(cout_20[3]),
    .sum(sum_20[3]));
  AL_FADD comp20_30 (
    .a(i20[30]),
    .b(sum_19[30]),
    .c(cout_20[29]),
    .cout(cout_20[30]),
    .sum(sum_20[30]));
  AL_FADD comp20_31 (
    .a(i20[31]),
    .b(sum_19[31]),
    .c(cout_20[30]),
    .cout(cout_20[31]),
    .sum(sum_20[31]));
  AL_FADD comp20_32 (
    .a(i20[32]),
    .b(sum_19[32]),
    .c(cout_20[31]),
    .cout(cout_20[32]),
    .sum(sum_20[32]));
  AL_FADD comp20_33 (
    .a(i20[33]),
    .b(sum_19[33]),
    .c(cout_20[32]),
    .cout(cout_20[33]),
    .sum(sum_20[33]));
  AL_FADD comp20_34 (
    .a(i20[34]),
    .b(sum_19[34]),
    .c(cout_20[33]),
    .cout(cout_20[34]),
    .sum(sum_20[34]));
  AL_FADD comp20_35 (
    .a(i20[35]),
    .b(sum_19[35]),
    .c(cout_20[34]),
    .cout(cout_20[35]),
    .sum(sum_20[35]));
  AL_FADD comp20_36 (
    .a(i20[36]),
    .b(sum_19[36]),
    .c(cout_20[35]),
    .cout(cout_20[36]),
    .sum(sum_20[36]));
  AL_FADD comp20_37 (
    .a(i20[37]),
    .b(sum_19[37]),
    .c(cout_20[36]),
    .cout(cout_20[37]),
    .sum(sum_20[37]));
  AL_FADD comp20_38 (
    .a(i20[38]),
    .b(sum_19[38]),
    .c(cout_20[37]),
    .cout(cout_20[38]),
    .sum(sum_20[38]));
  AL_FADD comp20_39 (
    .a(i20[39]),
    .b(sum_19[39]),
    .c(cout_20[38]),
    .cout(cout_20[39]),
    .sum(sum_20[39]));
  AL_FADD comp20_4 (
    .a(i20[4]),
    .b(sum_19[4]),
    .c(cout_20[3]),
    .cout(cout_20[4]),
    .sum(sum_20[4]));
  AL_FADD comp20_40 (
    .a(i20[40]),
    .b(sum_19[40]),
    .c(cout_20[39]),
    .cout(cout_20[40]),
    .sum(sum_20[40]));
  AL_FADD comp20_41 (
    .a(1'b0),
    .b(sum_19[41]),
    .c(cout_20[40]),
    .cout(cout_20[41]),
    .sum(sum_20[41]));
  AL_FADD comp20_42 (
    .a(1'b0),
    .b(sum_19[42]),
    .c(cout_20[41]),
    .cout(cout_20[42]),
    .sum(sum_20[42]));
  AL_FADD comp20_43 (
    .a(1'b0),
    .b(sum_19[43]),
    .c(cout_20[42]),
    .cout(cout_20[43]),
    .sum(sum_20[43]));
  AL_FADD comp20_44 (
    .a(1'b0),
    .b(sum_19[44]),
    .c(cout_20[43]),
    .cout(cout_20[44]),
    .sum(sum_20[44]));
  AL_FADD comp20_45 (
    .a(1'b0),
    .b(sum_19[45]),
    .c(cout_20[44]),
    .cout(cout_20[45]),
    .sum(sum_20[45]));
  AL_FADD comp20_46 (
    .a(1'b0),
    .b(sum_19[46]),
    .c(cout_20[45]),
    .cout(cout_20[46]),
    .sum(sum_20[46]));
  AL_FADD comp20_47 (
    .a(1'b0),
    .b(sum_19[47]),
    .c(cout_20[46]),
    .cout(cout_20[47]),
    .sum(sum_20[47]));
  AL_FADD comp20_48 (
    .a(1'b0),
    .b(sum_19[48]),
    .c(cout_20[47]),
    .cout(cout_20[48]),
    .sum(sum_20[48]));
  AL_FADD comp20_49 (
    .a(1'b0),
    .b(sum_19[49]),
    .c(cout_20[48]),
    .cout(cout_20[49]),
    .sum(sum_20[49]));
  AL_FADD comp20_5 (
    .a(i20[5]),
    .b(sum_19[5]),
    .c(cout_20[4]),
    .cout(cout_20[5]),
    .sum(sum_20[5]));
  AL_FADD comp20_50 (
    .a(1'b0),
    .b(sum_19[50]),
    .c(cout_20[49]),
    .cout(cout_20[50]),
    .sum(sum_20[50]));
  AL_FADD comp20_51 (
    .a(1'b0),
    .b(sum_19[51]),
    .c(cout_20[50]),
    .cout(cout_20[51]),
    .sum(sum_20[51]));
  AL_FADD comp20_52 (
    .a(1'b0),
    .b(sum_19[52]),
    .c(cout_20[51]),
    .cout(cout_20[52]),
    .sum(sum_20[52]));
  AL_FADD comp20_53 (
    .a(1'b0),
    .b(sum_19[53]),
    .c(cout_20[52]),
    .cout(cout_20[53]),
    .sum(sum_20[53]));
  AL_FADD comp20_54 (
    .a(1'b0),
    .b(sum_19[54]),
    .c(cout_20[53]),
    .cout(cout_20[54]),
    .sum(sum_20[54]));
  AL_FADD comp20_55 (
    .a(1'b0),
    .b(sum_19[55]),
    .c(cout_20[54]),
    .cout(cout_20[55]),
    .sum(sum_20[55]));
  AL_FADD comp20_56 (
    .a(1'b0),
    .b(sum_19[56]),
    .c(cout_20[55]),
    .cout(cout_20[56]),
    .sum(sum_20[56]));
  AL_FADD comp20_57 (
    .a(1'b0),
    .b(sum_19[57]),
    .c(cout_20[56]),
    .cout(cout_20[57]),
    .sum(sum_20[57]));
  AL_FADD comp20_58 (
    .a(1'b0),
    .b(sum_19[58]),
    .c(cout_20[57]),
    .cout(cout_20[58]),
    .sum(sum_20[58]));
  AL_FADD comp20_59 (
    .a(1'b0),
    .b(sum_19[59]),
    .c(cout_20[58]),
    .cout(cout_20[59]),
    .sum(sum_20[59]));
  AL_FADD comp20_6 (
    .a(i20[6]),
    .b(sum_19[6]),
    .c(cout_20[5]),
    .cout(cout_20[6]),
    .sum(sum_20[6]));
  AL_FADD comp20_60 (
    .a(1'b0),
    .b(sum_19[60]),
    .c(cout_20[59]),
    .cout(cout_20[60]),
    .sum(sum_20[60]));
  AL_FADD comp20_61 (
    .a(1'b0),
    .b(sum_19[61]),
    .c(cout_20[60]),
    .cout(cout_20[61]),
    .sum(sum_20[61]));
  AL_FADD comp20_62 (
    .a(1'b0),
    .b(sum_19[62]),
    .c(cout_20[61]),
    .cout(cout_20[62]),
    .sum(sum_20[62]));
  AL_FADD comp20_63 (
    .a(1'b0),
    .b(sum_19[63]),
    .c(cout_20[62]),
    .cout(cout_20[63]),
    .sum(sum_20[63]));
  AL_FADD comp20_7 (
    .a(i20[7]),
    .b(sum_19[7]),
    .c(cout_20[6]),
    .cout(cout_20[7]),
    .sum(sum_20[7]));
  AL_FADD comp20_8 (
    .a(i20[8]),
    .b(sum_19[8]),
    .c(cout_20[7]),
    .cout(cout_20[8]),
    .sum(sum_20[8]));
  AL_FADD comp20_9 (
    .a(i20[9]),
    .b(sum_19[9]),
    .c(cout_20[8]),
    .cout(cout_20[9]),
    .sum(sum_20[9]));
  AL_FADD comp21_0 (
    .a(i21[0]),
    .b(sum_20[0]),
    .c(1'b0),
    .cout(cout_21[0]),
    .sum(sum_21[0]));
  AL_FADD comp21_1 (
    .a(i21[1]),
    .b(sum_20[1]),
    .c(cout_21[0]),
    .cout(cout_21[1]),
    .sum(sum_21[1]));
  AL_FADD comp21_10 (
    .a(i21[10]),
    .b(sum_20[10]),
    .c(cout_21[9]),
    .cout(cout_21[10]),
    .sum(sum_21[10]));
  AL_FADD comp21_11 (
    .a(i21[11]),
    .b(sum_20[11]),
    .c(cout_21[10]),
    .cout(cout_21[11]),
    .sum(sum_21[11]));
  AL_FADD comp21_12 (
    .a(i21[12]),
    .b(sum_20[12]),
    .c(cout_21[11]),
    .cout(cout_21[12]),
    .sum(sum_21[12]));
  AL_FADD comp21_13 (
    .a(i21[13]),
    .b(sum_20[13]),
    .c(cout_21[12]),
    .cout(cout_21[13]),
    .sum(sum_21[13]));
  AL_FADD comp21_14 (
    .a(i21[14]),
    .b(sum_20[14]),
    .c(cout_21[13]),
    .cout(cout_21[14]),
    .sum(sum_21[14]));
  AL_FADD comp21_15 (
    .a(i21[15]),
    .b(sum_20[15]),
    .c(cout_21[14]),
    .cout(cout_21[15]),
    .sum(sum_21[15]));
  AL_FADD comp21_16 (
    .a(i21[16]),
    .b(sum_20[16]),
    .c(cout_21[15]),
    .cout(cout_21[16]),
    .sum(sum_21[16]));
  AL_FADD comp21_17 (
    .a(i21[17]),
    .b(sum_20[17]),
    .c(cout_21[16]),
    .cout(cout_21[17]),
    .sum(sum_21[17]));
  AL_FADD comp21_18 (
    .a(i21[18]),
    .b(sum_20[18]),
    .c(cout_21[17]),
    .cout(cout_21[18]),
    .sum(sum_21[18]));
  AL_FADD comp21_19 (
    .a(i21[19]),
    .b(sum_20[19]),
    .c(cout_21[18]),
    .cout(cout_21[19]),
    .sum(sum_21[19]));
  AL_FADD comp21_2 (
    .a(i21[2]),
    .b(sum_20[2]),
    .c(cout_21[1]),
    .cout(cout_21[2]),
    .sum(sum_21[2]));
  AL_FADD comp21_20 (
    .a(i21[20]),
    .b(sum_20[20]),
    .c(cout_21[19]),
    .cout(cout_21[20]),
    .sum(sum_21[20]));
  AL_FADD comp21_21 (
    .a(i21[21]),
    .b(sum_20[21]),
    .c(cout_21[20]),
    .cout(cout_21[21]),
    .sum(sum_21[21]));
  AL_FADD comp21_22 (
    .a(i21[22]),
    .b(sum_20[22]),
    .c(cout_21[21]),
    .cout(cout_21[22]),
    .sum(sum_21[22]));
  AL_FADD comp21_23 (
    .a(i21[23]),
    .b(sum_20[23]),
    .c(cout_21[22]),
    .cout(cout_21[23]),
    .sum(sum_21[23]));
  AL_FADD comp21_24 (
    .a(i21[24]),
    .b(sum_20[24]),
    .c(cout_21[23]),
    .cout(cout_21[24]),
    .sum(sum_21[24]));
  AL_FADD comp21_25 (
    .a(i21[25]),
    .b(sum_20[25]),
    .c(cout_21[24]),
    .cout(cout_21[25]),
    .sum(sum_21[25]));
  AL_FADD comp21_26 (
    .a(i21[26]),
    .b(sum_20[26]),
    .c(cout_21[25]),
    .cout(cout_21[26]),
    .sum(sum_21[26]));
  AL_FADD comp21_27 (
    .a(i21[27]),
    .b(sum_20[27]),
    .c(cout_21[26]),
    .cout(cout_21[27]),
    .sum(sum_21[27]));
  AL_FADD comp21_28 (
    .a(i21[28]),
    .b(sum_20[28]),
    .c(cout_21[27]),
    .cout(cout_21[28]),
    .sum(sum_21[28]));
  AL_FADD comp21_29 (
    .a(i21[29]),
    .b(sum_20[29]),
    .c(cout_21[28]),
    .cout(cout_21[29]),
    .sum(sum_21[29]));
  AL_FADD comp21_3 (
    .a(i21[3]),
    .b(sum_20[3]),
    .c(cout_21[2]),
    .cout(cout_21[3]),
    .sum(sum_21[3]));
  AL_FADD comp21_30 (
    .a(i21[30]),
    .b(sum_20[30]),
    .c(cout_21[29]),
    .cout(cout_21[30]),
    .sum(sum_21[30]));
  AL_FADD comp21_31 (
    .a(i21[31]),
    .b(sum_20[31]),
    .c(cout_21[30]),
    .cout(cout_21[31]),
    .sum(sum_21[31]));
  AL_FADD comp21_32 (
    .a(i21[32]),
    .b(sum_20[32]),
    .c(cout_21[31]),
    .cout(cout_21[32]),
    .sum(sum_21[32]));
  AL_FADD comp21_33 (
    .a(i21[33]),
    .b(sum_20[33]),
    .c(cout_21[32]),
    .cout(cout_21[33]),
    .sum(sum_21[33]));
  AL_FADD comp21_34 (
    .a(i21[34]),
    .b(sum_20[34]),
    .c(cout_21[33]),
    .cout(cout_21[34]),
    .sum(sum_21[34]));
  AL_FADD comp21_35 (
    .a(i21[35]),
    .b(sum_20[35]),
    .c(cout_21[34]),
    .cout(cout_21[35]),
    .sum(sum_21[35]));
  AL_FADD comp21_36 (
    .a(i21[36]),
    .b(sum_20[36]),
    .c(cout_21[35]),
    .cout(cout_21[36]),
    .sum(sum_21[36]));
  AL_FADD comp21_37 (
    .a(i21[37]),
    .b(sum_20[37]),
    .c(cout_21[36]),
    .cout(cout_21[37]),
    .sum(sum_21[37]));
  AL_FADD comp21_38 (
    .a(i21[38]),
    .b(sum_20[38]),
    .c(cout_21[37]),
    .cout(cout_21[38]),
    .sum(sum_21[38]));
  AL_FADD comp21_39 (
    .a(i21[39]),
    .b(sum_20[39]),
    .c(cout_21[38]),
    .cout(cout_21[39]),
    .sum(sum_21[39]));
  AL_FADD comp21_4 (
    .a(i21[4]),
    .b(sum_20[4]),
    .c(cout_21[3]),
    .cout(cout_21[4]),
    .sum(sum_21[4]));
  AL_FADD comp21_40 (
    .a(1'b0),
    .b(sum_20[40]),
    .c(cout_21[39]),
    .cout(cout_21[40]),
    .sum(sum_21[40]));
  AL_FADD comp21_41 (
    .a(1'b0),
    .b(sum_20[41]),
    .c(cout_21[40]),
    .cout(cout_21[41]),
    .sum(sum_21[41]));
  AL_FADD comp21_42 (
    .a(1'b0),
    .b(sum_20[42]),
    .c(cout_21[41]),
    .cout(cout_21[42]),
    .sum(sum_21[42]));
  AL_FADD comp21_43 (
    .a(1'b0),
    .b(sum_20[43]),
    .c(cout_21[42]),
    .cout(cout_21[43]),
    .sum(sum_21[43]));
  AL_FADD comp21_44 (
    .a(1'b0),
    .b(sum_20[44]),
    .c(cout_21[43]),
    .cout(cout_21[44]),
    .sum(sum_21[44]));
  AL_FADD comp21_45 (
    .a(1'b0),
    .b(sum_20[45]),
    .c(cout_21[44]),
    .cout(cout_21[45]),
    .sum(sum_21[45]));
  AL_FADD comp21_46 (
    .a(1'b0),
    .b(sum_20[46]),
    .c(cout_21[45]),
    .cout(cout_21[46]),
    .sum(sum_21[46]));
  AL_FADD comp21_47 (
    .a(1'b0),
    .b(sum_20[47]),
    .c(cout_21[46]),
    .cout(cout_21[47]),
    .sum(sum_21[47]));
  AL_FADD comp21_48 (
    .a(1'b0),
    .b(sum_20[48]),
    .c(cout_21[47]),
    .cout(cout_21[48]),
    .sum(sum_21[48]));
  AL_FADD comp21_49 (
    .a(1'b0),
    .b(sum_20[49]),
    .c(cout_21[48]),
    .cout(cout_21[49]),
    .sum(sum_21[49]));
  AL_FADD comp21_5 (
    .a(i21[5]),
    .b(sum_20[5]),
    .c(cout_21[4]),
    .cout(cout_21[5]),
    .sum(sum_21[5]));
  AL_FADD comp21_50 (
    .a(1'b0),
    .b(sum_20[50]),
    .c(cout_21[49]),
    .cout(cout_21[50]),
    .sum(sum_21[50]));
  AL_FADD comp21_51 (
    .a(1'b0),
    .b(sum_20[51]),
    .c(cout_21[50]),
    .cout(cout_21[51]),
    .sum(sum_21[51]));
  AL_FADD comp21_52 (
    .a(1'b0),
    .b(sum_20[52]),
    .c(cout_21[51]),
    .cout(cout_21[52]),
    .sum(sum_21[52]));
  AL_FADD comp21_53 (
    .a(1'b0),
    .b(sum_20[53]),
    .c(cout_21[52]),
    .cout(cout_21[53]),
    .sum(sum_21[53]));
  AL_FADD comp21_54 (
    .a(1'b0),
    .b(sum_20[54]),
    .c(cout_21[53]),
    .cout(cout_21[54]),
    .sum(sum_21[54]));
  AL_FADD comp21_55 (
    .a(1'b0),
    .b(sum_20[55]),
    .c(cout_21[54]),
    .cout(cout_21[55]),
    .sum(sum_21[55]));
  AL_FADD comp21_56 (
    .a(1'b0),
    .b(sum_20[56]),
    .c(cout_21[55]),
    .cout(cout_21[56]),
    .sum(sum_21[56]));
  AL_FADD comp21_57 (
    .a(1'b0),
    .b(sum_20[57]),
    .c(cout_21[56]),
    .cout(cout_21[57]),
    .sum(sum_21[57]));
  AL_FADD comp21_58 (
    .a(1'b0),
    .b(sum_20[58]),
    .c(cout_21[57]),
    .cout(cout_21[58]),
    .sum(sum_21[58]));
  AL_FADD comp21_59 (
    .a(1'b0),
    .b(sum_20[59]),
    .c(cout_21[58]),
    .cout(cout_21[59]),
    .sum(sum_21[59]));
  AL_FADD comp21_6 (
    .a(i21[6]),
    .b(sum_20[6]),
    .c(cout_21[5]),
    .cout(cout_21[6]),
    .sum(sum_21[6]));
  AL_FADD comp21_60 (
    .a(1'b0),
    .b(sum_20[60]),
    .c(cout_21[59]),
    .cout(cout_21[60]),
    .sum(sum_21[60]));
  AL_FADD comp21_61 (
    .a(1'b0),
    .b(sum_20[61]),
    .c(cout_21[60]),
    .cout(cout_21[61]),
    .sum(sum_21[61]));
  AL_FADD comp21_62 (
    .a(1'b0),
    .b(sum_20[62]),
    .c(cout_21[61]),
    .cout(cout_21[62]),
    .sum(sum_21[62]));
  AL_FADD comp21_63 (
    .a(1'b0),
    .b(sum_20[63]),
    .c(cout_21[62]),
    .cout(cout_21[63]),
    .sum(sum_21[63]));
  AL_FADD comp21_7 (
    .a(i21[7]),
    .b(sum_20[7]),
    .c(cout_21[6]),
    .cout(cout_21[7]),
    .sum(sum_21[7]));
  AL_FADD comp21_8 (
    .a(i21[8]),
    .b(sum_20[8]),
    .c(cout_21[7]),
    .cout(cout_21[8]),
    .sum(sum_21[8]));
  AL_FADD comp21_9 (
    .a(i21[9]),
    .b(sum_20[9]),
    .c(cout_21[8]),
    .cout(cout_21[9]),
    .sum(sum_21[9]));
  AL_FADD comp22_0 (
    .a(i22[0]),
    .b(sum_21[0]),
    .c(1'b0),
    .cout(cout_22[0]),
    .sum(sum_22[0]));
  AL_FADD comp22_1 (
    .a(i22[1]),
    .b(sum_21[1]),
    .c(cout_22[0]),
    .cout(cout_22[1]),
    .sum(sum_22[1]));
  AL_FADD comp22_10 (
    .a(i22[10]),
    .b(sum_21[10]),
    .c(cout_22[9]),
    .cout(cout_22[10]),
    .sum(sum_22[10]));
  AL_FADD comp22_11 (
    .a(i22[11]),
    .b(sum_21[11]),
    .c(cout_22[10]),
    .cout(cout_22[11]),
    .sum(sum_22[11]));
  AL_FADD comp22_12 (
    .a(i22[12]),
    .b(sum_21[12]),
    .c(cout_22[11]),
    .cout(cout_22[12]),
    .sum(sum_22[12]));
  AL_FADD comp22_13 (
    .a(i22[13]),
    .b(sum_21[13]),
    .c(cout_22[12]),
    .cout(cout_22[13]),
    .sum(sum_22[13]));
  AL_FADD comp22_14 (
    .a(i22[14]),
    .b(sum_21[14]),
    .c(cout_22[13]),
    .cout(cout_22[14]),
    .sum(sum_22[14]));
  AL_FADD comp22_15 (
    .a(i22[15]),
    .b(sum_21[15]),
    .c(cout_22[14]),
    .cout(cout_22[15]),
    .sum(sum_22[15]));
  AL_FADD comp22_16 (
    .a(i22[16]),
    .b(sum_21[16]),
    .c(cout_22[15]),
    .cout(cout_22[16]),
    .sum(sum_22[16]));
  AL_FADD comp22_17 (
    .a(i22[17]),
    .b(sum_21[17]),
    .c(cout_22[16]),
    .cout(cout_22[17]),
    .sum(sum_22[17]));
  AL_FADD comp22_18 (
    .a(i22[18]),
    .b(sum_21[18]),
    .c(cout_22[17]),
    .cout(cout_22[18]),
    .sum(sum_22[18]));
  AL_FADD comp22_19 (
    .a(i22[19]),
    .b(sum_21[19]),
    .c(cout_22[18]),
    .cout(cout_22[19]),
    .sum(sum_22[19]));
  AL_FADD comp22_2 (
    .a(i22[2]),
    .b(sum_21[2]),
    .c(cout_22[1]),
    .cout(cout_22[2]),
    .sum(sum_22[2]));
  AL_FADD comp22_20 (
    .a(i22[20]),
    .b(sum_21[20]),
    .c(cout_22[19]),
    .cout(cout_22[20]),
    .sum(sum_22[20]));
  AL_FADD comp22_21 (
    .a(i22[21]),
    .b(sum_21[21]),
    .c(cout_22[20]),
    .cout(cout_22[21]),
    .sum(sum_22[21]));
  AL_FADD comp22_22 (
    .a(i22[22]),
    .b(sum_21[22]),
    .c(cout_22[21]),
    .cout(cout_22[22]),
    .sum(sum_22[22]));
  AL_FADD comp22_23 (
    .a(i22[23]),
    .b(sum_21[23]),
    .c(cout_22[22]),
    .cout(cout_22[23]),
    .sum(sum_22[23]));
  AL_FADD comp22_24 (
    .a(i22[24]),
    .b(sum_21[24]),
    .c(cout_22[23]),
    .cout(cout_22[24]),
    .sum(sum_22[24]));
  AL_FADD comp22_25 (
    .a(i22[25]),
    .b(sum_21[25]),
    .c(cout_22[24]),
    .cout(cout_22[25]),
    .sum(sum_22[25]));
  AL_FADD comp22_26 (
    .a(i22[26]),
    .b(sum_21[26]),
    .c(cout_22[25]),
    .cout(cout_22[26]),
    .sum(sum_22[26]));
  AL_FADD comp22_27 (
    .a(i22[27]),
    .b(sum_21[27]),
    .c(cout_22[26]),
    .cout(cout_22[27]),
    .sum(sum_22[27]));
  AL_FADD comp22_28 (
    .a(i22[28]),
    .b(sum_21[28]),
    .c(cout_22[27]),
    .cout(cout_22[28]),
    .sum(sum_22[28]));
  AL_FADD comp22_29 (
    .a(i22[29]),
    .b(sum_21[29]),
    .c(cout_22[28]),
    .cout(cout_22[29]),
    .sum(sum_22[29]));
  AL_FADD comp22_3 (
    .a(i22[3]),
    .b(sum_21[3]),
    .c(cout_22[2]),
    .cout(cout_22[3]),
    .sum(sum_22[3]));
  AL_FADD comp22_30 (
    .a(i22[30]),
    .b(sum_21[30]),
    .c(cout_22[29]),
    .cout(cout_22[30]),
    .sum(sum_22[30]));
  AL_FADD comp22_31 (
    .a(i22[31]),
    .b(sum_21[31]),
    .c(cout_22[30]),
    .cout(cout_22[31]),
    .sum(sum_22[31]));
  AL_FADD comp22_32 (
    .a(i22[32]),
    .b(sum_21[32]),
    .c(cout_22[31]),
    .cout(cout_22[32]),
    .sum(sum_22[32]));
  AL_FADD comp22_33 (
    .a(i22[33]),
    .b(sum_21[33]),
    .c(cout_22[32]),
    .cout(cout_22[33]),
    .sum(sum_22[33]));
  AL_FADD comp22_34 (
    .a(i22[34]),
    .b(sum_21[34]),
    .c(cout_22[33]),
    .cout(cout_22[34]),
    .sum(sum_22[34]));
  AL_FADD comp22_35 (
    .a(i22[35]),
    .b(sum_21[35]),
    .c(cout_22[34]),
    .cout(cout_22[35]),
    .sum(sum_22[35]));
  AL_FADD comp22_36 (
    .a(i22[36]),
    .b(sum_21[36]),
    .c(cout_22[35]),
    .cout(cout_22[36]),
    .sum(sum_22[36]));
  AL_FADD comp22_37 (
    .a(i22[37]),
    .b(sum_21[37]),
    .c(cout_22[36]),
    .cout(cout_22[37]),
    .sum(sum_22[37]));
  AL_FADD comp22_38 (
    .a(i22[38]),
    .b(sum_21[38]),
    .c(cout_22[37]),
    .cout(cout_22[38]),
    .sum(sum_22[38]));
  AL_FADD comp22_39 (
    .a(1'b0),
    .b(sum_21[39]),
    .c(cout_22[38]),
    .cout(cout_22[39]),
    .sum(sum_22[39]));
  AL_FADD comp22_4 (
    .a(i22[4]),
    .b(sum_21[4]),
    .c(cout_22[3]),
    .cout(cout_22[4]),
    .sum(sum_22[4]));
  AL_FADD comp22_40 (
    .a(1'b0),
    .b(sum_21[40]),
    .c(cout_22[39]),
    .cout(cout_22[40]),
    .sum(sum_22[40]));
  AL_FADD comp22_41 (
    .a(1'b0),
    .b(sum_21[41]),
    .c(cout_22[40]),
    .cout(cout_22[41]),
    .sum(sum_22[41]));
  AL_FADD comp22_42 (
    .a(1'b0),
    .b(sum_21[42]),
    .c(cout_22[41]),
    .cout(cout_22[42]),
    .sum(sum_22[42]));
  AL_FADD comp22_43 (
    .a(1'b0),
    .b(sum_21[43]),
    .c(cout_22[42]),
    .cout(cout_22[43]),
    .sum(sum_22[43]));
  AL_FADD comp22_44 (
    .a(1'b0),
    .b(sum_21[44]),
    .c(cout_22[43]),
    .cout(cout_22[44]),
    .sum(sum_22[44]));
  AL_FADD comp22_45 (
    .a(1'b0),
    .b(sum_21[45]),
    .c(cout_22[44]),
    .cout(cout_22[45]),
    .sum(sum_22[45]));
  AL_FADD comp22_46 (
    .a(1'b0),
    .b(sum_21[46]),
    .c(cout_22[45]),
    .cout(cout_22[46]),
    .sum(sum_22[46]));
  AL_FADD comp22_47 (
    .a(1'b0),
    .b(sum_21[47]),
    .c(cout_22[46]),
    .cout(cout_22[47]),
    .sum(sum_22[47]));
  AL_FADD comp22_48 (
    .a(1'b0),
    .b(sum_21[48]),
    .c(cout_22[47]),
    .cout(cout_22[48]),
    .sum(sum_22[48]));
  AL_FADD comp22_49 (
    .a(1'b0),
    .b(sum_21[49]),
    .c(cout_22[48]),
    .cout(cout_22[49]),
    .sum(sum_22[49]));
  AL_FADD comp22_5 (
    .a(i22[5]),
    .b(sum_21[5]),
    .c(cout_22[4]),
    .cout(cout_22[5]),
    .sum(sum_22[5]));
  AL_FADD comp22_50 (
    .a(1'b0),
    .b(sum_21[50]),
    .c(cout_22[49]),
    .cout(cout_22[50]),
    .sum(sum_22[50]));
  AL_FADD comp22_51 (
    .a(1'b0),
    .b(sum_21[51]),
    .c(cout_22[50]),
    .cout(cout_22[51]),
    .sum(sum_22[51]));
  AL_FADD comp22_52 (
    .a(1'b0),
    .b(sum_21[52]),
    .c(cout_22[51]),
    .cout(cout_22[52]),
    .sum(sum_22[52]));
  AL_FADD comp22_53 (
    .a(1'b0),
    .b(sum_21[53]),
    .c(cout_22[52]),
    .cout(cout_22[53]),
    .sum(sum_22[53]));
  AL_FADD comp22_54 (
    .a(1'b0),
    .b(sum_21[54]),
    .c(cout_22[53]),
    .cout(cout_22[54]),
    .sum(sum_22[54]));
  AL_FADD comp22_55 (
    .a(1'b0),
    .b(sum_21[55]),
    .c(cout_22[54]),
    .cout(cout_22[55]),
    .sum(sum_22[55]));
  AL_FADD comp22_56 (
    .a(1'b0),
    .b(sum_21[56]),
    .c(cout_22[55]),
    .cout(cout_22[56]),
    .sum(sum_22[56]));
  AL_FADD comp22_57 (
    .a(1'b0),
    .b(sum_21[57]),
    .c(cout_22[56]),
    .cout(cout_22[57]),
    .sum(sum_22[57]));
  AL_FADD comp22_58 (
    .a(1'b0),
    .b(sum_21[58]),
    .c(cout_22[57]),
    .cout(cout_22[58]),
    .sum(sum_22[58]));
  AL_FADD comp22_59 (
    .a(1'b0),
    .b(sum_21[59]),
    .c(cout_22[58]),
    .cout(cout_22[59]),
    .sum(sum_22[59]));
  AL_FADD comp22_6 (
    .a(i22[6]),
    .b(sum_21[6]),
    .c(cout_22[5]),
    .cout(cout_22[6]),
    .sum(sum_22[6]));
  AL_FADD comp22_60 (
    .a(1'b0),
    .b(sum_21[60]),
    .c(cout_22[59]),
    .cout(cout_22[60]),
    .sum(sum_22[60]));
  AL_FADD comp22_61 (
    .a(1'b0),
    .b(sum_21[61]),
    .c(cout_22[60]),
    .cout(cout_22[61]),
    .sum(sum_22[61]));
  AL_FADD comp22_62 (
    .a(1'b0),
    .b(sum_21[62]),
    .c(cout_22[61]),
    .cout(cout_22[62]),
    .sum(sum_22[62]));
  AL_FADD comp22_63 (
    .a(1'b0),
    .b(sum_21[63]),
    .c(cout_22[62]),
    .cout(cout_22[63]),
    .sum(sum_22[63]));
  AL_FADD comp22_7 (
    .a(i22[7]),
    .b(sum_21[7]),
    .c(cout_22[6]),
    .cout(cout_22[7]),
    .sum(sum_22[7]));
  AL_FADD comp22_8 (
    .a(i22[8]),
    .b(sum_21[8]),
    .c(cout_22[7]),
    .cout(cout_22[8]),
    .sum(sum_22[8]));
  AL_FADD comp22_9 (
    .a(i22[9]),
    .b(sum_21[9]),
    .c(cout_22[8]),
    .cout(cout_22[9]),
    .sum(sum_22[9]));
  AL_FADD comp23_0 (
    .a(i23[0]),
    .b(sum_22[0]),
    .c(1'b0),
    .cout(cout_23[0]),
    .sum(sum_23[0]));
  AL_FADD comp23_1 (
    .a(i23[1]),
    .b(sum_22[1]),
    .c(cout_23[0]),
    .cout(cout_23[1]),
    .sum(sum_23[1]));
  AL_FADD comp23_10 (
    .a(i23[10]),
    .b(sum_22[10]),
    .c(cout_23[9]),
    .cout(cout_23[10]),
    .sum(sum_23[10]));
  AL_FADD comp23_11 (
    .a(i23[11]),
    .b(sum_22[11]),
    .c(cout_23[10]),
    .cout(cout_23[11]),
    .sum(sum_23[11]));
  AL_FADD comp23_12 (
    .a(i23[12]),
    .b(sum_22[12]),
    .c(cout_23[11]),
    .cout(cout_23[12]),
    .sum(sum_23[12]));
  AL_FADD comp23_13 (
    .a(i23[13]),
    .b(sum_22[13]),
    .c(cout_23[12]),
    .cout(cout_23[13]),
    .sum(sum_23[13]));
  AL_FADD comp23_14 (
    .a(i23[14]),
    .b(sum_22[14]),
    .c(cout_23[13]),
    .cout(cout_23[14]),
    .sum(sum_23[14]));
  AL_FADD comp23_15 (
    .a(i23[15]),
    .b(sum_22[15]),
    .c(cout_23[14]),
    .cout(cout_23[15]),
    .sum(sum_23[15]));
  AL_FADD comp23_16 (
    .a(i23[16]),
    .b(sum_22[16]),
    .c(cout_23[15]),
    .cout(cout_23[16]),
    .sum(sum_23[16]));
  AL_FADD comp23_17 (
    .a(i23[17]),
    .b(sum_22[17]),
    .c(cout_23[16]),
    .cout(cout_23[17]),
    .sum(sum_23[17]));
  AL_FADD comp23_18 (
    .a(i23[18]),
    .b(sum_22[18]),
    .c(cout_23[17]),
    .cout(cout_23[18]),
    .sum(sum_23[18]));
  AL_FADD comp23_19 (
    .a(i23[19]),
    .b(sum_22[19]),
    .c(cout_23[18]),
    .cout(cout_23[19]),
    .sum(sum_23[19]));
  AL_FADD comp23_2 (
    .a(i23[2]),
    .b(sum_22[2]),
    .c(cout_23[1]),
    .cout(cout_23[2]),
    .sum(sum_23[2]));
  AL_FADD comp23_20 (
    .a(i23[20]),
    .b(sum_22[20]),
    .c(cout_23[19]),
    .cout(cout_23[20]),
    .sum(sum_23[20]));
  AL_FADD comp23_21 (
    .a(i23[21]),
    .b(sum_22[21]),
    .c(cout_23[20]),
    .cout(cout_23[21]),
    .sum(sum_23[21]));
  AL_FADD comp23_22 (
    .a(i23[22]),
    .b(sum_22[22]),
    .c(cout_23[21]),
    .cout(cout_23[22]),
    .sum(sum_23[22]));
  AL_FADD comp23_23 (
    .a(i23[23]),
    .b(sum_22[23]),
    .c(cout_23[22]),
    .cout(cout_23[23]),
    .sum(sum_23[23]));
  AL_FADD comp23_24 (
    .a(i23[24]),
    .b(sum_22[24]),
    .c(cout_23[23]),
    .cout(cout_23[24]),
    .sum(sum_23[24]));
  AL_FADD comp23_25 (
    .a(i23[25]),
    .b(sum_22[25]),
    .c(cout_23[24]),
    .cout(cout_23[25]),
    .sum(sum_23[25]));
  AL_FADD comp23_26 (
    .a(i23[26]),
    .b(sum_22[26]),
    .c(cout_23[25]),
    .cout(cout_23[26]),
    .sum(sum_23[26]));
  AL_FADD comp23_27 (
    .a(i23[27]),
    .b(sum_22[27]),
    .c(cout_23[26]),
    .cout(cout_23[27]),
    .sum(sum_23[27]));
  AL_FADD comp23_28 (
    .a(i23[28]),
    .b(sum_22[28]),
    .c(cout_23[27]),
    .cout(cout_23[28]),
    .sum(sum_23[28]));
  AL_FADD comp23_29 (
    .a(i23[29]),
    .b(sum_22[29]),
    .c(cout_23[28]),
    .cout(cout_23[29]),
    .sum(sum_23[29]));
  AL_FADD comp23_3 (
    .a(i23[3]),
    .b(sum_22[3]),
    .c(cout_23[2]),
    .cout(cout_23[3]),
    .sum(sum_23[3]));
  AL_FADD comp23_30 (
    .a(i23[30]),
    .b(sum_22[30]),
    .c(cout_23[29]),
    .cout(cout_23[30]),
    .sum(sum_23[30]));
  AL_FADD comp23_31 (
    .a(i23[31]),
    .b(sum_22[31]),
    .c(cout_23[30]),
    .cout(cout_23[31]),
    .sum(sum_23[31]));
  AL_FADD comp23_32 (
    .a(i23[32]),
    .b(sum_22[32]),
    .c(cout_23[31]),
    .cout(cout_23[32]),
    .sum(sum_23[32]));
  AL_FADD comp23_33 (
    .a(i23[33]),
    .b(sum_22[33]),
    .c(cout_23[32]),
    .cout(cout_23[33]),
    .sum(sum_23[33]));
  AL_FADD comp23_34 (
    .a(i23[34]),
    .b(sum_22[34]),
    .c(cout_23[33]),
    .cout(cout_23[34]),
    .sum(sum_23[34]));
  AL_FADD comp23_35 (
    .a(i23[35]),
    .b(sum_22[35]),
    .c(cout_23[34]),
    .cout(cout_23[35]),
    .sum(sum_23[35]));
  AL_FADD comp23_36 (
    .a(i23[36]),
    .b(sum_22[36]),
    .c(cout_23[35]),
    .cout(cout_23[36]),
    .sum(sum_23[36]));
  AL_FADD comp23_37 (
    .a(i23[37]),
    .b(sum_22[37]),
    .c(cout_23[36]),
    .cout(cout_23[37]),
    .sum(sum_23[37]));
  AL_FADD comp23_38 (
    .a(1'b0),
    .b(sum_22[38]),
    .c(cout_23[37]),
    .cout(cout_23[38]),
    .sum(sum_23[38]));
  AL_FADD comp23_39 (
    .a(1'b0),
    .b(sum_22[39]),
    .c(cout_23[38]),
    .cout(cout_23[39]),
    .sum(sum_23[39]));
  AL_FADD comp23_4 (
    .a(i23[4]),
    .b(sum_22[4]),
    .c(cout_23[3]),
    .cout(cout_23[4]),
    .sum(sum_23[4]));
  AL_FADD comp23_40 (
    .a(1'b0),
    .b(sum_22[40]),
    .c(cout_23[39]),
    .cout(cout_23[40]),
    .sum(sum_23[40]));
  AL_FADD comp23_41 (
    .a(1'b0),
    .b(sum_22[41]),
    .c(cout_23[40]),
    .cout(cout_23[41]),
    .sum(sum_23[41]));
  AL_FADD comp23_42 (
    .a(1'b0),
    .b(sum_22[42]),
    .c(cout_23[41]),
    .cout(cout_23[42]),
    .sum(sum_23[42]));
  AL_FADD comp23_43 (
    .a(1'b0),
    .b(sum_22[43]),
    .c(cout_23[42]),
    .cout(cout_23[43]),
    .sum(sum_23[43]));
  AL_FADD comp23_44 (
    .a(1'b0),
    .b(sum_22[44]),
    .c(cout_23[43]),
    .cout(cout_23[44]),
    .sum(sum_23[44]));
  AL_FADD comp23_45 (
    .a(1'b0),
    .b(sum_22[45]),
    .c(cout_23[44]),
    .cout(cout_23[45]),
    .sum(sum_23[45]));
  AL_FADD comp23_46 (
    .a(1'b0),
    .b(sum_22[46]),
    .c(cout_23[45]),
    .cout(cout_23[46]),
    .sum(sum_23[46]));
  AL_FADD comp23_47 (
    .a(1'b0),
    .b(sum_22[47]),
    .c(cout_23[46]),
    .cout(cout_23[47]),
    .sum(sum_23[47]));
  AL_FADD comp23_48 (
    .a(1'b0),
    .b(sum_22[48]),
    .c(cout_23[47]),
    .cout(cout_23[48]),
    .sum(sum_23[48]));
  AL_FADD comp23_49 (
    .a(1'b0),
    .b(sum_22[49]),
    .c(cout_23[48]),
    .cout(cout_23[49]),
    .sum(sum_23[49]));
  AL_FADD comp23_5 (
    .a(i23[5]),
    .b(sum_22[5]),
    .c(cout_23[4]),
    .cout(cout_23[5]),
    .sum(sum_23[5]));
  AL_FADD comp23_50 (
    .a(1'b0),
    .b(sum_22[50]),
    .c(cout_23[49]),
    .cout(cout_23[50]),
    .sum(sum_23[50]));
  AL_FADD comp23_51 (
    .a(1'b0),
    .b(sum_22[51]),
    .c(cout_23[50]),
    .cout(cout_23[51]),
    .sum(sum_23[51]));
  AL_FADD comp23_52 (
    .a(1'b0),
    .b(sum_22[52]),
    .c(cout_23[51]),
    .cout(cout_23[52]),
    .sum(sum_23[52]));
  AL_FADD comp23_53 (
    .a(1'b0),
    .b(sum_22[53]),
    .c(cout_23[52]),
    .cout(cout_23[53]),
    .sum(sum_23[53]));
  AL_FADD comp23_54 (
    .a(1'b0),
    .b(sum_22[54]),
    .c(cout_23[53]),
    .cout(cout_23[54]),
    .sum(sum_23[54]));
  AL_FADD comp23_55 (
    .a(1'b0),
    .b(sum_22[55]),
    .c(cout_23[54]),
    .cout(cout_23[55]),
    .sum(sum_23[55]));
  AL_FADD comp23_56 (
    .a(1'b0),
    .b(sum_22[56]),
    .c(cout_23[55]),
    .cout(cout_23[56]),
    .sum(sum_23[56]));
  AL_FADD comp23_57 (
    .a(1'b0),
    .b(sum_22[57]),
    .c(cout_23[56]),
    .cout(cout_23[57]),
    .sum(sum_23[57]));
  AL_FADD comp23_58 (
    .a(1'b0),
    .b(sum_22[58]),
    .c(cout_23[57]),
    .cout(cout_23[58]),
    .sum(sum_23[58]));
  AL_FADD comp23_59 (
    .a(1'b0),
    .b(sum_22[59]),
    .c(cout_23[58]),
    .cout(cout_23[59]),
    .sum(sum_23[59]));
  AL_FADD comp23_6 (
    .a(i23[6]),
    .b(sum_22[6]),
    .c(cout_23[5]),
    .cout(cout_23[6]),
    .sum(sum_23[6]));
  AL_FADD comp23_60 (
    .a(1'b0),
    .b(sum_22[60]),
    .c(cout_23[59]),
    .cout(cout_23[60]),
    .sum(sum_23[60]));
  AL_FADD comp23_61 (
    .a(1'b0),
    .b(sum_22[61]),
    .c(cout_23[60]),
    .cout(cout_23[61]),
    .sum(sum_23[61]));
  AL_FADD comp23_62 (
    .a(1'b0),
    .b(sum_22[62]),
    .c(cout_23[61]),
    .cout(cout_23[62]),
    .sum(sum_23[62]));
  AL_FADD comp23_63 (
    .a(1'b0),
    .b(sum_22[63]),
    .c(cout_23[62]),
    .cout(cout_23[63]),
    .sum(sum_23[63]));
  AL_FADD comp23_7 (
    .a(i23[7]),
    .b(sum_22[7]),
    .c(cout_23[6]),
    .cout(cout_23[7]),
    .sum(sum_23[7]));
  AL_FADD comp23_8 (
    .a(i23[8]),
    .b(sum_22[8]),
    .c(cout_23[7]),
    .cout(cout_23[8]),
    .sum(sum_23[8]));
  AL_FADD comp23_9 (
    .a(i23[9]),
    .b(sum_22[9]),
    .c(cout_23[8]),
    .cout(cout_23[9]),
    .sum(sum_23[9]));
  AL_FADD comp24_0 (
    .a(i24[0]),
    .b(sum_23[0]),
    .c(1'b0),
    .cout(cout_24[0]),
    .sum(sum_24[0]));
  AL_FADD comp24_1 (
    .a(i24[1]),
    .b(sum_23[1]),
    .c(cout_24[0]),
    .cout(cout_24[1]),
    .sum(sum_24[1]));
  AL_FADD comp24_10 (
    .a(i24[10]),
    .b(sum_23[10]),
    .c(cout_24[9]),
    .cout(cout_24[10]),
    .sum(sum_24[10]));
  AL_FADD comp24_11 (
    .a(i24[11]),
    .b(sum_23[11]),
    .c(cout_24[10]),
    .cout(cout_24[11]),
    .sum(sum_24[11]));
  AL_FADD comp24_12 (
    .a(i24[12]),
    .b(sum_23[12]),
    .c(cout_24[11]),
    .cout(cout_24[12]),
    .sum(sum_24[12]));
  AL_FADD comp24_13 (
    .a(i24[13]),
    .b(sum_23[13]),
    .c(cout_24[12]),
    .cout(cout_24[13]),
    .sum(sum_24[13]));
  AL_FADD comp24_14 (
    .a(i24[14]),
    .b(sum_23[14]),
    .c(cout_24[13]),
    .cout(cout_24[14]),
    .sum(sum_24[14]));
  AL_FADD comp24_15 (
    .a(i24[15]),
    .b(sum_23[15]),
    .c(cout_24[14]),
    .cout(cout_24[15]),
    .sum(sum_24[15]));
  AL_FADD comp24_16 (
    .a(i24[16]),
    .b(sum_23[16]),
    .c(cout_24[15]),
    .cout(cout_24[16]),
    .sum(sum_24[16]));
  AL_FADD comp24_17 (
    .a(i24[17]),
    .b(sum_23[17]),
    .c(cout_24[16]),
    .cout(cout_24[17]),
    .sum(sum_24[17]));
  AL_FADD comp24_18 (
    .a(i24[18]),
    .b(sum_23[18]),
    .c(cout_24[17]),
    .cout(cout_24[18]),
    .sum(sum_24[18]));
  AL_FADD comp24_19 (
    .a(i24[19]),
    .b(sum_23[19]),
    .c(cout_24[18]),
    .cout(cout_24[19]),
    .sum(sum_24[19]));
  AL_FADD comp24_2 (
    .a(i24[2]),
    .b(sum_23[2]),
    .c(cout_24[1]),
    .cout(cout_24[2]),
    .sum(sum_24[2]));
  AL_FADD comp24_20 (
    .a(i24[20]),
    .b(sum_23[20]),
    .c(cout_24[19]),
    .cout(cout_24[20]),
    .sum(sum_24[20]));
  AL_FADD comp24_21 (
    .a(i24[21]),
    .b(sum_23[21]),
    .c(cout_24[20]),
    .cout(cout_24[21]),
    .sum(sum_24[21]));
  AL_FADD comp24_22 (
    .a(i24[22]),
    .b(sum_23[22]),
    .c(cout_24[21]),
    .cout(cout_24[22]),
    .sum(sum_24[22]));
  AL_FADD comp24_23 (
    .a(i24[23]),
    .b(sum_23[23]),
    .c(cout_24[22]),
    .cout(cout_24[23]),
    .sum(sum_24[23]));
  AL_FADD comp24_24 (
    .a(i24[24]),
    .b(sum_23[24]),
    .c(cout_24[23]),
    .cout(cout_24[24]),
    .sum(sum_24[24]));
  AL_FADD comp24_25 (
    .a(i24[25]),
    .b(sum_23[25]),
    .c(cout_24[24]),
    .cout(cout_24[25]),
    .sum(sum_24[25]));
  AL_FADD comp24_26 (
    .a(i24[26]),
    .b(sum_23[26]),
    .c(cout_24[25]),
    .cout(cout_24[26]),
    .sum(sum_24[26]));
  AL_FADD comp24_27 (
    .a(i24[27]),
    .b(sum_23[27]),
    .c(cout_24[26]),
    .cout(cout_24[27]),
    .sum(sum_24[27]));
  AL_FADD comp24_28 (
    .a(i24[28]),
    .b(sum_23[28]),
    .c(cout_24[27]),
    .cout(cout_24[28]),
    .sum(sum_24[28]));
  AL_FADD comp24_29 (
    .a(i24[29]),
    .b(sum_23[29]),
    .c(cout_24[28]),
    .cout(cout_24[29]),
    .sum(sum_24[29]));
  AL_FADD comp24_3 (
    .a(i24[3]),
    .b(sum_23[3]),
    .c(cout_24[2]),
    .cout(cout_24[3]),
    .sum(sum_24[3]));
  AL_FADD comp24_30 (
    .a(i24[30]),
    .b(sum_23[30]),
    .c(cout_24[29]),
    .cout(cout_24[30]),
    .sum(sum_24[30]));
  AL_FADD comp24_31 (
    .a(i24[31]),
    .b(sum_23[31]),
    .c(cout_24[30]),
    .cout(cout_24[31]),
    .sum(sum_24[31]));
  AL_FADD comp24_32 (
    .a(i24[32]),
    .b(sum_23[32]),
    .c(cout_24[31]),
    .cout(cout_24[32]),
    .sum(sum_24[32]));
  AL_FADD comp24_33 (
    .a(i24[33]),
    .b(sum_23[33]),
    .c(cout_24[32]),
    .cout(cout_24[33]),
    .sum(sum_24[33]));
  AL_FADD comp24_34 (
    .a(i24[34]),
    .b(sum_23[34]),
    .c(cout_24[33]),
    .cout(cout_24[34]),
    .sum(sum_24[34]));
  AL_FADD comp24_35 (
    .a(i24[35]),
    .b(sum_23[35]),
    .c(cout_24[34]),
    .cout(cout_24[35]),
    .sum(sum_24[35]));
  AL_FADD comp24_36 (
    .a(i24[36]),
    .b(sum_23[36]),
    .c(cout_24[35]),
    .cout(cout_24[36]),
    .sum(sum_24[36]));
  AL_FADD comp24_37 (
    .a(1'b0),
    .b(sum_23[37]),
    .c(cout_24[36]),
    .cout(cout_24[37]),
    .sum(sum_24[37]));
  AL_FADD comp24_38 (
    .a(1'b0),
    .b(sum_23[38]),
    .c(cout_24[37]),
    .cout(cout_24[38]),
    .sum(sum_24[38]));
  AL_FADD comp24_39 (
    .a(1'b0),
    .b(sum_23[39]),
    .c(cout_24[38]),
    .cout(cout_24[39]),
    .sum(sum_24[39]));
  AL_FADD comp24_4 (
    .a(i24[4]),
    .b(sum_23[4]),
    .c(cout_24[3]),
    .cout(cout_24[4]),
    .sum(sum_24[4]));
  AL_FADD comp24_40 (
    .a(1'b0),
    .b(sum_23[40]),
    .c(cout_24[39]),
    .cout(cout_24[40]),
    .sum(sum_24[40]));
  AL_FADD comp24_41 (
    .a(1'b0),
    .b(sum_23[41]),
    .c(cout_24[40]),
    .cout(cout_24[41]),
    .sum(sum_24[41]));
  AL_FADD comp24_42 (
    .a(1'b0),
    .b(sum_23[42]),
    .c(cout_24[41]),
    .cout(cout_24[42]),
    .sum(sum_24[42]));
  AL_FADD comp24_43 (
    .a(1'b0),
    .b(sum_23[43]),
    .c(cout_24[42]),
    .cout(cout_24[43]),
    .sum(sum_24[43]));
  AL_FADD comp24_44 (
    .a(1'b0),
    .b(sum_23[44]),
    .c(cout_24[43]),
    .cout(cout_24[44]),
    .sum(sum_24[44]));
  AL_FADD comp24_45 (
    .a(1'b0),
    .b(sum_23[45]),
    .c(cout_24[44]),
    .cout(cout_24[45]),
    .sum(sum_24[45]));
  AL_FADD comp24_46 (
    .a(1'b0),
    .b(sum_23[46]),
    .c(cout_24[45]),
    .cout(cout_24[46]),
    .sum(sum_24[46]));
  AL_FADD comp24_47 (
    .a(1'b0),
    .b(sum_23[47]),
    .c(cout_24[46]),
    .cout(cout_24[47]),
    .sum(sum_24[47]));
  AL_FADD comp24_48 (
    .a(1'b0),
    .b(sum_23[48]),
    .c(cout_24[47]),
    .cout(cout_24[48]),
    .sum(sum_24[48]));
  AL_FADD comp24_49 (
    .a(1'b0),
    .b(sum_23[49]),
    .c(cout_24[48]),
    .cout(cout_24[49]),
    .sum(sum_24[49]));
  AL_FADD comp24_5 (
    .a(i24[5]),
    .b(sum_23[5]),
    .c(cout_24[4]),
    .cout(cout_24[5]),
    .sum(sum_24[5]));
  AL_FADD comp24_50 (
    .a(1'b0),
    .b(sum_23[50]),
    .c(cout_24[49]),
    .cout(cout_24[50]),
    .sum(sum_24[50]));
  AL_FADD comp24_51 (
    .a(1'b0),
    .b(sum_23[51]),
    .c(cout_24[50]),
    .cout(cout_24[51]),
    .sum(sum_24[51]));
  AL_FADD comp24_52 (
    .a(1'b0),
    .b(sum_23[52]),
    .c(cout_24[51]),
    .cout(cout_24[52]),
    .sum(sum_24[52]));
  AL_FADD comp24_53 (
    .a(1'b0),
    .b(sum_23[53]),
    .c(cout_24[52]),
    .cout(cout_24[53]),
    .sum(sum_24[53]));
  AL_FADD comp24_54 (
    .a(1'b0),
    .b(sum_23[54]),
    .c(cout_24[53]),
    .cout(cout_24[54]),
    .sum(sum_24[54]));
  AL_FADD comp24_55 (
    .a(1'b0),
    .b(sum_23[55]),
    .c(cout_24[54]),
    .cout(cout_24[55]),
    .sum(sum_24[55]));
  AL_FADD comp24_56 (
    .a(1'b0),
    .b(sum_23[56]),
    .c(cout_24[55]),
    .cout(cout_24[56]),
    .sum(sum_24[56]));
  AL_FADD comp24_57 (
    .a(1'b0),
    .b(sum_23[57]),
    .c(cout_24[56]),
    .cout(cout_24[57]),
    .sum(sum_24[57]));
  AL_FADD comp24_58 (
    .a(1'b0),
    .b(sum_23[58]),
    .c(cout_24[57]),
    .cout(cout_24[58]),
    .sum(sum_24[58]));
  AL_FADD comp24_59 (
    .a(1'b0),
    .b(sum_23[59]),
    .c(cout_24[58]),
    .cout(cout_24[59]),
    .sum(sum_24[59]));
  AL_FADD comp24_6 (
    .a(i24[6]),
    .b(sum_23[6]),
    .c(cout_24[5]),
    .cout(cout_24[6]),
    .sum(sum_24[6]));
  AL_FADD comp24_60 (
    .a(1'b0),
    .b(sum_23[60]),
    .c(cout_24[59]),
    .cout(cout_24[60]),
    .sum(sum_24[60]));
  AL_FADD comp24_61 (
    .a(1'b0),
    .b(sum_23[61]),
    .c(cout_24[60]),
    .cout(cout_24[61]),
    .sum(sum_24[61]));
  AL_FADD comp24_62 (
    .a(1'b0),
    .b(sum_23[62]),
    .c(cout_24[61]),
    .cout(cout_24[62]),
    .sum(sum_24[62]));
  AL_FADD comp24_63 (
    .a(1'b0),
    .b(sum_23[63]),
    .c(cout_24[62]),
    .cout(cout_24[63]),
    .sum(sum_24[63]));
  AL_FADD comp24_7 (
    .a(i24[7]),
    .b(sum_23[7]),
    .c(cout_24[6]),
    .cout(cout_24[7]),
    .sum(sum_24[7]));
  AL_FADD comp24_8 (
    .a(i24[8]),
    .b(sum_23[8]),
    .c(cout_24[7]),
    .cout(cout_24[8]),
    .sum(sum_24[8]));
  AL_FADD comp24_9 (
    .a(i24[9]),
    .b(sum_23[9]),
    .c(cout_24[8]),
    .cout(cout_24[9]),
    .sum(sum_24[9]));
  AL_FADD comp25_0 (
    .a(i25[0]),
    .b(sum_24[0]),
    .c(1'b0),
    .cout(cout_25[0]),
    .sum(sum_25[0]));
  AL_FADD comp25_1 (
    .a(i25[1]),
    .b(sum_24[1]),
    .c(cout_25[0]),
    .cout(cout_25[1]),
    .sum(sum_25[1]));
  AL_FADD comp25_10 (
    .a(i25[10]),
    .b(sum_24[10]),
    .c(cout_25[9]),
    .cout(cout_25[10]),
    .sum(sum_25[10]));
  AL_FADD comp25_11 (
    .a(i25[11]),
    .b(sum_24[11]),
    .c(cout_25[10]),
    .cout(cout_25[11]),
    .sum(sum_25[11]));
  AL_FADD comp25_12 (
    .a(i25[12]),
    .b(sum_24[12]),
    .c(cout_25[11]),
    .cout(cout_25[12]),
    .sum(sum_25[12]));
  AL_FADD comp25_13 (
    .a(i25[13]),
    .b(sum_24[13]),
    .c(cout_25[12]),
    .cout(cout_25[13]),
    .sum(sum_25[13]));
  AL_FADD comp25_14 (
    .a(i25[14]),
    .b(sum_24[14]),
    .c(cout_25[13]),
    .cout(cout_25[14]),
    .sum(sum_25[14]));
  AL_FADD comp25_15 (
    .a(i25[15]),
    .b(sum_24[15]),
    .c(cout_25[14]),
    .cout(cout_25[15]),
    .sum(sum_25[15]));
  AL_FADD comp25_16 (
    .a(i25[16]),
    .b(sum_24[16]),
    .c(cout_25[15]),
    .cout(cout_25[16]),
    .sum(sum_25[16]));
  AL_FADD comp25_17 (
    .a(i25[17]),
    .b(sum_24[17]),
    .c(cout_25[16]),
    .cout(cout_25[17]),
    .sum(sum_25[17]));
  AL_FADD comp25_18 (
    .a(i25[18]),
    .b(sum_24[18]),
    .c(cout_25[17]),
    .cout(cout_25[18]),
    .sum(sum_25[18]));
  AL_FADD comp25_19 (
    .a(i25[19]),
    .b(sum_24[19]),
    .c(cout_25[18]),
    .cout(cout_25[19]),
    .sum(sum_25[19]));
  AL_FADD comp25_2 (
    .a(i25[2]),
    .b(sum_24[2]),
    .c(cout_25[1]),
    .cout(cout_25[2]),
    .sum(sum_25[2]));
  AL_FADD comp25_20 (
    .a(i25[20]),
    .b(sum_24[20]),
    .c(cout_25[19]),
    .cout(cout_25[20]),
    .sum(sum_25[20]));
  AL_FADD comp25_21 (
    .a(i25[21]),
    .b(sum_24[21]),
    .c(cout_25[20]),
    .cout(cout_25[21]),
    .sum(sum_25[21]));
  AL_FADD comp25_22 (
    .a(i25[22]),
    .b(sum_24[22]),
    .c(cout_25[21]),
    .cout(cout_25[22]),
    .sum(sum_25[22]));
  AL_FADD comp25_23 (
    .a(i25[23]),
    .b(sum_24[23]),
    .c(cout_25[22]),
    .cout(cout_25[23]),
    .sum(sum_25[23]));
  AL_FADD comp25_24 (
    .a(i25[24]),
    .b(sum_24[24]),
    .c(cout_25[23]),
    .cout(cout_25[24]),
    .sum(sum_25[24]));
  AL_FADD comp25_25 (
    .a(i25[25]),
    .b(sum_24[25]),
    .c(cout_25[24]),
    .cout(cout_25[25]),
    .sum(sum_25[25]));
  AL_FADD comp25_26 (
    .a(i25[26]),
    .b(sum_24[26]),
    .c(cout_25[25]),
    .cout(cout_25[26]),
    .sum(sum_25[26]));
  AL_FADD comp25_27 (
    .a(i25[27]),
    .b(sum_24[27]),
    .c(cout_25[26]),
    .cout(cout_25[27]),
    .sum(sum_25[27]));
  AL_FADD comp25_28 (
    .a(i25[28]),
    .b(sum_24[28]),
    .c(cout_25[27]),
    .cout(cout_25[28]),
    .sum(sum_25[28]));
  AL_FADD comp25_29 (
    .a(i25[29]),
    .b(sum_24[29]),
    .c(cout_25[28]),
    .cout(cout_25[29]),
    .sum(sum_25[29]));
  AL_FADD comp25_3 (
    .a(i25[3]),
    .b(sum_24[3]),
    .c(cout_25[2]),
    .cout(cout_25[3]),
    .sum(sum_25[3]));
  AL_FADD comp25_30 (
    .a(i25[30]),
    .b(sum_24[30]),
    .c(cout_25[29]),
    .cout(cout_25[30]),
    .sum(sum_25[30]));
  AL_FADD comp25_31 (
    .a(i25[31]),
    .b(sum_24[31]),
    .c(cout_25[30]),
    .cout(cout_25[31]),
    .sum(sum_25[31]));
  AL_FADD comp25_32 (
    .a(i25[32]),
    .b(sum_24[32]),
    .c(cout_25[31]),
    .cout(cout_25[32]),
    .sum(sum_25[32]));
  AL_FADD comp25_33 (
    .a(i25[33]),
    .b(sum_24[33]),
    .c(cout_25[32]),
    .cout(cout_25[33]),
    .sum(sum_25[33]));
  AL_FADD comp25_34 (
    .a(i25[34]),
    .b(sum_24[34]),
    .c(cout_25[33]),
    .cout(cout_25[34]),
    .sum(sum_25[34]));
  AL_FADD comp25_35 (
    .a(i25[35]),
    .b(sum_24[35]),
    .c(cout_25[34]),
    .cout(cout_25[35]),
    .sum(sum_25[35]));
  AL_FADD comp25_36 (
    .a(1'b0),
    .b(sum_24[36]),
    .c(cout_25[35]),
    .cout(cout_25[36]),
    .sum(sum_25[36]));
  AL_FADD comp25_37 (
    .a(1'b0),
    .b(sum_24[37]),
    .c(cout_25[36]),
    .cout(cout_25[37]),
    .sum(sum_25[37]));
  AL_FADD comp25_38 (
    .a(1'b0),
    .b(sum_24[38]),
    .c(cout_25[37]),
    .cout(cout_25[38]),
    .sum(sum_25[38]));
  AL_FADD comp25_39 (
    .a(1'b0),
    .b(sum_24[39]),
    .c(cout_25[38]),
    .cout(cout_25[39]),
    .sum(sum_25[39]));
  AL_FADD comp25_4 (
    .a(i25[4]),
    .b(sum_24[4]),
    .c(cout_25[3]),
    .cout(cout_25[4]),
    .sum(sum_25[4]));
  AL_FADD comp25_40 (
    .a(1'b0),
    .b(sum_24[40]),
    .c(cout_25[39]),
    .cout(cout_25[40]),
    .sum(sum_25[40]));
  AL_FADD comp25_41 (
    .a(1'b0),
    .b(sum_24[41]),
    .c(cout_25[40]),
    .cout(cout_25[41]),
    .sum(sum_25[41]));
  AL_FADD comp25_42 (
    .a(1'b0),
    .b(sum_24[42]),
    .c(cout_25[41]),
    .cout(cout_25[42]),
    .sum(sum_25[42]));
  AL_FADD comp25_43 (
    .a(1'b0),
    .b(sum_24[43]),
    .c(cout_25[42]),
    .cout(cout_25[43]),
    .sum(sum_25[43]));
  AL_FADD comp25_44 (
    .a(1'b0),
    .b(sum_24[44]),
    .c(cout_25[43]),
    .cout(cout_25[44]),
    .sum(sum_25[44]));
  AL_FADD comp25_45 (
    .a(1'b0),
    .b(sum_24[45]),
    .c(cout_25[44]),
    .cout(cout_25[45]),
    .sum(sum_25[45]));
  AL_FADD comp25_46 (
    .a(1'b0),
    .b(sum_24[46]),
    .c(cout_25[45]),
    .cout(cout_25[46]),
    .sum(sum_25[46]));
  AL_FADD comp25_47 (
    .a(1'b0),
    .b(sum_24[47]),
    .c(cout_25[46]),
    .cout(cout_25[47]),
    .sum(sum_25[47]));
  AL_FADD comp25_48 (
    .a(1'b0),
    .b(sum_24[48]),
    .c(cout_25[47]),
    .cout(cout_25[48]),
    .sum(sum_25[48]));
  AL_FADD comp25_49 (
    .a(1'b0),
    .b(sum_24[49]),
    .c(cout_25[48]),
    .cout(cout_25[49]),
    .sum(sum_25[49]));
  AL_FADD comp25_5 (
    .a(i25[5]),
    .b(sum_24[5]),
    .c(cout_25[4]),
    .cout(cout_25[5]),
    .sum(sum_25[5]));
  AL_FADD comp25_50 (
    .a(1'b0),
    .b(sum_24[50]),
    .c(cout_25[49]),
    .cout(cout_25[50]),
    .sum(sum_25[50]));
  AL_FADD comp25_51 (
    .a(1'b0),
    .b(sum_24[51]),
    .c(cout_25[50]),
    .cout(cout_25[51]),
    .sum(sum_25[51]));
  AL_FADD comp25_52 (
    .a(1'b0),
    .b(sum_24[52]),
    .c(cout_25[51]),
    .cout(cout_25[52]),
    .sum(sum_25[52]));
  AL_FADD comp25_53 (
    .a(1'b0),
    .b(sum_24[53]),
    .c(cout_25[52]),
    .cout(cout_25[53]),
    .sum(sum_25[53]));
  AL_FADD comp25_54 (
    .a(1'b0),
    .b(sum_24[54]),
    .c(cout_25[53]),
    .cout(cout_25[54]),
    .sum(sum_25[54]));
  AL_FADD comp25_55 (
    .a(1'b0),
    .b(sum_24[55]),
    .c(cout_25[54]),
    .cout(cout_25[55]),
    .sum(sum_25[55]));
  AL_FADD comp25_56 (
    .a(1'b0),
    .b(sum_24[56]),
    .c(cout_25[55]),
    .cout(cout_25[56]),
    .sum(sum_25[56]));
  AL_FADD comp25_57 (
    .a(1'b0),
    .b(sum_24[57]),
    .c(cout_25[56]),
    .cout(cout_25[57]),
    .sum(sum_25[57]));
  AL_FADD comp25_58 (
    .a(1'b0),
    .b(sum_24[58]),
    .c(cout_25[57]),
    .cout(cout_25[58]),
    .sum(sum_25[58]));
  AL_FADD comp25_59 (
    .a(1'b0),
    .b(sum_24[59]),
    .c(cout_25[58]),
    .cout(cout_25[59]),
    .sum(sum_25[59]));
  AL_FADD comp25_6 (
    .a(i25[6]),
    .b(sum_24[6]),
    .c(cout_25[5]),
    .cout(cout_25[6]),
    .sum(sum_25[6]));
  AL_FADD comp25_60 (
    .a(1'b0),
    .b(sum_24[60]),
    .c(cout_25[59]),
    .cout(cout_25[60]),
    .sum(sum_25[60]));
  AL_FADD comp25_61 (
    .a(1'b0),
    .b(sum_24[61]),
    .c(cout_25[60]),
    .cout(cout_25[61]),
    .sum(sum_25[61]));
  AL_FADD comp25_62 (
    .a(1'b0),
    .b(sum_24[62]),
    .c(cout_25[61]),
    .cout(cout_25[62]),
    .sum(sum_25[62]));
  AL_FADD comp25_63 (
    .a(1'b0),
    .b(sum_24[63]),
    .c(cout_25[62]),
    .cout(cout_25[63]),
    .sum(sum_25[63]));
  AL_FADD comp25_7 (
    .a(i25[7]),
    .b(sum_24[7]),
    .c(cout_25[6]),
    .cout(cout_25[7]),
    .sum(sum_25[7]));
  AL_FADD comp25_8 (
    .a(i25[8]),
    .b(sum_24[8]),
    .c(cout_25[7]),
    .cout(cout_25[8]),
    .sum(sum_25[8]));
  AL_FADD comp25_9 (
    .a(i25[9]),
    .b(sum_24[9]),
    .c(cout_25[8]),
    .cout(cout_25[9]),
    .sum(sum_25[9]));
  AL_FADD comp26_0 (
    .a(i26[0]),
    .b(sum_25[0]),
    .c(1'b0),
    .cout(cout_26[0]),
    .sum(sum_26[0]));
  AL_FADD comp26_1 (
    .a(i26[1]),
    .b(sum_25[1]),
    .c(cout_26[0]),
    .cout(cout_26[1]),
    .sum(sum_26[1]));
  AL_FADD comp26_10 (
    .a(i26[10]),
    .b(sum_25[10]),
    .c(cout_26[9]),
    .cout(cout_26[10]),
    .sum(sum_26[10]));
  AL_FADD comp26_11 (
    .a(i26[11]),
    .b(sum_25[11]),
    .c(cout_26[10]),
    .cout(cout_26[11]),
    .sum(sum_26[11]));
  AL_FADD comp26_12 (
    .a(i26[12]),
    .b(sum_25[12]),
    .c(cout_26[11]),
    .cout(cout_26[12]),
    .sum(sum_26[12]));
  AL_FADD comp26_13 (
    .a(i26[13]),
    .b(sum_25[13]),
    .c(cout_26[12]),
    .cout(cout_26[13]),
    .sum(sum_26[13]));
  AL_FADD comp26_14 (
    .a(i26[14]),
    .b(sum_25[14]),
    .c(cout_26[13]),
    .cout(cout_26[14]),
    .sum(sum_26[14]));
  AL_FADD comp26_15 (
    .a(i26[15]),
    .b(sum_25[15]),
    .c(cout_26[14]),
    .cout(cout_26[15]),
    .sum(sum_26[15]));
  AL_FADD comp26_16 (
    .a(i26[16]),
    .b(sum_25[16]),
    .c(cout_26[15]),
    .cout(cout_26[16]),
    .sum(sum_26[16]));
  AL_FADD comp26_17 (
    .a(i26[17]),
    .b(sum_25[17]),
    .c(cout_26[16]),
    .cout(cout_26[17]),
    .sum(sum_26[17]));
  AL_FADD comp26_18 (
    .a(i26[18]),
    .b(sum_25[18]),
    .c(cout_26[17]),
    .cout(cout_26[18]),
    .sum(sum_26[18]));
  AL_FADD comp26_19 (
    .a(i26[19]),
    .b(sum_25[19]),
    .c(cout_26[18]),
    .cout(cout_26[19]),
    .sum(sum_26[19]));
  AL_FADD comp26_2 (
    .a(i26[2]),
    .b(sum_25[2]),
    .c(cout_26[1]),
    .cout(cout_26[2]),
    .sum(sum_26[2]));
  AL_FADD comp26_20 (
    .a(i26[20]),
    .b(sum_25[20]),
    .c(cout_26[19]),
    .cout(cout_26[20]),
    .sum(sum_26[20]));
  AL_FADD comp26_21 (
    .a(i26[21]),
    .b(sum_25[21]),
    .c(cout_26[20]),
    .cout(cout_26[21]),
    .sum(sum_26[21]));
  AL_FADD comp26_22 (
    .a(i26[22]),
    .b(sum_25[22]),
    .c(cout_26[21]),
    .cout(cout_26[22]),
    .sum(sum_26[22]));
  AL_FADD comp26_23 (
    .a(i26[23]),
    .b(sum_25[23]),
    .c(cout_26[22]),
    .cout(cout_26[23]),
    .sum(sum_26[23]));
  AL_FADD comp26_24 (
    .a(i26[24]),
    .b(sum_25[24]),
    .c(cout_26[23]),
    .cout(cout_26[24]),
    .sum(sum_26[24]));
  AL_FADD comp26_25 (
    .a(i26[25]),
    .b(sum_25[25]),
    .c(cout_26[24]),
    .cout(cout_26[25]),
    .sum(sum_26[25]));
  AL_FADD comp26_26 (
    .a(i26[26]),
    .b(sum_25[26]),
    .c(cout_26[25]),
    .cout(cout_26[26]),
    .sum(sum_26[26]));
  AL_FADD comp26_27 (
    .a(i26[27]),
    .b(sum_25[27]),
    .c(cout_26[26]),
    .cout(cout_26[27]),
    .sum(sum_26[27]));
  AL_FADD comp26_28 (
    .a(i26[28]),
    .b(sum_25[28]),
    .c(cout_26[27]),
    .cout(cout_26[28]),
    .sum(sum_26[28]));
  AL_FADD comp26_29 (
    .a(i26[29]),
    .b(sum_25[29]),
    .c(cout_26[28]),
    .cout(cout_26[29]),
    .sum(sum_26[29]));
  AL_FADD comp26_3 (
    .a(i26[3]),
    .b(sum_25[3]),
    .c(cout_26[2]),
    .cout(cout_26[3]),
    .sum(sum_26[3]));
  AL_FADD comp26_30 (
    .a(i26[30]),
    .b(sum_25[30]),
    .c(cout_26[29]),
    .cout(cout_26[30]),
    .sum(sum_26[30]));
  AL_FADD comp26_31 (
    .a(i26[31]),
    .b(sum_25[31]),
    .c(cout_26[30]),
    .cout(cout_26[31]),
    .sum(sum_26[31]));
  AL_FADD comp26_32 (
    .a(i26[32]),
    .b(sum_25[32]),
    .c(cout_26[31]),
    .cout(cout_26[32]),
    .sum(sum_26[32]));
  AL_FADD comp26_33 (
    .a(i26[33]),
    .b(sum_25[33]),
    .c(cout_26[32]),
    .cout(cout_26[33]),
    .sum(sum_26[33]));
  AL_FADD comp26_34 (
    .a(i26[34]),
    .b(sum_25[34]),
    .c(cout_26[33]),
    .cout(cout_26[34]),
    .sum(sum_26[34]));
  AL_FADD comp26_35 (
    .a(1'b0),
    .b(sum_25[35]),
    .c(cout_26[34]),
    .cout(cout_26[35]),
    .sum(sum_26[35]));
  AL_FADD comp26_36 (
    .a(1'b0),
    .b(sum_25[36]),
    .c(cout_26[35]),
    .cout(cout_26[36]),
    .sum(sum_26[36]));
  AL_FADD comp26_37 (
    .a(1'b0),
    .b(sum_25[37]),
    .c(cout_26[36]),
    .cout(cout_26[37]),
    .sum(sum_26[37]));
  AL_FADD comp26_38 (
    .a(1'b0),
    .b(sum_25[38]),
    .c(cout_26[37]),
    .cout(cout_26[38]),
    .sum(sum_26[38]));
  AL_FADD comp26_39 (
    .a(1'b0),
    .b(sum_25[39]),
    .c(cout_26[38]),
    .cout(cout_26[39]),
    .sum(sum_26[39]));
  AL_FADD comp26_4 (
    .a(i26[4]),
    .b(sum_25[4]),
    .c(cout_26[3]),
    .cout(cout_26[4]),
    .sum(sum_26[4]));
  AL_FADD comp26_40 (
    .a(1'b0),
    .b(sum_25[40]),
    .c(cout_26[39]),
    .cout(cout_26[40]),
    .sum(sum_26[40]));
  AL_FADD comp26_41 (
    .a(1'b0),
    .b(sum_25[41]),
    .c(cout_26[40]),
    .cout(cout_26[41]),
    .sum(sum_26[41]));
  AL_FADD comp26_42 (
    .a(1'b0),
    .b(sum_25[42]),
    .c(cout_26[41]),
    .cout(cout_26[42]),
    .sum(sum_26[42]));
  AL_FADD comp26_43 (
    .a(1'b0),
    .b(sum_25[43]),
    .c(cout_26[42]),
    .cout(cout_26[43]),
    .sum(sum_26[43]));
  AL_FADD comp26_44 (
    .a(1'b0),
    .b(sum_25[44]),
    .c(cout_26[43]),
    .cout(cout_26[44]),
    .sum(sum_26[44]));
  AL_FADD comp26_45 (
    .a(1'b0),
    .b(sum_25[45]),
    .c(cout_26[44]),
    .cout(cout_26[45]),
    .sum(sum_26[45]));
  AL_FADD comp26_46 (
    .a(1'b0),
    .b(sum_25[46]),
    .c(cout_26[45]),
    .cout(cout_26[46]),
    .sum(sum_26[46]));
  AL_FADD comp26_47 (
    .a(1'b0),
    .b(sum_25[47]),
    .c(cout_26[46]),
    .cout(cout_26[47]),
    .sum(sum_26[47]));
  AL_FADD comp26_48 (
    .a(1'b0),
    .b(sum_25[48]),
    .c(cout_26[47]),
    .cout(cout_26[48]),
    .sum(sum_26[48]));
  AL_FADD comp26_49 (
    .a(1'b0),
    .b(sum_25[49]),
    .c(cout_26[48]),
    .cout(cout_26[49]),
    .sum(sum_26[49]));
  AL_FADD comp26_5 (
    .a(i26[5]),
    .b(sum_25[5]),
    .c(cout_26[4]),
    .cout(cout_26[5]),
    .sum(sum_26[5]));
  AL_FADD comp26_50 (
    .a(1'b0),
    .b(sum_25[50]),
    .c(cout_26[49]),
    .cout(cout_26[50]),
    .sum(sum_26[50]));
  AL_FADD comp26_51 (
    .a(1'b0),
    .b(sum_25[51]),
    .c(cout_26[50]),
    .cout(cout_26[51]),
    .sum(sum_26[51]));
  AL_FADD comp26_52 (
    .a(1'b0),
    .b(sum_25[52]),
    .c(cout_26[51]),
    .cout(cout_26[52]),
    .sum(sum_26[52]));
  AL_FADD comp26_53 (
    .a(1'b0),
    .b(sum_25[53]),
    .c(cout_26[52]),
    .cout(cout_26[53]),
    .sum(sum_26[53]));
  AL_FADD comp26_54 (
    .a(1'b0),
    .b(sum_25[54]),
    .c(cout_26[53]),
    .cout(cout_26[54]),
    .sum(sum_26[54]));
  AL_FADD comp26_55 (
    .a(1'b0),
    .b(sum_25[55]),
    .c(cout_26[54]),
    .cout(cout_26[55]),
    .sum(sum_26[55]));
  AL_FADD comp26_56 (
    .a(1'b0),
    .b(sum_25[56]),
    .c(cout_26[55]),
    .cout(cout_26[56]),
    .sum(sum_26[56]));
  AL_FADD comp26_57 (
    .a(1'b0),
    .b(sum_25[57]),
    .c(cout_26[56]),
    .cout(cout_26[57]),
    .sum(sum_26[57]));
  AL_FADD comp26_58 (
    .a(1'b0),
    .b(sum_25[58]),
    .c(cout_26[57]),
    .cout(cout_26[58]),
    .sum(sum_26[58]));
  AL_FADD comp26_59 (
    .a(1'b0),
    .b(sum_25[59]),
    .c(cout_26[58]),
    .cout(cout_26[59]),
    .sum(sum_26[59]));
  AL_FADD comp26_6 (
    .a(i26[6]),
    .b(sum_25[6]),
    .c(cout_26[5]),
    .cout(cout_26[6]),
    .sum(sum_26[6]));
  AL_FADD comp26_60 (
    .a(1'b0),
    .b(sum_25[60]),
    .c(cout_26[59]),
    .cout(cout_26[60]),
    .sum(sum_26[60]));
  AL_FADD comp26_61 (
    .a(1'b0),
    .b(sum_25[61]),
    .c(cout_26[60]),
    .cout(cout_26[61]),
    .sum(sum_26[61]));
  AL_FADD comp26_62 (
    .a(1'b0),
    .b(sum_25[62]),
    .c(cout_26[61]),
    .cout(cout_26[62]),
    .sum(sum_26[62]));
  AL_FADD comp26_63 (
    .a(1'b0),
    .b(sum_25[63]),
    .c(cout_26[62]),
    .cout(cout_26[63]),
    .sum(sum_26[63]));
  AL_FADD comp26_7 (
    .a(i26[7]),
    .b(sum_25[7]),
    .c(cout_26[6]),
    .cout(cout_26[7]),
    .sum(sum_26[7]));
  AL_FADD comp26_8 (
    .a(i26[8]),
    .b(sum_25[8]),
    .c(cout_26[7]),
    .cout(cout_26[8]),
    .sum(sum_26[8]));
  AL_FADD comp26_9 (
    .a(i26[9]),
    .b(sum_25[9]),
    .c(cout_26[8]),
    .cout(cout_26[9]),
    .sum(sum_26[9]));
  AL_FADD comp27_0 (
    .a(i27[0]),
    .b(sum_26[0]),
    .c(1'b0),
    .cout(cout_27[0]),
    .sum(sum_27[0]));
  AL_FADD comp27_1 (
    .a(i27[1]),
    .b(sum_26[1]),
    .c(cout_27[0]),
    .cout(cout_27[1]),
    .sum(sum_27[1]));
  AL_FADD comp27_10 (
    .a(i27[10]),
    .b(sum_26[10]),
    .c(cout_27[9]),
    .cout(cout_27[10]),
    .sum(sum_27[10]));
  AL_FADD comp27_11 (
    .a(i27[11]),
    .b(sum_26[11]),
    .c(cout_27[10]),
    .cout(cout_27[11]),
    .sum(sum_27[11]));
  AL_FADD comp27_12 (
    .a(i27[12]),
    .b(sum_26[12]),
    .c(cout_27[11]),
    .cout(cout_27[12]),
    .sum(sum_27[12]));
  AL_FADD comp27_13 (
    .a(i27[13]),
    .b(sum_26[13]),
    .c(cout_27[12]),
    .cout(cout_27[13]),
    .sum(sum_27[13]));
  AL_FADD comp27_14 (
    .a(i27[14]),
    .b(sum_26[14]),
    .c(cout_27[13]),
    .cout(cout_27[14]),
    .sum(sum_27[14]));
  AL_FADD comp27_15 (
    .a(i27[15]),
    .b(sum_26[15]),
    .c(cout_27[14]),
    .cout(cout_27[15]),
    .sum(sum_27[15]));
  AL_FADD comp27_16 (
    .a(i27[16]),
    .b(sum_26[16]),
    .c(cout_27[15]),
    .cout(cout_27[16]),
    .sum(sum_27[16]));
  AL_FADD comp27_17 (
    .a(i27[17]),
    .b(sum_26[17]),
    .c(cout_27[16]),
    .cout(cout_27[17]),
    .sum(sum_27[17]));
  AL_FADD comp27_18 (
    .a(i27[18]),
    .b(sum_26[18]),
    .c(cout_27[17]),
    .cout(cout_27[18]),
    .sum(sum_27[18]));
  AL_FADD comp27_19 (
    .a(i27[19]),
    .b(sum_26[19]),
    .c(cout_27[18]),
    .cout(cout_27[19]),
    .sum(sum_27[19]));
  AL_FADD comp27_2 (
    .a(i27[2]),
    .b(sum_26[2]),
    .c(cout_27[1]),
    .cout(cout_27[2]),
    .sum(sum_27[2]));
  AL_FADD comp27_20 (
    .a(i27[20]),
    .b(sum_26[20]),
    .c(cout_27[19]),
    .cout(cout_27[20]),
    .sum(sum_27[20]));
  AL_FADD comp27_21 (
    .a(i27[21]),
    .b(sum_26[21]),
    .c(cout_27[20]),
    .cout(cout_27[21]),
    .sum(sum_27[21]));
  AL_FADD comp27_22 (
    .a(i27[22]),
    .b(sum_26[22]),
    .c(cout_27[21]),
    .cout(cout_27[22]),
    .sum(sum_27[22]));
  AL_FADD comp27_23 (
    .a(i27[23]),
    .b(sum_26[23]),
    .c(cout_27[22]),
    .cout(cout_27[23]),
    .sum(sum_27[23]));
  AL_FADD comp27_24 (
    .a(i27[24]),
    .b(sum_26[24]),
    .c(cout_27[23]),
    .cout(cout_27[24]),
    .sum(sum_27[24]));
  AL_FADD comp27_25 (
    .a(i27[25]),
    .b(sum_26[25]),
    .c(cout_27[24]),
    .cout(cout_27[25]),
    .sum(sum_27[25]));
  AL_FADD comp27_26 (
    .a(i27[26]),
    .b(sum_26[26]),
    .c(cout_27[25]),
    .cout(cout_27[26]),
    .sum(sum_27[26]));
  AL_FADD comp27_27 (
    .a(i27[27]),
    .b(sum_26[27]),
    .c(cout_27[26]),
    .cout(cout_27[27]),
    .sum(sum_27[27]));
  AL_FADD comp27_28 (
    .a(i27[28]),
    .b(sum_26[28]),
    .c(cout_27[27]),
    .cout(cout_27[28]),
    .sum(sum_27[28]));
  AL_FADD comp27_29 (
    .a(i27[29]),
    .b(sum_26[29]),
    .c(cout_27[28]),
    .cout(cout_27[29]),
    .sum(sum_27[29]));
  AL_FADD comp27_3 (
    .a(i27[3]),
    .b(sum_26[3]),
    .c(cout_27[2]),
    .cout(cout_27[3]),
    .sum(sum_27[3]));
  AL_FADD comp27_30 (
    .a(i27[30]),
    .b(sum_26[30]),
    .c(cout_27[29]),
    .cout(cout_27[30]),
    .sum(sum_27[30]));
  AL_FADD comp27_31 (
    .a(i27[31]),
    .b(sum_26[31]),
    .c(cout_27[30]),
    .cout(cout_27[31]),
    .sum(sum_27[31]));
  AL_FADD comp27_32 (
    .a(i27[32]),
    .b(sum_26[32]),
    .c(cout_27[31]),
    .cout(cout_27[32]),
    .sum(sum_27[32]));
  AL_FADD comp27_33 (
    .a(i27[33]),
    .b(sum_26[33]),
    .c(cout_27[32]),
    .cout(cout_27[33]),
    .sum(sum_27[33]));
  AL_FADD comp27_34 (
    .a(1'b0),
    .b(sum_26[34]),
    .c(cout_27[33]),
    .cout(cout_27[34]),
    .sum(sum_27[34]));
  AL_FADD comp27_35 (
    .a(1'b0),
    .b(sum_26[35]),
    .c(cout_27[34]),
    .cout(cout_27[35]),
    .sum(sum_27[35]));
  AL_FADD comp27_36 (
    .a(1'b0),
    .b(sum_26[36]),
    .c(cout_27[35]),
    .cout(cout_27[36]),
    .sum(sum_27[36]));
  AL_FADD comp27_37 (
    .a(1'b0),
    .b(sum_26[37]),
    .c(cout_27[36]),
    .cout(cout_27[37]),
    .sum(sum_27[37]));
  AL_FADD comp27_38 (
    .a(1'b0),
    .b(sum_26[38]),
    .c(cout_27[37]),
    .cout(cout_27[38]),
    .sum(sum_27[38]));
  AL_FADD comp27_39 (
    .a(1'b0),
    .b(sum_26[39]),
    .c(cout_27[38]),
    .cout(cout_27[39]),
    .sum(sum_27[39]));
  AL_FADD comp27_4 (
    .a(i27[4]),
    .b(sum_26[4]),
    .c(cout_27[3]),
    .cout(cout_27[4]),
    .sum(sum_27[4]));
  AL_FADD comp27_40 (
    .a(1'b0),
    .b(sum_26[40]),
    .c(cout_27[39]),
    .cout(cout_27[40]),
    .sum(sum_27[40]));
  AL_FADD comp27_41 (
    .a(1'b0),
    .b(sum_26[41]),
    .c(cout_27[40]),
    .cout(cout_27[41]),
    .sum(sum_27[41]));
  AL_FADD comp27_42 (
    .a(1'b0),
    .b(sum_26[42]),
    .c(cout_27[41]),
    .cout(cout_27[42]),
    .sum(sum_27[42]));
  AL_FADD comp27_43 (
    .a(1'b0),
    .b(sum_26[43]),
    .c(cout_27[42]),
    .cout(cout_27[43]),
    .sum(sum_27[43]));
  AL_FADD comp27_44 (
    .a(1'b0),
    .b(sum_26[44]),
    .c(cout_27[43]),
    .cout(cout_27[44]),
    .sum(sum_27[44]));
  AL_FADD comp27_45 (
    .a(1'b0),
    .b(sum_26[45]),
    .c(cout_27[44]),
    .cout(cout_27[45]),
    .sum(sum_27[45]));
  AL_FADD comp27_46 (
    .a(1'b0),
    .b(sum_26[46]),
    .c(cout_27[45]),
    .cout(cout_27[46]),
    .sum(sum_27[46]));
  AL_FADD comp27_47 (
    .a(1'b0),
    .b(sum_26[47]),
    .c(cout_27[46]),
    .cout(cout_27[47]),
    .sum(sum_27[47]));
  AL_FADD comp27_48 (
    .a(1'b0),
    .b(sum_26[48]),
    .c(cout_27[47]),
    .cout(cout_27[48]),
    .sum(sum_27[48]));
  AL_FADD comp27_49 (
    .a(1'b0),
    .b(sum_26[49]),
    .c(cout_27[48]),
    .cout(cout_27[49]),
    .sum(sum_27[49]));
  AL_FADD comp27_5 (
    .a(i27[5]),
    .b(sum_26[5]),
    .c(cout_27[4]),
    .cout(cout_27[5]),
    .sum(sum_27[5]));
  AL_FADD comp27_50 (
    .a(1'b0),
    .b(sum_26[50]),
    .c(cout_27[49]),
    .cout(cout_27[50]),
    .sum(sum_27[50]));
  AL_FADD comp27_51 (
    .a(1'b0),
    .b(sum_26[51]),
    .c(cout_27[50]),
    .cout(cout_27[51]),
    .sum(sum_27[51]));
  AL_FADD comp27_52 (
    .a(1'b0),
    .b(sum_26[52]),
    .c(cout_27[51]),
    .cout(cout_27[52]),
    .sum(sum_27[52]));
  AL_FADD comp27_53 (
    .a(1'b0),
    .b(sum_26[53]),
    .c(cout_27[52]),
    .cout(cout_27[53]),
    .sum(sum_27[53]));
  AL_FADD comp27_54 (
    .a(1'b0),
    .b(sum_26[54]),
    .c(cout_27[53]),
    .cout(cout_27[54]),
    .sum(sum_27[54]));
  AL_FADD comp27_55 (
    .a(1'b0),
    .b(sum_26[55]),
    .c(cout_27[54]),
    .cout(cout_27[55]),
    .sum(sum_27[55]));
  AL_FADD comp27_56 (
    .a(1'b0),
    .b(sum_26[56]),
    .c(cout_27[55]),
    .cout(cout_27[56]),
    .sum(sum_27[56]));
  AL_FADD comp27_57 (
    .a(1'b0),
    .b(sum_26[57]),
    .c(cout_27[56]),
    .cout(cout_27[57]),
    .sum(sum_27[57]));
  AL_FADD comp27_58 (
    .a(1'b0),
    .b(sum_26[58]),
    .c(cout_27[57]),
    .cout(cout_27[58]),
    .sum(sum_27[58]));
  AL_FADD comp27_59 (
    .a(1'b0),
    .b(sum_26[59]),
    .c(cout_27[58]),
    .cout(cout_27[59]),
    .sum(sum_27[59]));
  AL_FADD comp27_6 (
    .a(i27[6]),
    .b(sum_26[6]),
    .c(cout_27[5]),
    .cout(cout_27[6]),
    .sum(sum_27[6]));
  AL_FADD comp27_60 (
    .a(1'b0),
    .b(sum_26[60]),
    .c(cout_27[59]),
    .cout(cout_27[60]),
    .sum(sum_27[60]));
  AL_FADD comp27_61 (
    .a(1'b0),
    .b(sum_26[61]),
    .c(cout_27[60]),
    .cout(cout_27[61]),
    .sum(sum_27[61]));
  AL_FADD comp27_62 (
    .a(1'b0),
    .b(sum_26[62]),
    .c(cout_27[61]),
    .cout(cout_27[62]),
    .sum(sum_27[62]));
  AL_FADD comp27_63 (
    .a(1'b0),
    .b(sum_26[63]),
    .c(cout_27[62]),
    .cout(cout_27[63]),
    .sum(sum_27[63]));
  AL_FADD comp27_7 (
    .a(i27[7]),
    .b(sum_26[7]),
    .c(cout_27[6]),
    .cout(cout_27[7]),
    .sum(sum_27[7]));
  AL_FADD comp27_8 (
    .a(i27[8]),
    .b(sum_26[8]),
    .c(cout_27[7]),
    .cout(cout_27[8]),
    .sum(sum_27[8]));
  AL_FADD comp27_9 (
    .a(i27[9]),
    .b(sum_26[9]),
    .c(cout_27[8]),
    .cout(cout_27[9]),
    .sum(sum_27[9]));
  AL_FADD comp28_0 (
    .a(i28[0]),
    .b(sum_27[0]),
    .c(1'b0),
    .cout(cout_28[0]),
    .sum(sum_28[0]));
  AL_FADD comp28_1 (
    .a(i28[1]),
    .b(sum_27[1]),
    .c(cout_28[0]),
    .cout(cout_28[1]),
    .sum(sum_28[1]));
  AL_FADD comp28_10 (
    .a(i28[10]),
    .b(sum_27[10]),
    .c(cout_28[9]),
    .cout(cout_28[10]),
    .sum(sum_28[10]));
  AL_FADD comp28_11 (
    .a(i28[11]),
    .b(sum_27[11]),
    .c(cout_28[10]),
    .cout(cout_28[11]),
    .sum(sum_28[11]));
  AL_FADD comp28_12 (
    .a(i28[12]),
    .b(sum_27[12]),
    .c(cout_28[11]),
    .cout(cout_28[12]),
    .sum(sum_28[12]));
  AL_FADD comp28_13 (
    .a(i28[13]),
    .b(sum_27[13]),
    .c(cout_28[12]),
    .cout(cout_28[13]),
    .sum(sum_28[13]));
  AL_FADD comp28_14 (
    .a(i28[14]),
    .b(sum_27[14]),
    .c(cout_28[13]),
    .cout(cout_28[14]),
    .sum(sum_28[14]));
  AL_FADD comp28_15 (
    .a(i28[15]),
    .b(sum_27[15]),
    .c(cout_28[14]),
    .cout(cout_28[15]),
    .sum(sum_28[15]));
  AL_FADD comp28_16 (
    .a(i28[16]),
    .b(sum_27[16]),
    .c(cout_28[15]),
    .cout(cout_28[16]),
    .sum(sum_28[16]));
  AL_FADD comp28_17 (
    .a(i28[17]),
    .b(sum_27[17]),
    .c(cout_28[16]),
    .cout(cout_28[17]),
    .sum(sum_28[17]));
  AL_FADD comp28_18 (
    .a(i28[18]),
    .b(sum_27[18]),
    .c(cout_28[17]),
    .cout(cout_28[18]),
    .sum(sum_28[18]));
  AL_FADD comp28_19 (
    .a(i28[19]),
    .b(sum_27[19]),
    .c(cout_28[18]),
    .cout(cout_28[19]),
    .sum(sum_28[19]));
  AL_FADD comp28_2 (
    .a(i28[2]),
    .b(sum_27[2]),
    .c(cout_28[1]),
    .cout(cout_28[2]),
    .sum(sum_28[2]));
  AL_FADD comp28_20 (
    .a(i28[20]),
    .b(sum_27[20]),
    .c(cout_28[19]),
    .cout(cout_28[20]),
    .sum(sum_28[20]));
  AL_FADD comp28_21 (
    .a(i28[21]),
    .b(sum_27[21]),
    .c(cout_28[20]),
    .cout(cout_28[21]),
    .sum(sum_28[21]));
  AL_FADD comp28_22 (
    .a(i28[22]),
    .b(sum_27[22]),
    .c(cout_28[21]),
    .cout(cout_28[22]),
    .sum(sum_28[22]));
  AL_FADD comp28_23 (
    .a(i28[23]),
    .b(sum_27[23]),
    .c(cout_28[22]),
    .cout(cout_28[23]),
    .sum(sum_28[23]));
  AL_FADD comp28_24 (
    .a(i28[24]),
    .b(sum_27[24]),
    .c(cout_28[23]),
    .cout(cout_28[24]),
    .sum(sum_28[24]));
  AL_FADD comp28_25 (
    .a(i28[25]),
    .b(sum_27[25]),
    .c(cout_28[24]),
    .cout(cout_28[25]),
    .sum(sum_28[25]));
  AL_FADD comp28_26 (
    .a(i28[26]),
    .b(sum_27[26]),
    .c(cout_28[25]),
    .cout(cout_28[26]),
    .sum(sum_28[26]));
  AL_FADD comp28_27 (
    .a(i28[27]),
    .b(sum_27[27]),
    .c(cout_28[26]),
    .cout(cout_28[27]),
    .sum(sum_28[27]));
  AL_FADD comp28_28 (
    .a(i28[28]),
    .b(sum_27[28]),
    .c(cout_28[27]),
    .cout(cout_28[28]),
    .sum(sum_28[28]));
  AL_FADD comp28_29 (
    .a(i28[29]),
    .b(sum_27[29]),
    .c(cout_28[28]),
    .cout(cout_28[29]),
    .sum(sum_28[29]));
  AL_FADD comp28_3 (
    .a(i28[3]),
    .b(sum_27[3]),
    .c(cout_28[2]),
    .cout(cout_28[3]),
    .sum(sum_28[3]));
  AL_FADD comp28_30 (
    .a(i28[30]),
    .b(sum_27[30]),
    .c(cout_28[29]),
    .cout(cout_28[30]),
    .sum(sum_28[30]));
  AL_FADD comp28_31 (
    .a(i28[31]),
    .b(sum_27[31]),
    .c(cout_28[30]),
    .cout(cout_28[31]),
    .sum(sum_28[31]));
  AL_FADD comp28_32 (
    .a(i28[32]),
    .b(sum_27[32]),
    .c(cout_28[31]),
    .cout(cout_28[32]),
    .sum(sum_28[32]));
  AL_FADD comp28_33 (
    .a(1'b0),
    .b(sum_27[33]),
    .c(cout_28[32]),
    .cout(cout_28[33]),
    .sum(sum_28[33]));
  AL_FADD comp28_34 (
    .a(1'b0),
    .b(sum_27[34]),
    .c(cout_28[33]),
    .cout(cout_28[34]),
    .sum(sum_28[34]));
  AL_FADD comp28_35 (
    .a(1'b0),
    .b(sum_27[35]),
    .c(cout_28[34]),
    .cout(cout_28[35]),
    .sum(sum_28[35]));
  AL_FADD comp28_36 (
    .a(1'b0),
    .b(sum_27[36]),
    .c(cout_28[35]),
    .cout(cout_28[36]),
    .sum(sum_28[36]));
  AL_FADD comp28_37 (
    .a(1'b0),
    .b(sum_27[37]),
    .c(cout_28[36]),
    .cout(cout_28[37]),
    .sum(sum_28[37]));
  AL_FADD comp28_38 (
    .a(1'b0),
    .b(sum_27[38]),
    .c(cout_28[37]),
    .cout(cout_28[38]),
    .sum(sum_28[38]));
  AL_FADD comp28_39 (
    .a(1'b0),
    .b(sum_27[39]),
    .c(cout_28[38]),
    .cout(cout_28[39]),
    .sum(sum_28[39]));
  AL_FADD comp28_4 (
    .a(i28[4]),
    .b(sum_27[4]),
    .c(cout_28[3]),
    .cout(cout_28[4]),
    .sum(sum_28[4]));
  AL_FADD comp28_40 (
    .a(1'b0),
    .b(sum_27[40]),
    .c(cout_28[39]),
    .cout(cout_28[40]),
    .sum(sum_28[40]));
  AL_FADD comp28_41 (
    .a(1'b0),
    .b(sum_27[41]),
    .c(cout_28[40]),
    .cout(cout_28[41]),
    .sum(sum_28[41]));
  AL_FADD comp28_42 (
    .a(1'b0),
    .b(sum_27[42]),
    .c(cout_28[41]),
    .cout(cout_28[42]),
    .sum(sum_28[42]));
  AL_FADD comp28_43 (
    .a(1'b0),
    .b(sum_27[43]),
    .c(cout_28[42]),
    .cout(cout_28[43]),
    .sum(sum_28[43]));
  AL_FADD comp28_44 (
    .a(1'b0),
    .b(sum_27[44]),
    .c(cout_28[43]),
    .cout(cout_28[44]),
    .sum(sum_28[44]));
  AL_FADD comp28_45 (
    .a(1'b0),
    .b(sum_27[45]),
    .c(cout_28[44]),
    .cout(cout_28[45]),
    .sum(sum_28[45]));
  AL_FADD comp28_46 (
    .a(1'b0),
    .b(sum_27[46]),
    .c(cout_28[45]),
    .cout(cout_28[46]),
    .sum(sum_28[46]));
  AL_FADD comp28_47 (
    .a(1'b0),
    .b(sum_27[47]),
    .c(cout_28[46]),
    .cout(cout_28[47]),
    .sum(sum_28[47]));
  AL_FADD comp28_48 (
    .a(1'b0),
    .b(sum_27[48]),
    .c(cout_28[47]),
    .cout(cout_28[48]),
    .sum(sum_28[48]));
  AL_FADD comp28_49 (
    .a(1'b0),
    .b(sum_27[49]),
    .c(cout_28[48]),
    .cout(cout_28[49]),
    .sum(sum_28[49]));
  AL_FADD comp28_5 (
    .a(i28[5]),
    .b(sum_27[5]),
    .c(cout_28[4]),
    .cout(cout_28[5]),
    .sum(sum_28[5]));
  AL_FADD comp28_50 (
    .a(1'b0),
    .b(sum_27[50]),
    .c(cout_28[49]),
    .cout(cout_28[50]),
    .sum(sum_28[50]));
  AL_FADD comp28_51 (
    .a(1'b0),
    .b(sum_27[51]),
    .c(cout_28[50]),
    .cout(cout_28[51]),
    .sum(sum_28[51]));
  AL_FADD comp28_52 (
    .a(1'b0),
    .b(sum_27[52]),
    .c(cout_28[51]),
    .cout(cout_28[52]),
    .sum(sum_28[52]));
  AL_FADD comp28_53 (
    .a(1'b0),
    .b(sum_27[53]),
    .c(cout_28[52]),
    .cout(cout_28[53]),
    .sum(sum_28[53]));
  AL_FADD comp28_54 (
    .a(1'b0),
    .b(sum_27[54]),
    .c(cout_28[53]),
    .cout(cout_28[54]),
    .sum(sum_28[54]));
  AL_FADD comp28_55 (
    .a(1'b0),
    .b(sum_27[55]),
    .c(cout_28[54]),
    .cout(cout_28[55]),
    .sum(sum_28[55]));
  AL_FADD comp28_56 (
    .a(1'b0),
    .b(sum_27[56]),
    .c(cout_28[55]),
    .cout(cout_28[56]),
    .sum(sum_28[56]));
  AL_FADD comp28_57 (
    .a(1'b0),
    .b(sum_27[57]),
    .c(cout_28[56]),
    .cout(cout_28[57]),
    .sum(sum_28[57]));
  AL_FADD comp28_58 (
    .a(1'b0),
    .b(sum_27[58]),
    .c(cout_28[57]),
    .cout(cout_28[58]),
    .sum(sum_28[58]));
  AL_FADD comp28_59 (
    .a(1'b0),
    .b(sum_27[59]),
    .c(cout_28[58]),
    .cout(cout_28[59]),
    .sum(sum_28[59]));
  AL_FADD comp28_6 (
    .a(i28[6]),
    .b(sum_27[6]),
    .c(cout_28[5]),
    .cout(cout_28[6]),
    .sum(sum_28[6]));
  AL_FADD comp28_60 (
    .a(1'b0),
    .b(sum_27[60]),
    .c(cout_28[59]),
    .cout(cout_28[60]),
    .sum(sum_28[60]));
  AL_FADD comp28_61 (
    .a(1'b0),
    .b(sum_27[61]),
    .c(cout_28[60]),
    .cout(cout_28[61]),
    .sum(sum_28[61]));
  AL_FADD comp28_62 (
    .a(1'b0),
    .b(sum_27[62]),
    .c(cout_28[61]),
    .cout(cout_28[62]),
    .sum(sum_28[62]));
  AL_FADD comp28_63 (
    .a(1'b0),
    .b(sum_27[63]),
    .c(cout_28[62]),
    .cout(cout_28[63]),
    .sum(sum_28[63]));
  AL_FADD comp28_7 (
    .a(i28[7]),
    .b(sum_27[7]),
    .c(cout_28[6]),
    .cout(cout_28[7]),
    .sum(sum_28[7]));
  AL_FADD comp28_8 (
    .a(i28[8]),
    .b(sum_27[8]),
    .c(cout_28[7]),
    .cout(cout_28[8]),
    .sum(sum_28[8]));
  AL_FADD comp28_9 (
    .a(i28[9]),
    .b(sum_27[9]),
    .c(cout_28[8]),
    .cout(cout_28[9]),
    .sum(sum_28[9]));
  AL_FADD comp29_0 (
    .a(i29[0]),
    .b(sum_28[0]),
    .c(1'b0),
    .cout(cout_29[0]),
    .sum(sum_29[0]));
  AL_FADD comp29_1 (
    .a(i29[1]),
    .b(sum_28[1]),
    .c(cout_29[0]),
    .cout(cout_29[1]),
    .sum(sum_29[1]));
  AL_FADD comp29_10 (
    .a(i29[10]),
    .b(sum_28[10]),
    .c(cout_29[9]),
    .cout(cout_29[10]),
    .sum(sum_29[10]));
  AL_FADD comp29_11 (
    .a(i29[11]),
    .b(sum_28[11]),
    .c(cout_29[10]),
    .cout(cout_29[11]),
    .sum(sum_29[11]));
  AL_FADD comp29_12 (
    .a(i29[12]),
    .b(sum_28[12]),
    .c(cout_29[11]),
    .cout(cout_29[12]),
    .sum(sum_29[12]));
  AL_FADD comp29_13 (
    .a(i29[13]),
    .b(sum_28[13]),
    .c(cout_29[12]),
    .cout(cout_29[13]),
    .sum(sum_29[13]));
  AL_FADD comp29_14 (
    .a(i29[14]),
    .b(sum_28[14]),
    .c(cout_29[13]),
    .cout(cout_29[14]),
    .sum(sum_29[14]));
  AL_FADD comp29_15 (
    .a(i29[15]),
    .b(sum_28[15]),
    .c(cout_29[14]),
    .cout(cout_29[15]),
    .sum(sum_29[15]));
  AL_FADD comp29_16 (
    .a(i29[16]),
    .b(sum_28[16]),
    .c(cout_29[15]),
    .cout(cout_29[16]),
    .sum(sum_29[16]));
  AL_FADD comp29_17 (
    .a(i29[17]),
    .b(sum_28[17]),
    .c(cout_29[16]),
    .cout(cout_29[17]),
    .sum(sum_29[17]));
  AL_FADD comp29_18 (
    .a(i29[18]),
    .b(sum_28[18]),
    .c(cout_29[17]),
    .cout(cout_29[18]),
    .sum(sum_29[18]));
  AL_FADD comp29_19 (
    .a(i29[19]),
    .b(sum_28[19]),
    .c(cout_29[18]),
    .cout(cout_29[19]),
    .sum(sum_29[19]));
  AL_FADD comp29_2 (
    .a(i29[2]),
    .b(sum_28[2]),
    .c(cout_29[1]),
    .cout(cout_29[2]),
    .sum(sum_29[2]));
  AL_FADD comp29_20 (
    .a(i29[20]),
    .b(sum_28[20]),
    .c(cout_29[19]),
    .cout(cout_29[20]),
    .sum(sum_29[20]));
  AL_FADD comp29_21 (
    .a(i29[21]),
    .b(sum_28[21]),
    .c(cout_29[20]),
    .cout(cout_29[21]),
    .sum(sum_29[21]));
  AL_FADD comp29_22 (
    .a(i29[22]),
    .b(sum_28[22]),
    .c(cout_29[21]),
    .cout(cout_29[22]),
    .sum(sum_29[22]));
  AL_FADD comp29_23 (
    .a(i29[23]),
    .b(sum_28[23]),
    .c(cout_29[22]),
    .cout(cout_29[23]),
    .sum(sum_29[23]));
  AL_FADD comp29_24 (
    .a(i29[24]),
    .b(sum_28[24]),
    .c(cout_29[23]),
    .cout(cout_29[24]),
    .sum(sum_29[24]));
  AL_FADD comp29_25 (
    .a(i29[25]),
    .b(sum_28[25]),
    .c(cout_29[24]),
    .cout(cout_29[25]),
    .sum(sum_29[25]));
  AL_FADD comp29_26 (
    .a(i29[26]),
    .b(sum_28[26]),
    .c(cout_29[25]),
    .cout(cout_29[26]),
    .sum(sum_29[26]));
  AL_FADD comp29_27 (
    .a(i29[27]),
    .b(sum_28[27]),
    .c(cout_29[26]),
    .cout(cout_29[27]),
    .sum(sum_29[27]));
  AL_FADD comp29_28 (
    .a(i29[28]),
    .b(sum_28[28]),
    .c(cout_29[27]),
    .cout(cout_29[28]),
    .sum(sum_29[28]));
  AL_FADD comp29_29 (
    .a(i29[29]),
    .b(sum_28[29]),
    .c(cout_29[28]),
    .cout(cout_29[29]),
    .sum(sum_29[29]));
  AL_FADD comp29_3 (
    .a(i29[3]),
    .b(sum_28[3]),
    .c(cout_29[2]),
    .cout(cout_29[3]),
    .sum(sum_29[3]));
  AL_FADD comp29_30 (
    .a(i29[30]),
    .b(sum_28[30]),
    .c(cout_29[29]),
    .cout(cout_29[30]),
    .sum(sum_29[30]));
  AL_FADD comp29_31 (
    .a(i29[31]),
    .b(sum_28[31]),
    .c(cout_29[30]),
    .cout(cout_29[31]),
    .sum(sum_29[31]));
  AL_FADD comp29_32 (
    .a(1'b0),
    .b(sum_28[32]),
    .c(cout_29[31]),
    .cout(cout_29[32]),
    .sum(sum_29[32]));
  AL_FADD comp29_33 (
    .a(1'b0),
    .b(sum_28[33]),
    .c(cout_29[32]),
    .cout(cout_29[33]),
    .sum(sum_29[33]));
  AL_FADD comp29_34 (
    .a(1'b0),
    .b(sum_28[34]),
    .c(cout_29[33]),
    .cout(cout_29[34]),
    .sum(sum_29[34]));
  AL_FADD comp29_35 (
    .a(1'b0),
    .b(sum_28[35]),
    .c(cout_29[34]),
    .cout(cout_29[35]),
    .sum(sum_29[35]));
  AL_FADD comp29_36 (
    .a(1'b0),
    .b(sum_28[36]),
    .c(cout_29[35]),
    .cout(cout_29[36]),
    .sum(sum_29[36]));
  AL_FADD comp29_37 (
    .a(1'b0),
    .b(sum_28[37]),
    .c(cout_29[36]),
    .cout(cout_29[37]),
    .sum(sum_29[37]));
  AL_FADD comp29_38 (
    .a(1'b0),
    .b(sum_28[38]),
    .c(cout_29[37]),
    .cout(cout_29[38]),
    .sum(sum_29[38]));
  AL_FADD comp29_39 (
    .a(1'b0),
    .b(sum_28[39]),
    .c(cout_29[38]),
    .cout(cout_29[39]),
    .sum(sum_29[39]));
  AL_FADD comp29_4 (
    .a(i29[4]),
    .b(sum_28[4]),
    .c(cout_29[3]),
    .cout(cout_29[4]),
    .sum(sum_29[4]));
  AL_FADD comp29_40 (
    .a(1'b0),
    .b(sum_28[40]),
    .c(cout_29[39]),
    .cout(cout_29[40]),
    .sum(sum_29[40]));
  AL_FADD comp29_41 (
    .a(1'b0),
    .b(sum_28[41]),
    .c(cout_29[40]),
    .cout(cout_29[41]),
    .sum(sum_29[41]));
  AL_FADD comp29_42 (
    .a(1'b0),
    .b(sum_28[42]),
    .c(cout_29[41]),
    .cout(cout_29[42]),
    .sum(sum_29[42]));
  AL_FADD comp29_43 (
    .a(1'b0),
    .b(sum_28[43]),
    .c(cout_29[42]),
    .cout(cout_29[43]),
    .sum(sum_29[43]));
  AL_FADD comp29_44 (
    .a(1'b0),
    .b(sum_28[44]),
    .c(cout_29[43]),
    .cout(cout_29[44]),
    .sum(sum_29[44]));
  AL_FADD comp29_45 (
    .a(1'b0),
    .b(sum_28[45]),
    .c(cout_29[44]),
    .cout(cout_29[45]),
    .sum(sum_29[45]));
  AL_FADD comp29_46 (
    .a(1'b0),
    .b(sum_28[46]),
    .c(cout_29[45]),
    .cout(cout_29[46]),
    .sum(sum_29[46]));
  AL_FADD comp29_47 (
    .a(1'b0),
    .b(sum_28[47]),
    .c(cout_29[46]),
    .cout(cout_29[47]),
    .sum(sum_29[47]));
  AL_FADD comp29_48 (
    .a(1'b0),
    .b(sum_28[48]),
    .c(cout_29[47]),
    .cout(cout_29[48]),
    .sum(sum_29[48]));
  AL_FADD comp29_49 (
    .a(1'b0),
    .b(sum_28[49]),
    .c(cout_29[48]),
    .cout(cout_29[49]),
    .sum(sum_29[49]));
  AL_FADD comp29_5 (
    .a(i29[5]),
    .b(sum_28[5]),
    .c(cout_29[4]),
    .cout(cout_29[5]),
    .sum(sum_29[5]));
  AL_FADD comp29_50 (
    .a(1'b0),
    .b(sum_28[50]),
    .c(cout_29[49]),
    .cout(cout_29[50]),
    .sum(sum_29[50]));
  AL_FADD comp29_51 (
    .a(1'b0),
    .b(sum_28[51]),
    .c(cout_29[50]),
    .cout(cout_29[51]),
    .sum(sum_29[51]));
  AL_FADD comp29_52 (
    .a(1'b0),
    .b(sum_28[52]),
    .c(cout_29[51]),
    .cout(cout_29[52]),
    .sum(sum_29[52]));
  AL_FADD comp29_53 (
    .a(1'b0),
    .b(sum_28[53]),
    .c(cout_29[52]),
    .cout(cout_29[53]),
    .sum(sum_29[53]));
  AL_FADD comp29_54 (
    .a(1'b0),
    .b(sum_28[54]),
    .c(cout_29[53]),
    .cout(cout_29[54]),
    .sum(sum_29[54]));
  AL_FADD comp29_55 (
    .a(1'b0),
    .b(sum_28[55]),
    .c(cout_29[54]),
    .cout(cout_29[55]),
    .sum(sum_29[55]));
  AL_FADD comp29_56 (
    .a(1'b0),
    .b(sum_28[56]),
    .c(cout_29[55]),
    .cout(cout_29[56]),
    .sum(sum_29[56]));
  AL_FADD comp29_57 (
    .a(1'b0),
    .b(sum_28[57]),
    .c(cout_29[56]),
    .cout(cout_29[57]),
    .sum(sum_29[57]));
  AL_FADD comp29_58 (
    .a(1'b0),
    .b(sum_28[58]),
    .c(cout_29[57]),
    .cout(cout_29[58]),
    .sum(sum_29[58]));
  AL_FADD comp29_59 (
    .a(1'b0),
    .b(sum_28[59]),
    .c(cout_29[58]),
    .cout(cout_29[59]),
    .sum(sum_29[59]));
  AL_FADD comp29_6 (
    .a(i29[6]),
    .b(sum_28[6]),
    .c(cout_29[5]),
    .cout(cout_29[6]),
    .sum(sum_29[6]));
  AL_FADD comp29_60 (
    .a(1'b0),
    .b(sum_28[60]),
    .c(cout_29[59]),
    .cout(cout_29[60]),
    .sum(sum_29[60]));
  AL_FADD comp29_61 (
    .a(1'b0),
    .b(sum_28[61]),
    .c(cout_29[60]),
    .cout(cout_29[61]),
    .sum(sum_29[61]));
  AL_FADD comp29_62 (
    .a(1'b0),
    .b(sum_28[62]),
    .c(cout_29[61]),
    .cout(cout_29[62]),
    .sum(sum_29[62]));
  AL_FADD comp29_63 (
    .a(1'b0),
    .b(sum_28[63]),
    .c(cout_29[62]),
    .cout(cout_29[63]),
    .sum(sum_29[63]));
  AL_FADD comp29_7 (
    .a(i29[7]),
    .b(sum_28[7]),
    .c(cout_29[6]),
    .cout(cout_29[7]),
    .sum(sum_29[7]));
  AL_FADD comp29_8 (
    .a(i29[8]),
    .b(sum_28[8]),
    .c(cout_29[7]),
    .cout(cout_29[8]),
    .sum(sum_29[8]));
  AL_FADD comp29_9 (
    .a(i29[9]),
    .b(sum_28[9]),
    .c(cout_29[8]),
    .cout(cout_29[9]),
    .sum(sum_29[9]));
  AL_FADD comp2_0 (
    .a(i2[0]),
    .b(sum_1[0]),
    .c(1'b0),
    .cout(cout_2[0]),
    .sum(sum_2[0]));
  AL_FADD comp2_1 (
    .a(i2[1]),
    .b(sum_1[1]),
    .c(cout_2[0]),
    .cout(cout_2[1]),
    .sum(sum_2[1]));
  AL_FADD comp2_10 (
    .a(i2[10]),
    .b(sum_1[10]),
    .c(cout_2[9]),
    .cout(cout_2[10]),
    .sum(sum_2[10]));
  AL_FADD comp2_11 (
    .a(i2[11]),
    .b(sum_1[11]),
    .c(cout_2[10]),
    .cout(cout_2[11]),
    .sum(sum_2[11]));
  AL_FADD comp2_12 (
    .a(i2[12]),
    .b(sum_1[12]),
    .c(cout_2[11]),
    .cout(cout_2[12]),
    .sum(sum_2[12]));
  AL_FADD comp2_13 (
    .a(i2[13]),
    .b(sum_1[13]),
    .c(cout_2[12]),
    .cout(cout_2[13]),
    .sum(sum_2[13]));
  AL_FADD comp2_14 (
    .a(i2[14]),
    .b(sum_1[14]),
    .c(cout_2[13]),
    .cout(cout_2[14]),
    .sum(sum_2[14]));
  AL_FADD comp2_15 (
    .a(i2[15]),
    .b(sum_1[15]),
    .c(cout_2[14]),
    .cout(cout_2[15]),
    .sum(sum_2[15]));
  AL_FADD comp2_16 (
    .a(i2[16]),
    .b(sum_1[16]),
    .c(cout_2[15]),
    .cout(cout_2[16]),
    .sum(sum_2[16]));
  AL_FADD comp2_17 (
    .a(i2[17]),
    .b(sum_1[17]),
    .c(cout_2[16]),
    .cout(cout_2[17]),
    .sum(sum_2[17]));
  AL_FADD comp2_18 (
    .a(i2[18]),
    .b(sum_1[18]),
    .c(cout_2[17]),
    .cout(cout_2[18]),
    .sum(sum_2[18]));
  AL_FADD comp2_19 (
    .a(i2[19]),
    .b(sum_1[19]),
    .c(cout_2[18]),
    .cout(cout_2[19]),
    .sum(sum_2[19]));
  AL_FADD comp2_2 (
    .a(i2[2]),
    .b(sum_1[2]),
    .c(cout_2[1]),
    .cout(cout_2[2]),
    .sum(sum_2[2]));
  AL_FADD comp2_20 (
    .a(i2[20]),
    .b(sum_1[20]),
    .c(cout_2[19]),
    .cout(cout_2[20]),
    .sum(sum_2[20]));
  AL_FADD comp2_21 (
    .a(i2[21]),
    .b(sum_1[21]),
    .c(cout_2[20]),
    .cout(cout_2[21]),
    .sum(sum_2[21]));
  AL_FADD comp2_22 (
    .a(i2[22]),
    .b(sum_1[22]),
    .c(cout_2[21]),
    .cout(cout_2[22]),
    .sum(sum_2[22]));
  AL_FADD comp2_23 (
    .a(i2[23]),
    .b(sum_1[23]),
    .c(cout_2[22]),
    .cout(cout_2[23]),
    .sum(sum_2[23]));
  AL_FADD comp2_24 (
    .a(i2[24]),
    .b(sum_1[24]),
    .c(cout_2[23]),
    .cout(cout_2[24]),
    .sum(sum_2[24]));
  AL_FADD comp2_25 (
    .a(i2[25]),
    .b(sum_1[25]),
    .c(cout_2[24]),
    .cout(cout_2[25]),
    .sum(sum_2[25]));
  AL_FADD comp2_26 (
    .a(i2[26]),
    .b(sum_1[26]),
    .c(cout_2[25]),
    .cout(cout_2[26]),
    .sum(sum_2[26]));
  AL_FADD comp2_27 (
    .a(i2[27]),
    .b(sum_1[27]),
    .c(cout_2[26]),
    .cout(cout_2[27]),
    .sum(sum_2[27]));
  AL_FADD comp2_28 (
    .a(i2[28]),
    .b(sum_1[28]),
    .c(cout_2[27]),
    .cout(cout_2[28]),
    .sum(sum_2[28]));
  AL_FADD comp2_29 (
    .a(i2[29]),
    .b(sum_1[29]),
    .c(cout_2[28]),
    .cout(cout_2[29]),
    .sum(sum_2[29]));
  AL_FADD comp2_3 (
    .a(i2[3]),
    .b(sum_1[3]),
    .c(cout_2[2]),
    .cout(cout_2[3]),
    .sum(sum_2[3]));
  AL_FADD comp2_30 (
    .a(i2[30]),
    .b(sum_1[30]),
    .c(cout_2[29]),
    .cout(cout_2[30]),
    .sum(sum_2[30]));
  AL_FADD comp2_31 (
    .a(i2[31]),
    .b(sum_1[31]),
    .c(cout_2[30]),
    .cout(cout_2[31]),
    .sum(sum_2[31]));
  AL_FADD comp2_32 (
    .a(i2[32]),
    .b(sum_1[32]),
    .c(cout_2[31]),
    .cout(cout_2[32]),
    .sum(sum_2[32]));
  AL_FADD comp2_33 (
    .a(i2[33]),
    .b(sum_1[33]),
    .c(cout_2[32]),
    .cout(cout_2[33]),
    .sum(sum_2[33]));
  AL_FADD comp2_34 (
    .a(i2[34]),
    .b(sum_1[34]),
    .c(cout_2[33]),
    .cout(cout_2[34]),
    .sum(sum_2[34]));
  AL_FADD comp2_35 (
    .a(i2[35]),
    .b(sum_1[35]),
    .c(cout_2[34]),
    .cout(cout_2[35]),
    .sum(sum_2[35]));
  AL_FADD comp2_36 (
    .a(i2[36]),
    .b(sum_1[36]),
    .c(cout_2[35]),
    .cout(cout_2[36]),
    .sum(sum_2[36]));
  AL_FADD comp2_37 (
    .a(i2[37]),
    .b(sum_1[37]),
    .c(cout_2[36]),
    .cout(cout_2[37]),
    .sum(sum_2[37]));
  AL_FADD comp2_38 (
    .a(i2[38]),
    .b(sum_1[38]),
    .c(cout_2[37]),
    .cout(cout_2[38]),
    .sum(sum_2[38]));
  AL_FADD comp2_39 (
    .a(i2[39]),
    .b(sum_1[39]),
    .c(cout_2[38]),
    .cout(cout_2[39]),
    .sum(sum_2[39]));
  AL_FADD comp2_4 (
    .a(i2[4]),
    .b(sum_1[4]),
    .c(cout_2[3]),
    .cout(cout_2[4]),
    .sum(sum_2[4]));
  AL_FADD comp2_40 (
    .a(i2[40]),
    .b(sum_1[40]),
    .c(cout_2[39]),
    .cout(cout_2[40]),
    .sum(sum_2[40]));
  AL_FADD comp2_41 (
    .a(i2[41]),
    .b(sum_1[41]),
    .c(cout_2[40]),
    .cout(cout_2[41]),
    .sum(sum_2[41]));
  AL_FADD comp2_42 (
    .a(i2[42]),
    .b(sum_1[42]),
    .c(cout_2[41]),
    .cout(cout_2[42]),
    .sum(sum_2[42]));
  AL_FADD comp2_43 (
    .a(i2[43]),
    .b(sum_1[43]),
    .c(cout_2[42]),
    .cout(cout_2[43]),
    .sum(sum_2[43]));
  AL_FADD comp2_44 (
    .a(i2[44]),
    .b(sum_1[44]),
    .c(cout_2[43]),
    .cout(cout_2[44]),
    .sum(sum_2[44]));
  AL_FADD comp2_45 (
    .a(i2[45]),
    .b(sum_1[45]),
    .c(cout_2[44]),
    .cout(cout_2[45]),
    .sum(sum_2[45]));
  AL_FADD comp2_46 (
    .a(i2[46]),
    .b(sum_1[46]),
    .c(cout_2[45]),
    .cout(cout_2[46]),
    .sum(sum_2[46]));
  AL_FADD comp2_47 (
    .a(i2[47]),
    .b(sum_1[47]),
    .c(cout_2[46]),
    .cout(cout_2[47]),
    .sum(sum_2[47]));
  AL_FADD comp2_48 (
    .a(i2[48]),
    .b(sum_1[48]),
    .c(cout_2[47]),
    .cout(cout_2[48]),
    .sum(sum_2[48]));
  AL_FADD comp2_49 (
    .a(i2[49]),
    .b(sum_1[49]),
    .c(cout_2[48]),
    .cout(cout_2[49]),
    .sum(sum_2[49]));
  AL_FADD comp2_5 (
    .a(i2[5]),
    .b(sum_1[5]),
    .c(cout_2[4]),
    .cout(cout_2[5]),
    .sum(sum_2[5]));
  AL_FADD comp2_50 (
    .a(i2[50]),
    .b(sum_1[50]),
    .c(cout_2[49]),
    .cout(cout_2[50]),
    .sum(sum_2[50]));
  AL_FADD comp2_51 (
    .a(i2[51]),
    .b(sum_1[51]),
    .c(cout_2[50]),
    .cout(cout_2[51]),
    .sum(sum_2[51]));
  AL_FADD comp2_52 (
    .a(i2[52]),
    .b(sum_1[52]),
    .c(cout_2[51]),
    .cout(cout_2[52]),
    .sum(sum_2[52]));
  AL_FADD comp2_53 (
    .a(i2[53]),
    .b(sum_1[53]),
    .c(cout_2[52]),
    .cout(cout_2[53]),
    .sum(sum_2[53]));
  AL_FADD comp2_54 (
    .a(i2[54]),
    .b(sum_1[54]),
    .c(cout_2[53]),
    .cout(cout_2[54]),
    .sum(sum_2[54]));
  AL_FADD comp2_55 (
    .a(i2[55]),
    .b(sum_1[55]),
    .c(cout_2[54]),
    .cout(cout_2[55]),
    .sum(sum_2[55]));
  AL_FADD comp2_56 (
    .a(i2[56]),
    .b(sum_1[56]),
    .c(cout_2[55]),
    .cout(cout_2[56]),
    .sum(sum_2[56]));
  AL_FADD comp2_57 (
    .a(i2[57]),
    .b(sum_1[57]),
    .c(cout_2[56]),
    .cout(cout_2[57]),
    .sum(sum_2[57]));
  AL_FADD comp2_58 (
    .a(i2[58]),
    .b(sum_1[58]),
    .c(cout_2[57]),
    .cout(cout_2[58]),
    .sum(sum_2[58]));
  AL_FADD comp2_59 (
    .a(1'b0),
    .b(sum_1[59]),
    .c(cout_2[58]),
    .cout(cout_2[59]),
    .sum(sum_2[59]));
  AL_FADD comp2_6 (
    .a(i2[6]),
    .b(sum_1[6]),
    .c(cout_2[5]),
    .cout(cout_2[6]),
    .sum(sum_2[6]));
  AL_FADD comp2_60 (
    .a(1'b0),
    .b(sum_1[60]),
    .c(cout_2[59]),
    .cout(cout_2[60]),
    .sum(sum_2[60]));
  AL_FADD comp2_61 (
    .a(1'b0),
    .b(sum_1[61]),
    .c(cout_2[60]),
    .cout(cout_2[61]),
    .sum(sum_2[61]));
  AL_FADD comp2_62 (
    .a(1'b0),
    .b(sum_1[62]),
    .c(cout_2[61]),
    .cout(cout_2[62]),
    .sum(sum_2[62]));
  AL_FADD comp2_63 (
    .a(1'b0),
    .b(cout_1[62]),
    .c(cout_2[62]),
    .cout(cout_2[63]),
    .sum(sum_2[63]));
  AL_FADD comp2_7 (
    .a(i2[7]),
    .b(sum_1[7]),
    .c(cout_2[6]),
    .cout(cout_2[7]),
    .sum(sum_2[7]));
  AL_FADD comp2_8 (
    .a(i2[8]),
    .b(sum_1[8]),
    .c(cout_2[7]),
    .cout(cout_2[8]),
    .sum(sum_2[8]));
  AL_FADD comp2_9 (
    .a(i2[9]),
    .b(sum_1[9]),
    .c(cout_2[8]),
    .cout(cout_2[9]),
    .sum(sum_2[9]));
  AL_FADD comp30_0 (
    .a(i30[0]),
    .b(sum_29[0]),
    .c(1'b0),
    .cout(cout_30[0]),
    .sum(sum_30[0]));
  AL_FADD comp30_1 (
    .a(i30[1]),
    .b(sum_29[1]),
    .c(cout_30[0]),
    .cout(cout_30[1]),
    .sum(sum_30[1]));
  AL_FADD comp30_10 (
    .a(i30[10]),
    .b(sum_29[10]),
    .c(cout_30[9]),
    .cout(cout_30[10]),
    .sum(sum_30[10]));
  AL_FADD comp30_11 (
    .a(i30[11]),
    .b(sum_29[11]),
    .c(cout_30[10]),
    .cout(cout_30[11]),
    .sum(sum_30[11]));
  AL_FADD comp30_12 (
    .a(i30[12]),
    .b(sum_29[12]),
    .c(cout_30[11]),
    .cout(cout_30[12]),
    .sum(sum_30[12]));
  AL_FADD comp30_13 (
    .a(i30[13]),
    .b(sum_29[13]),
    .c(cout_30[12]),
    .cout(cout_30[13]),
    .sum(sum_30[13]));
  AL_FADD comp30_14 (
    .a(i30[14]),
    .b(sum_29[14]),
    .c(cout_30[13]),
    .cout(cout_30[14]),
    .sum(sum_30[14]));
  AL_FADD comp30_15 (
    .a(i30[15]),
    .b(sum_29[15]),
    .c(cout_30[14]),
    .cout(cout_30[15]),
    .sum(sum_30[15]));
  AL_FADD comp30_16 (
    .a(i30[16]),
    .b(sum_29[16]),
    .c(cout_30[15]),
    .cout(cout_30[16]),
    .sum(sum_30[16]));
  AL_FADD comp30_17 (
    .a(i30[17]),
    .b(sum_29[17]),
    .c(cout_30[16]),
    .cout(cout_30[17]),
    .sum(sum_30[17]));
  AL_FADD comp30_18 (
    .a(i30[18]),
    .b(sum_29[18]),
    .c(cout_30[17]),
    .cout(cout_30[18]),
    .sum(sum_30[18]));
  AL_FADD comp30_19 (
    .a(i30[19]),
    .b(sum_29[19]),
    .c(cout_30[18]),
    .cout(cout_30[19]),
    .sum(sum_30[19]));
  AL_FADD comp30_2 (
    .a(i30[2]),
    .b(sum_29[2]),
    .c(cout_30[1]),
    .cout(cout_30[2]),
    .sum(sum_30[2]));
  AL_FADD comp30_20 (
    .a(i30[20]),
    .b(sum_29[20]),
    .c(cout_30[19]),
    .cout(cout_30[20]),
    .sum(sum_30[20]));
  AL_FADD comp30_21 (
    .a(i30[21]),
    .b(sum_29[21]),
    .c(cout_30[20]),
    .cout(cout_30[21]),
    .sum(sum_30[21]));
  AL_FADD comp30_22 (
    .a(i30[22]),
    .b(sum_29[22]),
    .c(cout_30[21]),
    .cout(cout_30[22]),
    .sum(sum_30[22]));
  AL_FADD comp30_23 (
    .a(i30[23]),
    .b(sum_29[23]),
    .c(cout_30[22]),
    .cout(cout_30[23]),
    .sum(sum_30[23]));
  AL_FADD comp30_24 (
    .a(i30[24]),
    .b(sum_29[24]),
    .c(cout_30[23]),
    .cout(cout_30[24]),
    .sum(sum_30[24]));
  AL_FADD comp30_25 (
    .a(i30[25]),
    .b(sum_29[25]),
    .c(cout_30[24]),
    .cout(cout_30[25]),
    .sum(sum_30[25]));
  AL_FADD comp30_26 (
    .a(i30[26]),
    .b(sum_29[26]),
    .c(cout_30[25]),
    .cout(cout_30[26]),
    .sum(sum_30[26]));
  AL_FADD comp30_27 (
    .a(i30[27]),
    .b(sum_29[27]),
    .c(cout_30[26]),
    .cout(cout_30[27]),
    .sum(sum_30[27]));
  AL_FADD comp30_28 (
    .a(i30[28]),
    .b(sum_29[28]),
    .c(cout_30[27]),
    .cout(cout_30[28]),
    .sum(sum_30[28]));
  AL_FADD comp30_29 (
    .a(i30[29]),
    .b(sum_29[29]),
    .c(cout_30[28]),
    .cout(cout_30[29]),
    .sum(sum_30[29]));
  AL_FADD comp30_3 (
    .a(i30[3]),
    .b(sum_29[3]),
    .c(cout_30[2]),
    .cout(cout_30[3]),
    .sum(sum_30[3]));
  AL_FADD comp30_30 (
    .a(i30[30]),
    .b(sum_29[30]),
    .c(cout_30[29]),
    .cout(cout_30[30]),
    .sum(sum_30[30]));
  AL_FADD comp30_31 (
    .a(1'b0),
    .b(sum_29[31]),
    .c(cout_30[30]),
    .cout(cout_30[31]),
    .sum(sum_30[31]));
  AL_FADD comp30_32 (
    .a(1'b0),
    .b(sum_29[32]),
    .c(cout_30[31]),
    .cout(cout_30[32]),
    .sum(sum_30[32]));
  AL_FADD comp30_33 (
    .a(1'b0),
    .b(sum_29[33]),
    .c(cout_30[32]),
    .cout(cout_30[33]),
    .sum(sum_30[33]));
  AL_FADD comp30_34 (
    .a(1'b0),
    .b(sum_29[34]),
    .c(cout_30[33]),
    .cout(cout_30[34]),
    .sum(sum_30[34]));
  AL_FADD comp30_35 (
    .a(1'b0),
    .b(sum_29[35]),
    .c(cout_30[34]),
    .cout(cout_30[35]),
    .sum(sum_30[35]));
  AL_FADD comp30_36 (
    .a(1'b0),
    .b(sum_29[36]),
    .c(cout_30[35]),
    .cout(cout_30[36]),
    .sum(sum_30[36]));
  AL_FADD comp30_37 (
    .a(1'b0),
    .b(sum_29[37]),
    .c(cout_30[36]),
    .cout(cout_30[37]),
    .sum(sum_30[37]));
  AL_FADD comp30_38 (
    .a(1'b0),
    .b(sum_29[38]),
    .c(cout_30[37]),
    .cout(cout_30[38]),
    .sum(sum_30[38]));
  AL_FADD comp30_39 (
    .a(1'b0),
    .b(sum_29[39]),
    .c(cout_30[38]),
    .cout(cout_30[39]),
    .sum(sum_30[39]));
  AL_FADD comp30_4 (
    .a(i30[4]),
    .b(sum_29[4]),
    .c(cout_30[3]),
    .cout(cout_30[4]),
    .sum(sum_30[4]));
  AL_FADD comp30_40 (
    .a(1'b0),
    .b(sum_29[40]),
    .c(cout_30[39]),
    .cout(cout_30[40]),
    .sum(sum_30[40]));
  AL_FADD comp30_41 (
    .a(1'b0),
    .b(sum_29[41]),
    .c(cout_30[40]),
    .cout(cout_30[41]),
    .sum(sum_30[41]));
  AL_FADD comp30_42 (
    .a(1'b0),
    .b(sum_29[42]),
    .c(cout_30[41]),
    .cout(cout_30[42]),
    .sum(sum_30[42]));
  AL_FADD comp30_43 (
    .a(1'b0),
    .b(sum_29[43]),
    .c(cout_30[42]),
    .cout(cout_30[43]),
    .sum(sum_30[43]));
  AL_FADD comp30_44 (
    .a(1'b0),
    .b(sum_29[44]),
    .c(cout_30[43]),
    .cout(cout_30[44]),
    .sum(sum_30[44]));
  AL_FADD comp30_45 (
    .a(1'b0),
    .b(sum_29[45]),
    .c(cout_30[44]),
    .cout(cout_30[45]),
    .sum(sum_30[45]));
  AL_FADD comp30_46 (
    .a(1'b0),
    .b(sum_29[46]),
    .c(cout_30[45]),
    .cout(cout_30[46]),
    .sum(sum_30[46]));
  AL_FADD comp30_47 (
    .a(1'b0),
    .b(sum_29[47]),
    .c(cout_30[46]),
    .cout(cout_30[47]),
    .sum(sum_30[47]));
  AL_FADD comp30_48 (
    .a(1'b0),
    .b(sum_29[48]),
    .c(cout_30[47]),
    .cout(cout_30[48]),
    .sum(sum_30[48]));
  AL_FADD comp30_49 (
    .a(1'b0),
    .b(sum_29[49]),
    .c(cout_30[48]),
    .cout(cout_30[49]),
    .sum(sum_30[49]));
  AL_FADD comp30_5 (
    .a(i30[5]),
    .b(sum_29[5]),
    .c(cout_30[4]),
    .cout(cout_30[5]),
    .sum(sum_30[5]));
  AL_FADD comp30_50 (
    .a(1'b0),
    .b(sum_29[50]),
    .c(cout_30[49]),
    .cout(cout_30[50]),
    .sum(sum_30[50]));
  AL_FADD comp30_51 (
    .a(1'b0),
    .b(sum_29[51]),
    .c(cout_30[50]),
    .cout(cout_30[51]),
    .sum(sum_30[51]));
  AL_FADD comp30_52 (
    .a(1'b0),
    .b(sum_29[52]),
    .c(cout_30[51]),
    .cout(cout_30[52]),
    .sum(sum_30[52]));
  AL_FADD comp30_53 (
    .a(1'b0),
    .b(sum_29[53]),
    .c(cout_30[52]),
    .cout(cout_30[53]),
    .sum(sum_30[53]));
  AL_FADD comp30_54 (
    .a(1'b0),
    .b(sum_29[54]),
    .c(cout_30[53]),
    .cout(cout_30[54]),
    .sum(sum_30[54]));
  AL_FADD comp30_55 (
    .a(1'b0),
    .b(sum_29[55]),
    .c(cout_30[54]),
    .cout(cout_30[55]),
    .sum(sum_30[55]));
  AL_FADD comp30_56 (
    .a(1'b0),
    .b(sum_29[56]),
    .c(cout_30[55]),
    .cout(cout_30[56]),
    .sum(sum_30[56]));
  AL_FADD comp30_57 (
    .a(1'b0),
    .b(sum_29[57]),
    .c(cout_30[56]),
    .cout(cout_30[57]),
    .sum(sum_30[57]));
  AL_FADD comp30_58 (
    .a(1'b0),
    .b(sum_29[58]),
    .c(cout_30[57]),
    .cout(cout_30[58]),
    .sum(sum_30[58]));
  AL_FADD comp30_59 (
    .a(1'b0),
    .b(sum_29[59]),
    .c(cout_30[58]),
    .cout(cout_30[59]),
    .sum(sum_30[59]));
  AL_FADD comp30_6 (
    .a(i30[6]),
    .b(sum_29[6]),
    .c(cout_30[5]),
    .cout(cout_30[6]),
    .sum(sum_30[6]));
  AL_FADD comp30_60 (
    .a(1'b0),
    .b(sum_29[60]),
    .c(cout_30[59]),
    .cout(cout_30[60]),
    .sum(sum_30[60]));
  AL_FADD comp30_61 (
    .a(1'b0),
    .b(sum_29[61]),
    .c(cout_30[60]),
    .cout(cout_30[61]),
    .sum(sum_30[61]));
  AL_FADD comp30_62 (
    .a(1'b0),
    .b(sum_29[62]),
    .c(cout_30[61]),
    .cout(cout_30[62]),
    .sum(sum_30[62]));
  AL_FADD comp30_63 (
    .a(1'b0),
    .b(sum_29[63]),
    .c(cout_30[62]),
    .cout(cout_30[63]),
    .sum(sum_30[63]));
  AL_FADD comp30_7 (
    .a(i30[7]),
    .b(sum_29[7]),
    .c(cout_30[6]),
    .cout(cout_30[7]),
    .sum(sum_30[7]));
  AL_FADD comp30_8 (
    .a(i30[8]),
    .b(sum_29[8]),
    .c(cout_30[7]),
    .cout(cout_30[8]),
    .sum(sum_30[8]));
  AL_FADD comp30_9 (
    .a(i30[9]),
    .b(sum_29[9]),
    .c(cout_30[8]),
    .cout(cout_30[9]),
    .sum(sum_30[9]));
  AL_FADD comp31_0 (
    .a(sum_30[0]),
    .b(net_nb31_0),
    .c(1'b1),
    .cout(cout_31[0]),
    .sum(sum_31[0]));
  AL_FADD comp31_1 (
    .a(sum_30[1]),
    .b(net_nb31_1),
    .c(cout_31[0]),
    .cout(cout_31[1]),
    .sum(sum_31[1]));
  AL_FADD comp31_10 (
    .a(sum_30[10]),
    .b(net_nb31_10),
    .c(cout_31[9]),
    .cout(cout_31[10]),
    .sum(sum_31[10]));
  AL_FADD comp31_11 (
    .a(sum_30[11]),
    .b(net_nb31_11),
    .c(cout_31[10]),
    .cout(cout_31[11]),
    .sum(sum_31[11]));
  AL_FADD comp31_12 (
    .a(sum_30[12]),
    .b(net_nb31_12),
    .c(cout_31[11]),
    .cout(cout_31[12]),
    .sum(sum_31[12]));
  AL_FADD comp31_13 (
    .a(sum_30[13]),
    .b(net_nb31_13),
    .c(cout_31[12]),
    .cout(cout_31[13]),
    .sum(sum_31[13]));
  AL_FADD comp31_14 (
    .a(sum_30[14]),
    .b(net_nb31_14),
    .c(cout_31[13]),
    .cout(cout_31[14]),
    .sum(sum_31[14]));
  AL_FADD comp31_15 (
    .a(sum_30[15]),
    .b(net_nb31_15),
    .c(cout_31[14]),
    .cout(cout_31[15]),
    .sum(sum_31[15]));
  AL_FADD comp31_16 (
    .a(sum_30[16]),
    .b(net_nb31_16),
    .c(cout_31[15]),
    .cout(cout_31[16]),
    .sum(sum_31[16]));
  AL_FADD comp31_17 (
    .a(sum_30[17]),
    .b(net_nb31_17),
    .c(cout_31[16]),
    .cout(cout_31[17]),
    .sum(sum_31[17]));
  AL_FADD comp31_18 (
    .a(sum_30[18]),
    .b(net_nb31_18),
    .c(cout_31[17]),
    .cout(cout_31[18]),
    .sum(sum_31[18]));
  AL_FADD comp31_19 (
    .a(sum_30[19]),
    .b(net_nb31_19),
    .c(cout_31[18]),
    .cout(cout_31[19]),
    .sum(sum_31[19]));
  AL_FADD comp31_2 (
    .a(sum_30[2]),
    .b(net_nb31_2),
    .c(cout_31[1]),
    .cout(cout_31[2]),
    .sum(sum_31[2]));
  AL_FADD comp31_20 (
    .a(sum_30[20]),
    .b(net_nb31_20),
    .c(cout_31[19]),
    .cout(cout_31[20]),
    .sum(sum_31[20]));
  AL_FADD comp31_21 (
    .a(sum_30[21]),
    .b(net_nb31_21),
    .c(cout_31[20]),
    .cout(cout_31[21]),
    .sum(sum_31[21]));
  AL_FADD comp31_22 (
    .a(sum_30[22]),
    .b(net_nb31_22),
    .c(cout_31[21]),
    .cout(cout_31[22]),
    .sum(sum_31[22]));
  AL_FADD comp31_23 (
    .a(sum_30[23]),
    .b(net_nb31_23),
    .c(cout_31[22]),
    .cout(cout_31[23]),
    .sum(sum_31[23]));
  AL_FADD comp31_24 (
    .a(sum_30[24]),
    .b(net_nb31_24),
    .c(cout_31[23]),
    .cout(cout_31[24]),
    .sum(sum_31[24]));
  AL_FADD comp31_25 (
    .a(sum_30[25]),
    .b(net_nb31_25),
    .c(cout_31[24]),
    .cout(cout_31[25]),
    .sum(sum_31[25]));
  AL_FADD comp31_26 (
    .a(sum_30[26]),
    .b(net_nb31_26),
    .c(cout_31[25]),
    .cout(cout_31[26]),
    .sum(sum_31[26]));
  AL_FADD comp31_27 (
    .a(sum_30[27]),
    .b(net_nb31_27),
    .c(cout_31[26]),
    .cout(cout_31[27]),
    .sum(sum_31[27]));
  AL_FADD comp31_28 (
    .a(sum_30[28]),
    .b(net_nb31_28),
    .c(cout_31[27]),
    .cout(cout_31[28]),
    .sum(sum_31[28]));
  AL_FADD comp31_29 (
    .a(sum_30[29]),
    .b(net_nb31_29),
    .c(cout_31[28]),
    .cout(cout_31[29]),
    .sum(sum_31[29]));
  AL_FADD comp31_3 (
    .a(sum_30[3]),
    .b(net_nb31_3),
    .c(cout_31[2]),
    .cout(cout_31[3]),
    .sum(sum_31[3]));
  AL_FADD comp31_30 (
    .a(sum_30[30]),
    .b(net_nb31_30),
    .c(cout_31[29]),
    .cout(cout_31[30]),
    .sum(sum_31[30]));
  AL_FADD comp31_31 (
    .a(sum_30[31]),
    .b(net_nb31_31),
    .c(cout_31[30]),
    .cout(cout_31[31]),
    .sum(sum_31[31]));
  AL_FADD comp31_32 (
    .a(sum_30[32]),
    .b(net_nb31_32),
    .c(cout_31[31]),
    .cout(cout_31[32]),
    .sum(sum_31[32]));
  AL_FADD comp31_33 (
    .a(sum_30[33]),
    .b(net_nb31_33),
    .c(cout_31[32]),
    .cout(cout_31[33]),
    .sum(sum_31[33]));
  AL_FADD comp31_34 (
    .a(sum_30[34]),
    .b(net_nb31_34),
    .c(cout_31[33]),
    .cout(cout_31[34]),
    .sum(sum_31[34]));
  AL_FADD comp31_35 (
    .a(sum_30[35]),
    .b(net_nb31_35),
    .c(cout_31[34]),
    .cout(cout_31[35]),
    .sum(sum_31[35]));
  AL_FADD comp31_36 (
    .a(sum_30[36]),
    .b(net_nb31_36),
    .c(cout_31[35]),
    .cout(cout_31[36]),
    .sum(sum_31[36]));
  AL_FADD comp31_37 (
    .a(sum_30[37]),
    .b(net_nb31_37),
    .c(cout_31[36]),
    .cout(cout_31[37]),
    .sum(sum_31[37]));
  AL_FADD comp31_38 (
    .a(sum_30[38]),
    .b(net_nb31_38),
    .c(cout_31[37]),
    .cout(cout_31[38]),
    .sum(sum_31[38]));
  AL_FADD comp31_39 (
    .a(sum_30[39]),
    .b(net_nb31_39),
    .c(cout_31[38]),
    .cout(cout_31[39]),
    .sum(sum_31[39]));
  AL_FADD comp31_4 (
    .a(sum_30[4]),
    .b(net_nb31_4),
    .c(cout_31[3]),
    .cout(cout_31[4]),
    .sum(sum_31[4]));
  AL_FADD comp31_40 (
    .a(sum_30[40]),
    .b(net_nb31_40),
    .c(cout_31[39]),
    .cout(cout_31[40]),
    .sum(sum_31[40]));
  AL_FADD comp31_41 (
    .a(sum_30[41]),
    .b(net_nb31_41),
    .c(cout_31[40]),
    .cout(cout_31[41]),
    .sum(sum_31[41]));
  AL_FADD comp31_42 (
    .a(sum_30[42]),
    .b(net_nb31_42),
    .c(cout_31[41]),
    .cout(cout_31[42]),
    .sum(sum_31[42]));
  AL_FADD comp31_43 (
    .a(sum_30[43]),
    .b(net_nb31_43),
    .c(cout_31[42]),
    .cout(cout_31[43]),
    .sum(sum_31[43]));
  AL_FADD comp31_44 (
    .a(sum_30[44]),
    .b(net_nb31_44),
    .c(cout_31[43]),
    .cout(cout_31[44]),
    .sum(sum_31[44]));
  AL_FADD comp31_45 (
    .a(sum_30[45]),
    .b(net_nb31_45),
    .c(cout_31[44]),
    .cout(cout_31[45]),
    .sum(sum_31[45]));
  AL_FADD comp31_46 (
    .a(sum_30[46]),
    .b(net_nb31_46),
    .c(cout_31[45]),
    .cout(cout_31[46]),
    .sum(sum_31[46]));
  AL_FADD comp31_47 (
    .a(sum_30[47]),
    .b(net_nb31_47),
    .c(cout_31[46]),
    .cout(cout_31[47]),
    .sum(sum_31[47]));
  AL_FADD comp31_48 (
    .a(sum_30[48]),
    .b(net_nb31_48),
    .c(cout_31[47]),
    .cout(cout_31[48]),
    .sum(sum_31[48]));
  AL_FADD comp31_49 (
    .a(sum_30[49]),
    .b(net_nb31_49),
    .c(cout_31[48]),
    .cout(cout_31[49]),
    .sum(sum_31[49]));
  AL_FADD comp31_5 (
    .a(sum_30[5]),
    .b(net_nb31_5),
    .c(cout_31[4]),
    .cout(cout_31[5]),
    .sum(sum_31[5]));
  AL_FADD comp31_50 (
    .a(sum_30[50]),
    .b(net_nb31_50),
    .c(cout_31[49]),
    .cout(cout_31[50]),
    .sum(sum_31[50]));
  AL_FADD comp31_51 (
    .a(sum_30[51]),
    .b(net_nb31_51),
    .c(cout_31[50]),
    .cout(cout_31[51]),
    .sum(sum_31[51]));
  AL_FADD comp31_52 (
    .a(sum_30[52]),
    .b(net_nb31_52),
    .c(cout_31[51]),
    .cout(cout_31[52]),
    .sum(sum_31[52]));
  AL_FADD comp31_53 (
    .a(sum_30[53]),
    .b(net_nb31_53),
    .c(cout_31[52]),
    .cout(cout_31[53]),
    .sum(sum_31[53]));
  AL_FADD comp31_54 (
    .a(sum_30[54]),
    .b(net_nb31_54),
    .c(cout_31[53]),
    .cout(cout_31[54]),
    .sum(sum_31[54]));
  AL_FADD comp31_55 (
    .a(sum_30[55]),
    .b(net_nb31_55),
    .c(cout_31[54]),
    .cout(cout_31[55]),
    .sum(sum_31[55]));
  AL_FADD comp31_56 (
    .a(sum_30[56]),
    .b(net_nb31_56),
    .c(cout_31[55]),
    .cout(cout_31[56]),
    .sum(sum_31[56]));
  AL_FADD comp31_57 (
    .a(sum_30[57]),
    .b(net_nb31_57),
    .c(cout_31[56]),
    .cout(cout_31[57]),
    .sum(sum_31[57]));
  AL_FADD comp31_58 (
    .a(sum_30[58]),
    .b(net_nb31_58),
    .c(cout_31[57]),
    .cout(cout_31[58]),
    .sum(sum_31[58]));
  AL_FADD comp31_59 (
    .a(sum_30[59]),
    .b(net_nb31_59),
    .c(cout_31[58]),
    .cout(cout_31[59]),
    .sum(sum_31[59]));
  AL_FADD comp31_6 (
    .a(sum_30[6]),
    .b(net_nb31_6),
    .c(cout_31[5]),
    .cout(cout_31[6]),
    .sum(sum_31[6]));
  AL_FADD comp31_60 (
    .a(sum_30[60]),
    .b(net_nb31_60),
    .c(cout_31[59]),
    .cout(cout_31[60]),
    .sum(sum_31[60]));
  AL_FADD comp31_61 (
    .a(sum_30[61]),
    .b(net_nb31_61),
    .c(cout_31[60]),
    .cout(cout_31[61]),
    .sum(sum_31[61]));
  AL_FADD comp31_62 (
    .a(sum_30[62]),
    .b(net_nb31_62),
    .c(cout_31[61]),
    .cout(cout_31[62]),
    .sum(sum_31[62]));
  AL_FADD comp31_63 (
    .a(sum_30[63]),
    .b(net_nb31_63),
    .c(cout_31[62]),
    .cout(cout_31[63]),
    .sum(sum_31[63]));
  AL_FADD comp31_7 (
    .a(sum_30[7]),
    .b(net_nb31_7),
    .c(cout_31[6]),
    .cout(cout_31[7]),
    .sum(sum_31[7]));
  AL_FADD comp31_8 (
    .a(sum_30[8]),
    .b(net_nb31_8),
    .c(cout_31[7]),
    .cout(cout_31[8]),
    .sum(sum_31[8]));
  AL_FADD comp31_9 (
    .a(sum_30[9]),
    .b(net_nb31_9),
    .c(cout_31[8]),
    .cout(cout_31[9]),
    .sum(sum_31[9]));
  AL_FADD comp32_0 (
    .a(sum_31[0]),
    .b(net_nb32_0),
    .c(1'b1),
    .cout(cout_32[0]),
    .sum(sum_32[0]));
  AL_FADD comp32_1 (
    .a(sum_31[1]),
    .b(net_nb32_1),
    .c(cout_32[0]),
    .cout(cout_32[1]),
    .sum(sum_32[1]));
  AL_FADD comp32_10 (
    .a(sum_31[10]),
    .b(net_nb32_10),
    .c(cout_32[9]),
    .cout(cout_32[10]),
    .sum(sum_32[10]));
  AL_FADD comp32_11 (
    .a(sum_31[11]),
    .b(net_nb32_11),
    .c(cout_32[10]),
    .cout(cout_32[11]),
    .sum(sum_32[11]));
  AL_FADD comp32_12 (
    .a(sum_31[12]),
    .b(net_nb32_12),
    .c(cout_32[11]),
    .cout(cout_32[12]),
    .sum(sum_32[12]));
  AL_FADD comp32_13 (
    .a(sum_31[13]),
    .b(net_nb32_13),
    .c(cout_32[12]),
    .cout(cout_32[13]),
    .sum(sum_32[13]));
  AL_FADD comp32_14 (
    .a(sum_31[14]),
    .b(net_nb32_14),
    .c(cout_32[13]),
    .cout(cout_32[14]),
    .sum(sum_32[14]));
  AL_FADD comp32_15 (
    .a(sum_31[15]),
    .b(net_nb32_15),
    .c(cout_32[14]),
    .cout(cout_32[15]),
    .sum(sum_32[15]));
  AL_FADD comp32_16 (
    .a(sum_31[16]),
    .b(net_nb32_16),
    .c(cout_32[15]),
    .cout(cout_32[16]),
    .sum(sum_32[16]));
  AL_FADD comp32_17 (
    .a(sum_31[17]),
    .b(net_nb32_17),
    .c(cout_32[16]),
    .cout(cout_32[17]),
    .sum(sum_32[17]));
  AL_FADD comp32_18 (
    .a(sum_31[18]),
    .b(net_nb32_18),
    .c(cout_32[17]),
    .cout(cout_32[18]),
    .sum(sum_32[18]));
  AL_FADD comp32_19 (
    .a(sum_31[19]),
    .b(net_nb32_19),
    .c(cout_32[18]),
    .cout(cout_32[19]),
    .sum(sum_32[19]));
  AL_FADD comp32_2 (
    .a(sum_31[2]),
    .b(net_nb32_2),
    .c(cout_32[1]),
    .cout(cout_32[2]),
    .sum(sum_32[2]));
  AL_FADD comp32_20 (
    .a(sum_31[20]),
    .b(net_nb32_20),
    .c(cout_32[19]),
    .cout(cout_32[20]),
    .sum(sum_32[20]));
  AL_FADD comp32_21 (
    .a(sum_31[21]),
    .b(net_nb32_21),
    .c(cout_32[20]),
    .cout(cout_32[21]),
    .sum(sum_32[21]));
  AL_FADD comp32_22 (
    .a(sum_31[22]),
    .b(net_nb32_22),
    .c(cout_32[21]),
    .cout(cout_32[22]),
    .sum(sum_32[22]));
  AL_FADD comp32_23 (
    .a(sum_31[23]),
    .b(net_nb32_23),
    .c(cout_32[22]),
    .cout(cout_32[23]),
    .sum(sum_32[23]));
  AL_FADD comp32_24 (
    .a(sum_31[24]),
    .b(net_nb32_24),
    .c(cout_32[23]),
    .cout(cout_32[24]),
    .sum(sum_32[24]));
  AL_FADD comp32_25 (
    .a(sum_31[25]),
    .b(net_nb32_25),
    .c(cout_32[24]),
    .cout(cout_32[25]),
    .sum(sum_32[25]));
  AL_FADD comp32_26 (
    .a(sum_31[26]),
    .b(net_nb32_26),
    .c(cout_32[25]),
    .cout(cout_32[26]),
    .sum(sum_32[26]));
  AL_FADD comp32_27 (
    .a(sum_31[27]),
    .b(net_nb32_27),
    .c(cout_32[26]),
    .cout(cout_32[27]),
    .sum(sum_32[27]));
  AL_FADD comp32_28 (
    .a(sum_31[28]),
    .b(net_nb32_28),
    .c(cout_32[27]),
    .cout(cout_32[28]),
    .sum(sum_32[28]));
  AL_FADD comp32_29 (
    .a(sum_31[29]),
    .b(net_nb32_29),
    .c(cout_32[28]),
    .cout(cout_32[29]),
    .sum(sum_32[29]));
  AL_FADD comp32_3 (
    .a(sum_31[3]),
    .b(net_nb32_3),
    .c(cout_32[2]),
    .cout(cout_32[3]),
    .sum(sum_32[3]));
  AL_FADD comp32_30 (
    .a(sum_31[30]),
    .b(net_nb32_30),
    .c(cout_32[29]),
    .cout(cout_32[30]),
    .sum(sum_32[30]));
  AL_FADD comp32_31 (
    .a(sum_31[31]),
    .b(net_nb32_31),
    .c(cout_32[30]),
    .cout(cout_32[31]),
    .sum(sum_32[31]));
  AL_FADD comp32_32 (
    .a(sum_31[32]),
    .b(net_nb32_32),
    .c(cout_32[31]),
    .cout(cout_32[32]),
    .sum(sum_32[32]));
  AL_FADD comp32_33 (
    .a(sum_31[33]),
    .b(net_nb32_33),
    .c(cout_32[32]),
    .cout(cout_32[33]),
    .sum(sum_32[33]));
  AL_FADD comp32_34 (
    .a(sum_31[34]),
    .b(net_nb32_34),
    .c(cout_32[33]),
    .cout(cout_32[34]),
    .sum(sum_32[34]));
  AL_FADD comp32_35 (
    .a(sum_31[35]),
    .b(net_nb32_35),
    .c(cout_32[34]),
    .cout(cout_32[35]),
    .sum(sum_32[35]));
  AL_FADD comp32_36 (
    .a(sum_31[36]),
    .b(net_nb32_36),
    .c(cout_32[35]),
    .cout(cout_32[36]),
    .sum(sum_32[36]));
  AL_FADD comp32_37 (
    .a(sum_31[37]),
    .b(net_nb32_37),
    .c(cout_32[36]),
    .cout(cout_32[37]),
    .sum(sum_32[37]));
  AL_FADD comp32_38 (
    .a(sum_31[38]),
    .b(net_nb32_38),
    .c(cout_32[37]),
    .cout(cout_32[38]),
    .sum(sum_32[38]));
  AL_FADD comp32_39 (
    .a(sum_31[39]),
    .b(net_nb32_39),
    .c(cout_32[38]),
    .cout(cout_32[39]),
    .sum(sum_32[39]));
  AL_FADD comp32_4 (
    .a(sum_31[4]),
    .b(net_nb32_4),
    .c(cout_32[3]),
    .cout(cout_32[4]),
    .sum(sum_32[4]));
  AL_FADD comp32_40 (
    .a(sum_31[40]),
    .b(net_nb32_40),
    .c(cout_32[39]),
    .cout(cout_32[40]),
    .sum(sum_32[40]));
  AL_FADD comp32_41 (
    .a(sum_31[41]),
    .b(net_nb32_41),
    .c(cout_32[40]),
    .cout(cout_32[41]),
    .sum(sum_32[41]));
  AL_FADD comp32_42 (
    .a(sum_31[42]),
    .b(net_nb32_42),
    .c(cout_32[41]),
    .cout(cout_32[42]),
    .sum(sum_32[42]));
  AL_FADD comp32_43 (
    .a(sum_31[43]),
    .b(net_nb32_43),
    .c(cout_32[42]),
    .cout(cout_32[43]),
    .sum(sum_32[43]));
  AL_FADD comp32_44 (
    .a(sum_31[44]),
    .b(net_nb32_44),
    .c(cout_32[43]),
    .cout(cout_32[44]),
    .sum(sum_32[44]));
  AL_FADD comp32_45 (
    .a(sum_31[45]),
    .b(net_nb32_45),
    .c(cout_32[44]),
    .cout(cout_32[45]),
    .sum(sum_32[45]));
  AL_FADD comp32_46 (
    .a(sum_31[46]),
    .b(net_nb32_46),
    .c(cout_32[45]),
    .cout(cout_32[46]),
    .sum(sum_32[46]));
  AL_FADD comp32_47 (
    .a(sum_31[47]),
    .b(net_nb32_47),
    .c(cout_32[46]),
    .cout(cout_32[47]),
    .sum(sum_32[47]));
  AL_FADD comp32_48 (
    .a(sum_31[48]),
    .b(net_nb32_48),
    .c(cout_32[47]),
    .cout(cout_32[48]),
    .sum(sum_32[48]));
  AL_FADD comp32_49 (
    .a(sum_31[49]),
    .b(net_nb32_49),
    .c(cout_32[48]),
    .cout(cout_32[49]),
    .sum(sum_32[49]));
  AL_FADD comp32_5 (
    .a(sum_31[5]),
    .b(net_nb32_5),
    .c(cout_32[4]),
    .cout(cout_32[5]),
    .sum(sum_32[5]));
  AL_FADD comp32_50 (
    .a(sum_31[50]),
    .b(net_nb32_50),
    .c(cout_32[49]),
    .cout(cout_32[50]),
    .sum(sum_32[50]));
  AL_FADD comp32_51 (
    .a(sum_31[51]),
    .b(net_nb32_51),
    .c(cout_32[50]),
    .cout(cout_32[51]),
    .sum(sum_32[51]));
  AL_FADD comp32_52 (
    .a(sum_31[52]),
    .b(net_nb32_52),
    .c(cout_32[51]),
    .cout(cout_32[52]),
    .sum(sum_32[52]));
  AL_FADD comp32_53 (
    .a(sum_31[53]),
    .b(net_nb32_53),
    .c(cout_32[52]),
    .cout(cout_32[53]),
    .sum(sum_32[53]));
  AL_FADD comp32_54 (
    .a(sum_31[54]),
    .b(net_nb32_54),
    .c(cout_32[53]),
    .cout(cout_32[54]),
    .sum(sum_32[54]));
  AL_FADD comp32_55 (
    .a(sum_31[55]),
    .b(net_nb32_55),
    .c(cout_32[54]),
    .cout(cout_32[55]),
    .sum(sum_32[55]));
  AL_FADD comp32_56 (
    .a(sum_31[56]),
    .b(net_nb32_56),
    .c(cout_32[55]),
    .cout(cout_32[56]),
    .sum(sum_32[56]));
  AL_FADD comp32_57 (
    .a(sum_31[57]),
    .b(net_nb32_57),
    .c(cout_32[56]),
    .cout(cout_32[57]),
    .sum(sum_32[57]));
  AL_FADD comp32_58 (
    .a(sum_31[58]),
    .b(net_nb32_58),
    .c(cout_32[57]),
    .cout(cout_32[58]),
    .sum(sum_32[58]));
  AL_FADD comp32_59 (
    .a(sum_31[59]),
    .b(net_nb32_59),
    .c(cout_32[58]),
    .cout(cout_32[59]),
    .sum(sum_32[59]));
  AL_FADD comp32_6 (
    .a(sum_31[6]),
    .b(net_nb32_6),
    .c(cout_32[5]),
    .cout(cout_32[6]),
    .sum(sum_32[6]));
  AL_FADD comp32_60 (
    .a(sum_31[60]),
    .b(net_nb32_60),
    .c(cout_32[59]),
    .cout(cout_32[60]),
    .sum(sum_32[60]));
  AL_FADD comp32_61 (
    .a(sum_31[61]),
    .b(net_nb32_61),
    .c(cout_32[60]),
    .cout(cout_32[61]),
    .sum(sum_32[61]));
  AL_FADD comp32_62 (
    .a(sum_31[62]),
    .b(net_nb32_62),
    .c(cout_32[61]),
    .cout(cout_32[62]),
    .sum(sum_32[62]));
  AL_FADD comp32_63 (
    .a(sum_31[63]),
    .b(net_nb32_63),
    .c(cout_32[62]),
    .cout(cout_32[63]),
    .sum(sum_32[63]));
  AL_FADD comp32_7 (
    .a(sum_31[7]),
    .b(net_nb32_7),
    .c(cout_32[6]),
    .cout(cout_32[7]),
    .sum(sum_32[7]));
  AL_FADD comp32_8 (
    .a(sum_31[8]),
    .b(net_nb32_8),
    .c(cout_32[7]),
    .cout(cout_32[8]),
    .sum(sum_32[8]));
  AL_FADD comp32_9 (
    .a(sum_31[9]),
    .b(net_nb32_9),
    .c(cout_32[8]),
    .cout(cout_32[9]),
    .sum(sum_32[9]));
  AL_FADD comp3_0 (
    .a(i3[0]),
    .b(sum_2[0]),
    .c(1'b0),
    .cout(cout_3[0]),
    .sum(sum_3[0]));
  AL_FADD comp3_1 (
    .a(i3[1]),
    .b(sum_2[1]),
    .c(cout_3[0]),
    .cout(cout_3[1]),
    .sum(sum_3[1]));
  AL_FADD comp3_10 (
    .a(i3[10]),
    .b(sum_2[10]),
    .c(cout_3[9]),
    .cout(cout_3[10]),
    .sum(sum_3[10]));
  AL_FADD comp3_11 (
    .a(i3[11]),
    .b(sum_2[11]),
    .c(cout_3[10]),
    .cout(cout_3[11]),
    .sum(sum_3[11]));
  AL_FADD comp3_12 (
    .a(i3[12]),
    .b(sum_2[12]),
    .c(cout_3[11]),
    .cout(cout_3[12]),
    .sum(sum_3[12]));
  AL_FADD comp3_13 (
    .a(i3[13]),
    .b(sum_2[13]),
    .c(cout_3[12]),
    .cout(cout_3[13]),
    .sum(sum_3[13]));
  AL_FADD comp3_14 (
    .a(i3[14]),
    .b(sum_2[14]),
    .c(cout_3[13]),
    .cout(cout_3[14]),
    .sum(sum_3[14]));
  AL_FADD comp3_15 (
    .a(i3[15]),
    .b(sum_2[15]),
    .c(cout_3[14]),
    .cout(cout_3[15]),
    .sum(sum_3[15]));
  AL_FADD comp3_16 (
    .a(i3[16]),
    .b(sum_2[16]),
    .c(cout_3[15]),
    .cout(cout_3[16]),
    .sum(sum_3[16]));
  AL_FADD comp3_17 (
    .a(i3[17]),
    .b(sum_2[17]),
    .c(cout_3[16]),
    .cout(cout_3[17]),
    .sum(sum_3[17]));
  AL_FADD comp3_18 (
    .a(i3[18]),
    .b(sum_2[18]),
    .c(cout_3[17]),
    .cout(cout_3[18]),
    .sum(sum_3[18]));
  AL_FADD comp3_19 (
    .a(i3[19]),
    .b(sum_2[19]),
    .c(cout_3[18]),
    .cout(cout_3[19]),
    .sum(sum_3[19]));
  AL_FADD comp3_2 (
    .a(i3[2]),
    .b(sum_2[2]),
    .c(cout_3[1]),
    .cout(cout_3[2]),
    .sum(sum_3[2]));
  AL_FADD comp3_20 (
    .a(i3[20]),
    .b(sum_2[20]),
    .c(cout_3[19]),
    .cout(cout_3[20]),
    .sum(sum_3[20]));
  AL_FADD comp3_21 (
    .a(i3[21]),
    .b(sum_2[21]),
    .c(cout_3[20]),
    .cout(cout_3[21]),
    .sum(sum_3[21]));
  AL_FADD comp3_22 (
    .a(i3[22]),
    .b(sum_2[22]),
    .c(cout_3[21]),
    .cout(cout_3[22]),
    .sum(sum_3[22]));
  AL_FADD comp3_23 (
    .a(i3[23]),
    .b(sum_2[23]),
    .c(cout_3[22]),
    .cout(cout_3[23]),
    .sum(sum_3[23]));
  AL_FADD comp3_24 (
    .a(i3[24]),
    .b(sum_2[24]),
    .c(cout_3[23]),
    .cout(cout_3[24]),
    .sum(sum_3[24]));
  AL_FADD comp3_25 (
    .a(i3[25]),
    .b(sum_2[25]),
    .c(cout_3[24]),
    .cout(cout_3[25]),
    .sum(sum_3[25]));
  AL_FADD comp3_26 (
    .a(i3[26]),
    .b(sum_2[26]),
    .c(cout_3[25]),
    .cout(cout_3[26]),
    .sum(sum_3[26]));
  AL_FADD comp3_27 (
    .a(i3[27]),
    .b(sum_2[27]),
    .c(cout_3[26]),
    .cout(cout_3[27]),
    .sum(sum_3[27]));
  AL_FADD comp3_28 (
    .a(i3[28]),
    .b(sum_2[28]),
    .c(cout_3[27]),
    .cout(cout_3[28]),
    .sum(sum_3[28]));
  AL_FADD comp3_29 (
    .a(i3[29]),
    .b(sum_2[29]),
    .c(cout_3[28]),
    .cout(cout_3[29]),
    .sum(sum_3[29]));
  AL_FADD comp3_3 (
    .a(i3[3]),
    .b(sum_2[3]),
    .c(cout_3[2]),
    .cout(cout_3[3]),
    .sum(sum_3[3]));
  AL_FADD comp3_30 (
    .a(i3[30]),
    .b(sum_2[30]),
    .c(cout_3[29]),
    .cout(cout_3[30]),
    .sum(sum_3[30]));
  AL_FADD comp3_31 (
    .a(i3[31]),
    .b(sum_2[31]),
    .c(cout_3[30]),
    .cout(cout_3[31]),
    .sum(sum_3[31]));
  AL_FADD comp3_32 (
    .a(i3[32]),
    .b(sum_2[32]),
    .c(cout_3[31]),
    .cout(cout_3[32]),
    .sum(sum_3[32]));
  AL_FADD comp3_33 (
    .a(i3[33]),
    .b(sum_2[33]),
    .c(cout_3[32]),
    .cout(cout_3[33]),
    .sum(sum_3[33]));
  AL_FADD comp3_34 (
    .a(i3[34]),
    .b(sum_2[34]),
    .c(cout_3[33]),
    .cout(cout_3[34]),
    .sum(sum_3[34]));
  AL_FADD comp3_35 (
    .a(i3[35]),
    .b(sum_2[35]),
    .c(cout_3[34]),
    .cout(cout_3[35]),
    .sum(sum_3[35]));
  AL_FADD comp3_36 (
    .a(i3[36]),
    .b(sum_2[36]),
    .c(cout_3[35]),
    .cout(cout_3[36]),
    .sum(sum_3[36]));
  AL_FADD comp3_37 (
    .a(i3[37]),
    .b(sum_2[37]),
    .c(cout_3[36]),
    .cout(cout_3[37]),
    .sum(sum_3[37]));
  AL_FADD comp3_38 (
    .a(i3[38]),
    .b(sum_2[38]),
    .c(cout_3[37]),
    .cout(cout_3[38]),
    .sum(sum_3[38]));
  AL_FADD comp3_39 (
    .a(i3[39]),
    .b(sum_2[39]),
    .c(cout_3[38]),
    .cout(cout_3[39]),
    .sum(sum_3[39]));
  AL_FADD comp3_4 (
    .a(i3[4]),
    .b(sum_2[4]),
    .c(cout_3[3]),
    .cout(cout_3[4]),
    .sum(sum_3[4]));
  AL_FADD comp3_40 (
    .a(i3[40]),
    .b(sum_2[40]),
    .c(cout_3[39]),
    .cout(cout_3[40]),
    .sum(sum_3[40]));
  AL_FADD comp3_41 (
    .a(i3[41]),
    .b(sum_2[41]),
    .c(cout_3[40]),
    .cout(cout_3[41]),
    .sum(sum_3[41]));
  AL_FADD comp3_42 (
    .a(i3[42]),
    .b(sum_2[42]),
    .c(cout_3[41]),
    .cout(cout_3[42]),
    .sum(sum_3[42]));
  AL_FADD comp3_43 (
    .a(i3[43]),
    .b(sum_2[43]),
    .c(cout_3[42]),
    .cout(cout_3[43]),
    .sum(sum_3[43]));
  AL_FADD comp3_44 (
    .a(i3[44]),
    .b(sum_2[44]),
    .c(cout_3[43]),
    .cout(cout_3[44]),
    .sum(sum_3[44]));
  AL_FADD comp3_45 (
    .a(i3[45]),
    .b(sum_2[45]),
    .c(cout_3[44]),
    .cout(cout_3[45]),
    .sum(sum_3[45]));
  AL_FADD comp3_46 (
    .a(i3[46]),
    .b(sum_2[46]),
    .c(cout_3[45]),
    .cout(cout_3[46]),
    .sum(sum_3[46]));
  AL_FADD comp3_47 (
    .a(i3[47]),
    .b(sum_2[47]),
    .c(cout_3[46]),
    .cout(cout_3[47]),
    .sum(sum_3[47]));
  AL_FADD comp3_48 (
    .a(i3[48]),
    .b(sum_2[48]),
    .c(cout_3[47]),
    .cout(cout_3[48]),
    .sum(sum_3[48]));
  AL_FADD comp3_49 (
    .a(i3[49]),
    .b(sum_2[49]),
    .c(cout_3[48]),
    .cout(cout_3[49]),
    .sum(sum_3[49]));
  AL_FADD comp3_5 (
    .a(i3[5]),
    .b(sum_2[5]),
    .c(cout_3[4]),
    .cout(cout_3[5]),
    .sum(sum_3[5]));
  AL_FADD comp3_50 (
    .a(i3[50]),
    .b(sum_2[50]),
    .c(cout_3[49]),
    .cout(cout_3[50]),
    .sum(sum_3[50]));
  AL_FADD comp3_51 (
    .a(i3[51]),
    .b(sum_2[51]),
    .c(cout_3[50]),
    .cout(cout_3[51]),
    .sum(sum_3[51]));
  AL_FADD comp3_52 (
    .a(i3[52]),
    .b(sum_2[52]),
    .c(cout_3[51]),
    .cout(cout_3[52]),
    .sum(sum_3[52]));
  AL_FADD comp3_53 (
    .a(i3[53]),
    .b(sum_2[53]),
    .c(cout_3[52]),
    .cout(cout_3[53]),
    .sum(sum_3[53]));
  AL_FADD comp3_54 (
    .a(i3[54]),
    .b(sum_2[54]),
    .c(cout_3[53]),
    .cout(cout_3[54]),
    .sum(sum_3[54]));
  AL_FADD comp3_55 (
    .a(i3[55]),
    .b(sum_2[55]),
    .c(cout_3[54]),
    .cout(cout_3[55]),
    .sum(sum_3[55]));
  AL_FADD comp3_56 (
    .a(i3[56]),
    .b(sum_2[56]),
    .c(cout_3[55]),
    .cout(cout_3[56]),
    .sum(sum_3[56]));
  AL_FADD comp3_57 (
    .a(i3[57]),
    .b(sum_2[57]),
    .c(cout_3[56]),
    .cout(cout_3[57]),
    .sum(sum_3[57]));
  AL_FADD comp3_58 (
    .a(1'b0),
    .b(sum_2[58]),
    .c(cout_3[57]),
    .cout(cout_3[58]),
    .sum(sum_3[58]));
  AL_FADD comp3_59 (
    .a(1'b0),
    .b(sum_2[59]),
    .c(cout_3[58]),
    .cout(cout_3[59]),
    .sum(sum_3[59]));
  AL_FADD comp3_6 (
    .a(i3[6]),
    .b(sum_2[6]),
    .c(cout_3[5]),
    .cout(cout_3[6]),
    .sum(sum_3[6]));
  AL_FADD comp3_60 (
    .a(1'b0),
    .b(sum_2[60]),
    .c(cout_3[59]),
    .cout(cout_3[60]),
    .sum(sum_3[60]));
  AL_FADD comp3_61 (
    .a(1'b0),
    .b(sum_2[61]),
    .c(cout_3[60]),
    .cout(cout_3[61]),
    .sum(sum_3[61]));
  AL_FADD comp3_62 (
    .a(1'b0),
    .b(sum_2[62]),
    .c(cout_3[61]),
    .cout(cout_3[62]),
    .sum(sum_3[62]));
  AL_FADD comp3_63 (
    .a(1'b0),
    .b(sum_2[63]),
    .c(cout_3[62]),
    .cout(cout_3[63]),
    .sum(sum_3[63]));
  AL_FADD comp3_7 (
    .a(i3[7]),
    .b(sum_2[7]),
    .c(cout_3[6]),
    .cout(cout_3[7]),
    .sum(sum_3[7]));
  AL_FADD comp3_8 (
    .a(i3[8]),
    .b(sum_2[8]),
    .c(cout_3[7]),
    .cout(cout_3[8]),
    .sum(sum_3[8]));
  AL_FADD comp3_9 (
    .a(i3[9]),
    .b(sum_2[9]),
    .c(cout_3[8]),
    .cout(cout_3[9]),
    .sum(sum_3[9]));
  AL_FADD comp4_0 (
    .a(i4[0]),
    .b(sum_3[0]),
    .c(1'b0),
    .cout(cout_4[0]),
    .sum(sum_4[0]));
  AL_FADD comp4_1 (
    .a(i4[1]),
    .b(sum_3[1]),
    .c(cout_4[0]),
    .cout(cout_4[1]),
    .sum(sum_4[1]));
  AL_FADD comp4_10 (
    .a(i4[10]),
    .b(sum_3[10]),
    .c(cout_4[9]),
    .cout(cout_4[10]),
    .sum(sum_4[10]));
  AL_FADD comp4_11 (
    .a(i4[11]),
    .b(sum_3[11]),
    .c(cout_4[10]),
    .cout(cout_4[11]),
    .sum(sum_4[11]));
  AL_FADD comp4_12 (
    .a(i4[12]),
    .b(sum_3[12]),
    .c(cout_4[11]),
    .cout(cout_4[12]),
    .sum(sum_4[12]));
  AL_FADD comp4_13 (
    .a(i4[13]),
    .b(sum_3[13]),
    .c(cout_4[12]),
    .cout(cout_4[13]),
    .sum(sum_4[13]));
  AL_FADD comp4_14 (
    .a(i4[14]),
    .b(sum_3[14]),
    .c(cout_4[13]),
    .cout(cout_4[14]),
    .sum(sum_4[14]));
  AL_FADD comp4_15 (
    .a(i4[15]),
    .b(sum_3[15]),
    .c(cout_4[14]),
    .cout(cout_4[15]),
    .sum(sum_4[15]));
  AL_FADD comp4_16 (
    .a(i4[16]),
    .b(sum_3[16]),
    .c(cout_4[15]),
    .cout(cout_4[16]),
    .sum(sum_4[16]));
  AL_FADD comp4_17 (
    .a(i4[17]),
    .b(sum_3[17]),
    .c(cout_4[16]),
    .cout(cout_4[17]),
    .sum(sum_4[17]));
  AL_FADD comp4_18 (
    .a(i4[18]),
    .b(sum_3[18]),
    .c(cout_4[17]),
    .cout(cout_4[18]),
    .sum(sum_4[18]));
  AL_FADD comp4_19 (
    .a(i4[19]),
    .b(sum_3[19]),
    .c(cout_4[18]),
    .cout(cout_4[19]),
    .sum(sum_4[19]));
  AL_FADD comp4_2 (
    .a(i4[2]),
    .b(sum_3[2]),
    .c(cout_4[1]),
    .cout(cout_4[2]),
    .sum(sum_4[2]));
  AL_FADD comp4_20 (
    .a(i4[20]),
    .b(sum_3[20]),
    .c(cout_4[19]),
    .cout(cout_4[20]),
    .sum(sum_4[20]));
  AL_FADD comp4_21 (
    .a(i4[21]),
    .b(sum_3[21]),
    .c(cout_4[20]),
    .cout(cout_4[21]),
    .sum(sum_4[21]));
  AL_FADD comp4_22 (
    .a(i4[22]),
    .b(sum_3[22]),
    .c(cout_4[21]),
    .cout(cout_4[22]),
    .sum(sum_4[22]));
  AL_FADD comp4_23 (
    .a(i4[23]),
    .b(sum_3[23]),
    .c(cout_4[22]),
    .cout(cout_4[23]),
    .sum(sum_4[23]));
  AL_FADD comp4_24 (
    .a(i4[24]),
    .b(sum_3[24]),
    .c(cout_4[23]),
    .cout(cout_4[24]),
    .sum(sum_4[24]));
  AL_FADD comp4_25 (
    .a(i4[25]),
    .b(sum_3[25]),
    .c(cout_4[24]),
    .cout(cout_4[25]),
    .sum(sum_4[25]));
  AL_FADD comp4_26 (
    .a(i4[26]),
    .b(sum_3[26]),
    .c(cout_4[25]),
    .cout(cout_4[26]),
    .sum(sum_4[26]));
  AL_FADD comp4_27 (
    .a(i4[27]),
    .b(sum_3[27]),
    .c(cout_4[26]),
    .cout(cout_4[27]),
    .sum(sum_4[27]));
  AL_FADD comp4_28 (
    .a(i4[28]),
    .b(sum_3[28]),
    .c(cout_4[27]),
    .cout(cout_4[28]),
    .sum(sum_4[28]));
  AL_FADD comp4_29 (
    .a(i4[29]),
    .b(sum_3[29]),
    .c(cout_4[28]),
    .cout(cout_4[29]),
    .sum(sum_4[29]));
  AL_FADD comp4_3 (
    .a(i4[3]),
    .b(sum_3[3]),
    .c(cout_4[2]),
    .cout(cout_4[3]),
    .sum(sum_4[3]));
  AL_FADD comp4_30 (
    .a(i4[30]),
    .b(sum_3[30]),
    .c(cout_4[29]),
    .cout(cout_4[30]),
    .sum(sum_4[30]));
  AL_FADD comp4_31 (
    .a(i4[31]),
    .b(sum_3[31]),
    .c(cout_4[30]),
    .cout(cout_4[31]),
    .sum(sum_4[31]));
  AL_FADD comp4_32 (
    .a(i4[32]),
    .b(sum_3[32]),
    .c(cout_4[31]),
    .cout(cout_4[32]),
    .sum(sum_4[32]));
  AL_FADD comp4_33 (
    .a(i4[33]),
    .b(sum_3[33]),
    .c(cout_4[32]),
    .cout(cout_4[33]),
    .sum(sum_4[33]));
  AL_FADD comp4_34 (
    .a(i4[34]),
    .b(sum_3[34]),
    .c(cout_4[33]),
    .cout(cout_4[34]),
    .sum(sum_4[34]));
  AL_FADD comp4_35 (
    .a(i4[35]),
    .b(sum_3[35]),
    .c(cout_4[34]),
    .cout(cout_4[35]),
    .sum(sum_4[35]));
  AL_FADD comp4_36 (
    .a(i4[36]),
    .b(sum_3[36]),
    .c(cout_4[35]),
    .cout(cout_4[36]),
    .sum(sum_4[36]));
  AL_FADD comp4_37 (
    .a(i4[37]),
    .b(sum_3[37]),
    .c(cout_4[36]),
    .cout(cout_4[37]),
    .sum(sum_4[37]));
  AL_FADD comp4_38 (
    .a(i4[38]),
    .b(sum_3[38]),
    .c(cout_4[37]),
    .cout(cout_4[38]),
    .sum(sum_4[38]));
  AL_FADD comp4_39 (
    .a(i4[39]),
    .b(sum_3[39]),
    .c(cout_4[38]),
    .cout(cout_4[39]),
    .sum(sum_4[39]));
  AL_FADD comp4_4 (
    .a(i4[4]),
    .b(sum_3[4]),
    .c(cout_4[3]),
    .cout(cout_4[4]),
    .sum(sum_4[4]));
  AL_FADD comp4_40 (
    .a(i4[40]),
    .b(sum_3[40]),
    .c(cout_4[39]),
    .cout(cout_4[40]),
    .sum(sum_4[40]));
  AL_FADD comp4_41 (
    .a(i4[41]),
    .b(sum_3[41]),
    .c(cout_4[40]),
    .cout(cout_4[41]),
    .sum(sum_4[41]));
  AL_FADD comp4_42 (
    .a(i4[42]),
    .b(sum_3[42]),
    .c(cout_4[41]),
    .cout(cout_4[42]),
    .sum(sum_4[42]));
  AL_FADD comp4_43 (
    .a(i4[43]),
    .b(sum_3[43]),
    .c(cout_4[42]),
    .cout(cout_4[43]),
    .sum(sum_4[43]));
  AL_FADD comp4_44 (
    .a(i4[44]),
    .b(sum_3[44]),
    .c(cout_4[43]),
    .cout(cout_4[44]),
    .sum(sum_4[44]));
  AL_FADD comp4_45 (
    .a(i4[45]),
    .b(sum_3[45]),
    .c(cout_4[44]),
    .cout(cout_4[45]),
    .sum(sum_4[45]));
  AL_FADD comp4_46 (
    .a(i4[46]),
    .b(sum_3[46]),
    .c(cout_4[45]),
    .cout(cout_4[46]),
    .sum(sum_4[46]));
  AL_FADD comp4_47 (
    .a(i4[47]),
    .b(sum_3[47]),
    .c(cout_4[46]),
    .cout(cout_4[47]),
    .sum(sum_4[47]));
  AL_FADD comp4_48 (
    .a(i4[48]),
    .b(sum_3[48]),
    .c(cout_4[47]),
    .cout(cout_4[48]),
    .sum(sum_4[48]));
  AL_FADD comp4_49 (
    .a(i4[49]),
    .b(sum_3[49]),
    .c(cout_4[48]),
    .cout(cout_4[49]),
    .sum(sum_4[49]));
  AL_FADD comp4_5 (
    .a(i4[5]),
    .b(sum_3[5]),
    .c(cout_4[4]),
    .cout(cout_4[5]),
    .sum(sum_4[5]));
  AL_FADD comp4_50 (
    .a(i4[50]),
    .b(sum_3[50]),
    .c(cout_4[49]),
    .cout(cout_4[50]),
    .sum(sum_4[50]));
  AL_FADD comp4_51 (
    .a(i4[51]),
    .b(sum_3[51]),
    .c(cout_4[50]),
    .cout(cout_4[51]),
    .sum(sum_4[51]));
  AL_FADD comp4_52 (
    .a(i4[52]),
    .b(sum_3[52]),
    .c(cout_4[51]),
    .cout(cout_4[52]),
    .sum(sum_4[52]));
  AL_FADD comp4_53 (
    .a(i4[53]),
    .b(sum_3[53]),
    .c(cout_4[52]),
    .cout(cout_4[53]),
    .sum(sum_4[53]));
  AL_FADD comp4_54 (
    .a(i4[54]),
    .b(sum_3[54]),
    .c(cout_4[53]),
    .cout(cout_4[54]),
    .sum(sum_4[54]));
  AL_FADD comp4_55 (
    .a(i4[55]),
    .b(sum_3[55]),
    .c(cout_4[54]),
    .cout(cout_4[55]),
    .sum(sum_4[55]));
  AL_FADD comp4_56 (
    .a(i4[56]),
    .b(sum_3[56]),
    .c(cout_4[55]),
    .cout(cout_4[56]),
    .sum(sum_4[56]));
  AL_FADD comp4_57 (
    .a(1'b0),
    .b(sum_3[57]),
    .c(cout_4[56]),
    .cout(cout_4[57]),
    .sum(sum_4[57]));
  AL_FADD comp4_58 (
    .a(1'b0),
    .b(sum_3[58]),
    .c(cout_4[57]),
    .cout(cout_4[58]),
    .sum(sum_4[58]));
  AL_FADD comp4_59 (
    .a(1'b0),
    .b(sum_3[59]),
    .c(cout_4[58]),
    .cout(cout_4[59]),
    .sum(sum_4[59]));
  AL_FADD comp4_6 (
    .a(i4[6]),
    .b(sum_3[6]),
    .c(cout_4[5]),
    .cout(cout_4[6]),
    .sum(sum_4[6]));
  AL_FADD comp4_60 (
    .a(1'b0),
    .b(sum_3[60]),
    .c(cout_4[59]),
    .cout(cout_4[60]),
    .sum(sum_4[60]));
  AL_FADD comp4_61 (
    .a(1'b0),
    .b(sum_3[61]),
    .c(cout_4[60]),
    .cout(cout_4[61]),
    .sum(sum_4[61]));
  AL_FADD comp4_62 (
    .a(1'b0),
    .b(sum_3[62]),
    .c(cout_4[61]),
    .cout(cout_4[62]),
    .sum(sum_4[62]));
  AL_FADD comp4_63 (
    .a(1'b0),
    .b(sum_3[63]),
    .c(cout_4[62]),
    .cout(cout_4[63]),
    .sum(sum_4[63]));
  AL_FADD comp4_7 (
    .a(i4[7]),
    .b(sum_3[7]),
    .c(cout_4[6]),
    .cout(cout_4[7]),
    .sum(sum_4[7]));
  AL_FADD comp4_8 (
    .a(i4[8]),
    .b(sum_3[8]),
    .c(cout_4[7]),
    .cout(cout_4[8]),
    .sum(sum_4[8]));
  AL_FADD comp4_9 (
    .a(i4[9]),
    .b(sum_3[9]),
    .c(cout_4[8]),
    .cout(cout_4[9]),
    .sum(sum_4[9]));
  AL_FADD comp5_0 (
    .a(i5[0]),
    .b(sum_4[0]),
    .c(1'b0),
    .cout(cout_5[0]),
    .sum(sum_5[0]));
  AL_FADD comp5_1 (
    .a(i5[1]),
    .b(sum_4[1]),
    .c(cout_5[0]),
    .cout(cout_5[1]),
    .sum(sum_5[1]));
  AL_FADD comp5_10 (
    .a(i5[10]),
    .b(sum_4[10]),
    .c(cout_5[9]),
    .cout(cout_5[10]),
    .sum(sum_5[10]));
  AL_FADD comp5_11 (
    .a(i5[11]),
    .b(sum_4[11]),
    .c(cout_5[10]),
    .cout(cout_5[11]),
    .sum(sum_5[11]));
  AL_FADD comp5_12 (
    .a(i5[12]),
    .b(sum_4[12]),
    .c(cout_5[11]),
    .cout(cout_5[12]),
    .sum(sum_5[12]));
  AL_FADD comp5_13 (
    .a(i5[13]),
    .b(sum_4[13]),
    .c(cout_5[12]),
    .cout(cout_5[13]),
    .sum(sum_5[13]));
  AL_FADD comp5_14 (
    .a(i5[14]),
    .b(sum_4[14]),
    .c(cout_5[13]),
    .cout(cout_5[14]),
    .sum(sum_5[14]));
  AL_FADD comp5_15 (
    .a(i5[15]),
    .b(sum_4[15]),
    .c(cout_5[14]),
    .cout(cout_5[15]),
    .sum(sum_5[15]));
  AL_FADD comp5_16 (
    .a(i5[16]),
    .b(sum_4[16]),
    .c(cout_5[15]),
    .cout(cout_5[16]),
    .sum(sum_5[16]));
  AL_FADD comp5_17 (
    .a(i5[17]),
    .b(sum_4[17]),
    .c(cout_5[16]),
    .cout(cout_5[17]),
    .sum(sum_5[17]));
  AL_FADD comp5_18 (
    .a(i5[18]),
    .b(sum_4[18]),
    .c(cout_5[17]),
    .cout(cout_5[18]),
    .sum(sum_5[18]));
  AL_FADD comp5_19 (
    .a(i5[19]),
    .b(sum_4[19]),
    .c(cout_5[18]),
    .cout(cout_5[19]),
    .sum(sum_5[19]));
  AL_FADD comp5_2 (
    .a(i5[2]),
    .b(sum_4[2]),
    .c(cout_5[1]),
    .cout(cout_5[2]),
    .sum(sum_5[2]));
  AL_FADD comp5_20 (
    .a(i5[20]),
    .b(sum_4[20]),
    .c(cout_5[19]),
    .cout(cout_5[20]),
    .sum(sum_5[20]));
  AL_FADD comp5_21 (
    .a(i5[21]),
    .b(sum_4[21]),
    .c(cout_5[20]),
    .cout(cout_5[21]),
    .sum(sum_5[21]));
  AL_FADD comp5_22 (
    .a(i5[22]),
    .b(sum_4[22]),
    .c(cout_5[21]),
    .cout(cout_5[22]),
    .sum(sum_5[22]));
  AL_FADD comp5_23 (
    .a(i5[23]),
    .b(sum_4[23]),
    .c(cout_5[22]),
    .cout(cout_5[23]),
    .sum(sum_5[23]));
  AL_FADD comp5_24 (
    .a(i5[24]),
    .b(sum_4[24]),
    .c(cout_5[23]),
    .cout(cout_5[24]),
    .sum(sum_5[24]));
  AL_FADD comp5_25 (
    .a(i5[25]),
    .b(sum_4[25]),
    .c(cout_5[24]),
    .cout(cout_5[25]),
    .sum(sum_5[25]));
  AL_FADD comp5_26 (
    .a(i5[26]),
    .b(sum_4[26]),
    .c(cout_5[25]),
    .cout(cout_5[26]),
    .sum(sum_5[26]));
  AL_FADD comp5_27 (
    .a(i5[27]),
    .b(sum_4[27]),
    .c(cout_5[26]),
    .cout(cout_5[27]),
    .sum(sum_5[27]));
  AL_FADD comp5_28 (
    .a(i5[28]),
    .b(sum_4[28]),
    .c(cout_5[27]),
    .cout(cout_5[28]),
    .sum(sum_5[28]));
  AL_FADD comp5_29 (
    .a(i5[29]),
    .b(sum_4[29]),
    .c(cout_5[28]),
    .cout(cout_5[29]),
    .sum(sum_5[29]));
  AL_FADD comp5_3 (
    .a(i5[3]),
    .b(sum_4[3]),
    .c(cout_5[2]),
    .cout(cout_5[3]),
    .sum(sum_5[3]));
  AL_FADD comp5_30 (
    .a(i5[30]),
    .b(sum_4[30]),
    .c(cout_5[29]),
    .cout(cout_5[30]),
    .sum(sum_5[30]));
  AL_FADD comp5_31 (
    .a(i5[31]),
    .b(sum_4[31]),
    .c(cout_5[30]),
    .cout(cout_5[31]),
    .sum(sum_5[31]));
  AL_FADD comp5_32 (
    .a(i5[32]),
    .b(sum_4[32]),
    .c(cout_5[31]),
    .cout(cout_5[32]),
    .sum(sum_5[32]));
  AL_FADD comp5_33 (
    .a(i5[33]),
    .b(sum_4[33]),
    .c(cout_5[32]),
    .cout(cout_5[33]),
    .sum(sum_5[33]));
  AL_FADD comp5_34 (
    .a(i5[34]),
    .b(sum_4[34]),
    .c(cout_5[33]),
    .cout(cout_5[34]),
    .sum(sum_5[34]));
  AL_FADD comp5_35 (
    .a(i5[35]),
    .b(sum_4[35]),
    .c(cout_5[34]),
    .cout(cout_5[35]),
    .sum(sum_5[35]));
  AL_FADD comp5_36 (
    .a(i5[36]),
    .b(sum_4[36]),
    .c(cout_5[35]),
    .cout(cout_5[36]),
    .sum(sum_5[36]));
  AL_FADD comp5_37 (
    .a(i5[37]),
    .b(sum_4[37]),
    .c(cout_5[36]),
    .cout(cout_5[37]),
    .sum(sum_5[37]));
  AL_FADD comp5_38 (
    .a(i5[38]),
    .b(sum_4[38]),
    .c(cout_5[37]),
    .cout(cout_5[38]),
    .sum(sum_5[38]));
  AL_FADD comp5_39 (
    .a(i5[39]),
    .b(sum_4[39]),
    .c(cout_5[38]),
    .cout(cout_5[39]),
    .sum(sum_5[39]));
  AL_FADD comp5_4 (
    .a(i5[4]),
    .b(sum_4[4]),
    .c(cout_5[3]),
    .cout(cout_5[4]),
    .sum(sum_5[4]));
  AL_FADD comp5_40 (
    .a(i5[40]),
    .b(sum_4[40]),
    .c(cout_5[39]),
    .cout(cout_5[40]),
    .sum(sum_5[40]));
  AL_FADD comp5_41 (
    .a(i5[41]),
    .b(sum_4[41]),
    .c(cout_5[40]),
    .cout(cout_5[41]),
    .sum(sum_5[41]));
  AL_FADD comp5_42 (
    .a(i5[42]),
    .b(sum_4[42]),
    .c(cout_5[41]),
    .cout(cout_5[42]),
    .sum(sum_5[42]));
  AL_FADD comp5_43 (
    .a(i5[43]),
    .b(sum_4[43]),
    .c(cout_5[42]),
    .cout(cout_5[43]),
    .sum(sum_5[43]));
  AL_FADD comp5_44 (
    .a(i5[44]),
    .b(sum_4[44]),
    .c(cout_5[43]),
    .cout(cout_5[44]),
    .sum(sum_5[44]));
  AL_FADD comp5_45 (
    .a(i5[45]),
    .b(sum_4[45]),
    .c(cout_5[44]),
    .cout(cout_5[45]),
    .sum(sum_5[45]));
  AL_FADD comp5_46 (
    .a(i5[46]),
    .b(sum_4[46]),
    .c(cout_5[45]),
    .cout(cout_5[46]),
    .sum(sum_5[46]));
  AL_FADD comp5_47 (
    .a(i5[47]),
    .b(sum_4[47]),
    .c(cout_5[46]),
    .cout(cout_5[47]),
    .sum(sum_5[47]));
  AL_FADD comp5_48 (
    .a(i5[48]),
    .b(sum_4[48]),
    .c(cout_5[47]),
    .cout(cout_5[48]),
    .sum(sum_5[48]));
  AL_FADD comp5_49 (
    .a(i5[49]),
    .b(sum_4[49]),
    .c(cout_5[48]),
    .cout(cout_5[49]),
    .sum(sum_5[49]));
  AL_FADD comp5_5 (
    .a(i5[5]),
    .b(sum_4[5]),
    .c(cout_5[4]),
    .cout(cout_5[5]),
    .sum(sum_5[5]));
  AL_FADD comp5_50 (
    .a(i5[50]),
    .b(sum_4[50]),
    .c(cout_5[49]),
    .cout(cout_5[50]),
    .sum(sum_5[50]));
  AL_FADD comp5_51 (
    .a(i5[51]),
    .b(sum_4[51]),
    .c(cout_5[50]),
    .cout(cout_5[51]),
    .sum(sum_5[51]));
  AL_FADD comp5_52 (
    .a(i5[52]),
    .b(sum_4[52]),
    .c(cout_5[51]),
    .cout(cout_5[52]),
    .sum(sum_5[52]));
  AL_FADD comp5_53 (
    .a(i5[53]),
    .b(sum_4[53]),
    .c(cout_5[52]),
    .cout(cout_5[53]),
    .sum(sum_5[53]));
  AL_FADD comp5_54 (
    .a(i5[54]),
    .b(sum_4[54]),
    .c(cout_5[53]),
    .cout(cout_5[54]),
    .sum(sum_5[54]));
  AL_FADD comp5_55 (
    .a(i5[55]),
    .b(sum_4[55]),
    .c(cout_5[54]),
    .cout(cout_5[55]),
    .sum(sum_5[55]));
  AL_FADD comp5_56 (
    .a(1'b0),
    .b(sum_4[56]),
    .c(cout_5[55]),
    .cout(cout_5[56]),
    .sum(sum_5[56]));
  AL_FADD comp5_57 (
    .a(1'b0),
    .b(sum_4[57]),
    .c(cout_5[56]),
    .cout(cout_5[57]),
    .sum(sum_5[57]));
  AL_FADD comp5_58 (
    .a(1'b0),
    .b(sum_4[58]),
    .c(cout_5[57]),
    .cout(cout_5[58]),
    .sum(sum_5[58]));
  AL_FADD comp5_59 (
    .a(1'b0),
    .b(sum_4[59]),
    .c(cout_5[58]),
    .cout(cout_5[59]),
    .sum(sum_5[59]));
  AL_FADD comp5_6 (
    .a(i5[6]),
    .b(sum_4[6]),
    .c(cout_5[5]),
    .cout(cout_5[6]),
    .sum(sum_5[6]));
  AL_FADD comp5_60 (
    .a(1'b0),
    .b(sum_4[60]),
    .c(cout_5[59]),
    .cout(cout_5[60]),
    .sum(sum_5[60]));
  AL_FADD comp5_61 (
    .a(1'b0),
    .b(sum_4[61]),
    .c(cout_5[60]),
    .cout(cout_5[61]),
    .sum(sum_5[61]));
  AL_FADD comp5_62 (
    .a(1'b0),
    .b(sum_4[62]),
    .c(cout_5[61]),
    .cout(cout_5[62]),
    .sum(sum_5[62]));
  AL_FADD comp5_63 (
    .a(1'b0),
    .b(sum_4[63]),
    .c(cout_5[62]),
    .cout(cout_5[63]),
    .sum(sum_5[63]));
  AL_FADD comp5_7 (
    .a(i5[7]),
    .b(sum_4[7]),
    .c(cout_5[6]),
    .cout(cout_5[7]),
    .sum(sum_5[7]));
  AL_FADD comp5_8 (
    .a(i5[8]),
    .b(sum_4[8]),
    .c(cout_5[7]),
    .cout(cout_5[8]),
    .sum(sum_5[8]));
  AL_FADD comp5_9 (
    .a(i5[9]),
    .b(sum_4[9]),
    .c(cout_5[8]),
    .cout(cout_5[9]),
    .sum(sum_5[9]));
  AL_FADD comp6_0 (
    .a(i6[0]),
    .b(sum_5[0]),
    .c(1'b0),
    .cout(cout_6[0]),
    .sum(sum_6[0]));
  AL_FADD comp6_1 (
    .a(i6[1]),
    .b(sum_5[1]),
    .c(cout_6[0]),
    .cout(cout_6[1]),
    .sum(sum_6[1]));
  AL_FADD comp6_10 (
    .a(i6[10]),
    .b(sum_5[10]),
    .c(cout_6[9]),
    .cout(cout_6[10]),
    .sum(sum_6[10]));
  AL_FADD comp6_11 (
    .a(i6[11]),
    .b(sum_5[11]),
    .c(cout_6[10]),
    .cout(cout_6[11]),
    .sum(sum_6[11]));
  AL_FADD comp6_12 (
    .a(i6[12]),
    .b(sum_5[12]),
    .c(cout_6[11]),
    .cout(cout_6[12]),
    .sum(sum_6[12]));
  AL_FADD comp6_13 (
    .a(i6[13]),
    .b(sum_5[13]),
    .c(cout_6[12]),
    .cout(cout_6[13]),
    .sum(sum_6[13]));
  AL_FADD comp6_14 (
    .a(i6[14]),
    .b(sum_5[14]),
    .c(cout_6[13]),
    .cout(cout_6[14]),
    .sum(sum_6[14]));
  AL_FADD comp6_15 (
    .a(i6[15]),
    .b(sum_5[15]),
    .c(cout_6[14]),
    .cout(cout_6[15]),
    .sum(sum_6[15]));
  AL_FADD comp6_16 (
    .a(i6[16]),
    .b(sum_5[16]),
    .c(cout_6[15]),
    .cout(cout_6[16]),
    .sum(sum_6[16]));
  AL_FADD comp6_17 (
    .a(i6[17]),
    .b(sum_5[17]),
    .c(cout_6[16]),
    .cout(cout_6[17]),
    .sum(sum_6[17]));
  AL_FADD comp6_18 (
    .a(i6[18]),
    .b(sum_5[18]),
    .c(cout_6[17]),
    .cout(cout_6[18]),
    .sum(sum_6[18]));
  AL_FADD comp6_19 (
    .a(i6[19]),
    .b(sum_5[19]),
    .c(cout_6[18]),
    .cout(cout_6[19]),
    .sum(sum_6[19]));
  AL_FADD comp6_2 (
    .a(i6[2]),
    .b(sum_5[2]),
    .c(cout_6[1]),
    .cout(cout_6[2]),
    .sum(sum_6[2]));
  AL_FADD comp6_20 (
    .a(i6[20]),
    .b(sum_5[20]),
    .c(cout_6[19]),
    .cout(cout_6[20]),
    .sum(sum_6[20]));
  AL_FADD comp6_21 (
    .a(i6[21]),
    .b(sum_5[21]),
    .c(cout_6[20]),
    .cout(cout_6[21]),
    .sum(sum_6[21]));
  AL_FADD comp6_22 (
    .a(i6[22]),
    .b(sum_5[22]),
    .c(cout_6[21]),
    .cout(cout_6[22]),
    .sum(sum_6[22]));
  AL_FADD comp6_23 (
    .a(i6[23]),
    .b(sum_5[23]),
    .c(cout_6[22]),
    .cout(cout_6[23]),
    .sum(sum_6[23]));
  AL_FADD comp6_24 (
    .a(i6[24]),
    .b(sum_5[24]),
    .c(cout_6[23]),
    .cout(cout_6[24]),
    .sum(sum_6[24]));
  AL_FADD comp6_25 (
    .a(i6[25]),
    .b(sum_5[25]),
    .c(cout_6[24]),
    .cout(cout_6[25]),
    .sum(sum_6[25]));
  AL_FADD comp6_26 (
    .a(i6[26]),
    .b(sum_5[26]),
    .c(cout_6[25]),
    .cout(cout_6[26]),
    .sum(sum_6[26]));
  AL_FADD comp6_27 (
    .a(i6[27]),
    .b(sum_5[27]),
    .c(cout_6[26]),
    .cout(cout_6[27]),
    .sum(sum_6[27]));
  AL_FADD comp6_28 (
    .a(i6[28]),
    .b(sum_5[28]),
    .c(cout_6[27]),
    .cout(cout_6[28]),
    .sum(sum_6[28]));
  AL_FADD comp6_29 (
    .a(i6[29]),
    .b(sum_5[29]),
    .c(cout_6[28]),
    .cout(cout_6[29]),
    .sum(sum_6[29]));
  AL_FADD comp6_3 (
    .a(i6[3]),
    .b(sum_5[3]),
    .c(cout_6[2]),
    .cout(cout_6[3]),
    .sum(sum_6[3]));
  AL_FADD comp6_30 (
    .a(i6[30]),
    .b(sum_5[30]),
    .c(cout_6[29]),
    .cout(cout_6[30]),
    .sum(sum_6[30]));
  AL_FADD comp6_31 (
    .a(i6[31]),
    .b(sum_5[31]),
    .c(cout_6[30]),
    .cout(cout_6[31]),
    .sum(sum_6[31]));
  AL_FADD comp6_32 (
    .a(i6[32]),
    .b(sum_5[32]),
    .c(cout_6[31]),
    .cout(cout_6[32]),
    .sum(sum_6[32]));
  AL_FADD comp6_33 (
    .a(i6[33]),
    .b(sum_5[33]),
    .c(cout_6[32]),
    .cout(cout_6[33]),
    .sum(sum_6[33]));
  AL_FADD comp6_34 (
    .a(i6[34]),
    .b(sum_5[34]),
    .c(cout_6[33]),
    .cout(cout_6[34]),
    .sum(sum_6[34]));
  AL_FADD comp6_35 (
    .a(i6[35]),
    .b(sum_5[35]),
    .c(cout_6[34]),
    .cout(cout_6[35]),
    .sum(sum_6[35]));
  AL_FADD comp6_36 (
    .a(i6[36]),
    .b(sum_5[36]),
    .c(cout_6[35]),
    .cout(cout_6[36]),
    .sum(sum_6[36]));
  AL_FADD comp6_37 (
    .a(i6[37]),
    .b(sum_5[37]),
    .c(cout_6[36]),
    .cout(cout_6[37]),
    .sum(sum_6[37]));
  AL_FADD comp6_38 (
    .a(i6[38]),
    .b(sum_5[38]),
    .c(cout_6[37]),
    .cout(cout_6[38]),
    .sum(sum_6[38]));
  AL_FADD comp6_39 (
    .a(i6[39]),
    .b(sum_5[39]),
    .c(cout_6[38]),
    .cout(cout_6[39]),
    .sum(sum_6[39]));
  AL_FADD comp6_4 (
    .a(i6[4]),
    .b(sum_5[4]),
    .c(cout_6[3]),
    .cout(cout_6[4]),
    .sum(sum_6[4]));
  AL_FADD comp6_40 (
    .a(i6[40]),
    .b(sum_5[40]),
    .c(cout_6[39]),
    .cout(cout_6[40]),
    .sum(sum_6[40]));
  AL_FADD comp6_41 (
    .a(i6[41]),
    .b(sum_5[41]),
    .c(cout_6[40]),
    .cout(cout_6[41]),
    .sum(sum_6[41]));
  AL_FADD comp6_42 (
    .a(i6[42]),
    .b(sum_5[42]),
    .c(cout_6[41]),
    .cout(cout_6[42]),
    .sum(sum_6[42]));
  AL_FADD comp6_43 (
    .a(i6[43]),
    .b(sum_5[43]),
    .c(cout_6[42]),
    .cout(cout_6[43]),
    .sum(sum_6[43]));
  AL_FADD comp6_44 (
    .a(i6[44]),
    .b(sum_5[44]),
    .c(cout_6[43]),
    .cout(cout_6[44]),
    .sum(sum_6[44]));
  AL_FADD comp6_45 (
    .a(i6[45]),
    .b(sum_5[45]),
    .c(cout_6[44]),
    .cout(cout_6[45]),
    .sum(sum_6[45]));
  AL_FADD comp6_46 (
    .a(i6[46]),
    .b(sum_5[46]),
    .c(cout_6[45]),
    .cout(cout_6[46]),
    .sum(sum_6[46]));
  AL_FADD comp6_47 (
    .a(i6[47]),
    .b(sum_5[47]),
    .c(cout_6[46]),
    .cout(cout_6[47]),
    .sum(sum_6[47]));
  AL_FADD comp6_48 (
    .a(i6[48]),
    .b(sum_5[48]),
    .c(cout_6[47]),
    .cout(cout_6[48]),
    .sum(sum_6[48]));
  AL_FADD comp6_49 (
    .a(i6[49]),
    .b(sum_5[49]),
    .c(cout_6[48]),
    .cout(cout_6[49]),
    .sum(sum_6[49]));
  AL_FADD comp6_5 (
    .a(i6[5]),
    .b(sum_5[5]),
    .c(cout_6[4]),
    .cout(cout_6[5]),
    .sum(sum_6[5]));
  AL_FADD comp6_50 (
    .a(i6[50]),
    .b(sum_5[50]),
    .c(cout_6[49]),
    .cout(cout_6[50]),
    .sum(sum_6[50]));
  AL_FADD comp6_51 (
    .a(i6[51]),
    .b(sum_5[51]),
    .c(cout_6[50]),
    .cout(cout_6[51]),
    .sum(sum_6[51]));
  AL_FADD comp6_52 (
    .a(i6[52]),
    .b(sum_5[52]),
    .c(cout_6[51]),
    .cout(cout_6[52]),
    .sum(sum_6[52]));
  AL_FADD comp6_53 (
    .a(i6[53]),
    .b(sum_5[53]),
    .c(cout_6[52]),
    .cout(cout_6[53]),
    .sum(sum_6[53]));
  AL_FADD comp6_54 (
    .a(i6[54]),
    .b(sum_5[54]),
    .c(cout_6[53]),
    .cout(cout_6[54]),
    .sum(sum_6[54]));
  AL_FADD comp6_55 (
    .a(1'b0),
    .b(sum_5[55]),
    .c(cout_6[54]),
    .cout(cout_6[55]),
    .sum(sum_6[55]));
  AL_FADD comp6_56 (
    .a(1'b0),
    .b(sum_5[56]),
    .c(cout_6[55]),
    .cout(cout_6[56]),
    .sum(sum_6[56]));
  AL_FADD comp6_57 (
    .a(1'b0),
    .b(sum_5[57]),
    .c(cout_6[56]),
    .cout(cout_6[57]),
    .sum(sum_6[57]));
  AL_FADD comp6_58 (
    .a(1'b0),
    .b(sum_5[58]),
    .c(cout_6[57]),
    .cout(cout_6[58]),
    .sum(sum_6[58]));
  AL_FADD comp6_59 (
    .a(1'b0),
    .b(sum_5[59]),
    .c(cout_6[58]),
    .cout(cout_6[59]),
    .sum(sum_6[59]));
  AL_FADD comp6_6 (
    .a(i6[6]),
    .b(sum_5[6]),
    .c(cout_6[5]),
    .cout(cout_6[6]),
    .sum(sum_6[6]));
  AL_FADD comp6_60 (
    .a(1'b0),
    .b(sum_5[60]),
    .c(cout_6[59]),
    .cout(cout_6[60]),
    .sum(sum_6[60]));
  AL_FADD comp6_61 (
    .a(1'b0),
    .b(sum_5[61]),
    .c(cout_6[60]),
    .cout(cout_6[61]),
    .sum(sum_6[61]));
  AL_FADD comp6_62 (
    .a(1'b0),
    .b(sum_5[62]),
    .c(cout_6[61]),
    .cout(cout_6[62]),
    .sum(sum_6[62]));
  AL_FADD comp6_63 (
    .a(1'b0),
    .b(sum_5[63]),
    .c(cout_6[62]),
    .cout(cout_6[63]),
    .sum(sum_6[63]));
  AL_FADD comp6_7 (
    .a(i6[7]),
    .b(sum_5[7]),
    .c(cout_6[6]),
    .cout(cout_6[7]),
    .sum(sum_6[7]));
  AL_FADD comp6_8 (
    .a(i6[8]),
    .b(sum_5[8]),
    .c(cout_6[7]),
    .cout(cout_6[8]),
    .sum(sum_6[8]));
  AL_FADD comp6_9 (
    .a(i6[9]),
    .b(sum_5[9]),
    .c(cout_6[8]),
    .cout(cout_6[9]),
    .sum(sum_6[9]));
  AL_FADD comp7_0 (
    .a(i7[0]),
    .b(sum_6[0]),
    .c(1'b0),
    .cout(cout_7[0]),
    .sum(sum_7[0]));
  AL_FADD comp7_1 (
    .a(i7[1]),
    .b(sum_6[1]),
    .c(cout_7[0]),
    .cout(cout_7[1]),
    .sum(sum_7[1]));
  AL_FADD comp7_10 (
    .a(i7[10]),
    .b(sum_6[10]),
    .c(cout_7[9]),
    .cout(cout_7[10]),
    .sum(sum_7[10]));
  AL_FADD comp7_11 (
    .a(i7[11]),
    .b(sum_6[11]),
    .c(cout_7[10]),
    .cout(cout_7[11]),
    .sum(sum_7[11]));
  AL_FADD comp7_12 (
    .a(i7[12]),
    .b(sum_6[12]),
    .c(cout_7[11]),
    .cout(cout_7[12]),
    .sum(sum_7[12]));
  AL_FADD comp7_13 (
    .a(i7[13]),
    .b(sum_6[13]),
    .c(cout_7[12]),
    .cout(cout_7[13]),
    .sum(sum_7[13]));
  AL_FADD comp7_14 (
    .a(i7[14]),
    .b(sum_6[14]),
    .c(cout_7[13]),
    .cout(cout_7[14]),
    .sum(sum_7[14]));
  AL_FADD comp7_15 (
    .a(i7[15]),
    .b(sum_6[15]),
    .c(cout_7[14]),
    .cout(cout_7[15]),
    .sum(sum_7[15]));
  AL_FADD comp7_16 (
    .a(i7[16]),
    .b(sum_6[16]),
    .c(cout_7[15]),
    .cout(cout_7[16]),
    .sum(sum_7[16]));
  AL_FADD comp7_17 (
    .a(i7[17]),
    .b(sum_6[17]),
    .c(cout_7[16]),
    .cout(cout_7[17]),
    .sum(sum_7[17]));
  AL_FADD comp7_18 (
    .a(i7[18]),
    .b(sum_6[18]),
    .c(cout_7[17]),
    .cout(cout_7[18]),
    .sum(sum_7[18]));
  AL_FADD comp7_19 (
    .a(i7[19]),
    .b(sum_6[19]),
    .c(cout_7[18]),
    .cout(cout_7[19]),
    .sum(sum_7[19]));
  AL_FADD comp7_2 (
    .a(i7[2]),
    .b(sum_6[2]),
    .c(cout_7[1]),
    .cout(cout_7[2]),
    .sum(sum_7[2]));
  AL_FADD comp7_20 (
    .a(i7[20]),
    .b(sum_6[20]),
    .c(cout_7[19]),
    .cout(cout_7[20]),
    .sum(sum_7[20]));
  AL_FADD comp7_21 (
    .a(i7[21]),
    .b(sum_6[21]),
    .c(cout_7[20]),
    .cout(cout_7[21]),
    .sum(sum_7[21]));
  AL_FADD comp7_22 (
    .a(i7[22]),
    .b(sum_6[22]),
    .c(cout_7[21]),
    .cout(cout_7[22]),
    .sum(sum_7[22]));
  AL_FADD comp7_23 (
    .a(i7[23]),
    .b(sum_6[23]),
    .c(cout_7[22]),
    .cout(cout_7[23]),
    .sum(sum_7[23]));
  AL_FADD comp7_24 (
    .a(i7[24]),
    .b(sum_6[24]),
    .c(cout_7[23]),
    .cout(cout_7[24]),
    .sum(sum_7[24]));
  AL_FADD comp7_25 (
    .a(i7[25]),
    .b(sum_6[25]),
    .c(cout_7[24]),
    .cout(cout_7[25]),
    .sum(sum_7[25]));
  AL_FADD comp7_26 (
    .a(i7[26]),
    .b(sum_6[26]),
    .c(cout_7[25]),
    .cout(cout_7[26]),
    .sum(sum_7[26]));
  AL_FADD comp7_27 (
    .a(i7[27]),
    .b(sum_6[27]),
    .c(cout_7[26]),
    .cout(cout_7[27]),
    .sum(sum_7[27]));
  AL_FADD comp7_28 (
    .a(i7[28]),
    .b(sum_6[28]),
    .c(cout_7[27]),
    .cout(cout_7[28]),
    .sum(sum_7[28]));
  AL_FADD comp7_29 (
    .a(i7[29]),
    .b(sum_6[29]),
    .c(cout_7[28]),
    .cout(cout_7[29]),
    .sum(sum_7[29]));
  AL_FADD comp7_3 (
    .a(i7[3]),
    .b(sum_6[3]),
    .c(cout_7[2]),
    .cout(cout_7[3]),
    .sum(sum_7[3]));
  AL_FADD comp7_30 (
    .a(i7[30]),
    .b(sum_6[30]),
    .c(cout_7[29]),
    .cout(cout_7[30]),
    .sum(sum_7[30]));
  AL_FADD comp7_31 (
    .a(i7[31]),
    .b(sum_6[31]),
    .c(cout_7[30]),
    .cout(cout_7[31]),
    .sum(sum_7[31]));
  AL_FADD comp7_32 (
    .a(i7[32]),
    .b(sum_6[32]),
    .c(cout_7[31]),
    .cout(cout_7[32]),
    .sum(sum_7[32]));
  AL_FADD comp7_33 (
    .a(i7[33]),
    .b(sum_6[33]),
    .c(cout_7[32]),
    .cout(cout_7[33]),
    .sum(sum_7[33]));
  AL_FADD comp7_34 (
    .a(i7[34]),
    .b(sum_6[34]),
    .c(cout_7[33]),
    .cout(cout_7[34]),
    .sum(sum_7[34]));
  AL_FADD comp7_35 (
    .a(i7[35]),
    .b(sum_6[35]),
    .c(cout_7[34]),
    .cout(cout_7[35]),
    .sum(sum_7[35]));
  AL_FADD comp7_36 (
    .a(i7[36]),
    .b(sum_6[36]),
    .c(cout_7[35]),
    .cout(cout_7[36]),
    .sum(sum_7[36]));
  AL_FADD comp7_37 (
    .a(i7[37]),
    .b(sum_6[37]),
    .c(cout_7[36]),
    .cout(cout_7[37]),
    .sum(sum_7[37]));
  AL_FADD comp7_38 (
    .a(i7[38]),
    .b(sum_6[38]),
    .c(cout_7[37]),
    .cout(cout_7[38]),
    .sum(sum_7[38]));
  AL_FADD comp7_39 (
    .a(i7[39]),
    .b(sum_6[39]),
    .c(cout_7[38]),
    .cout(cout_7[39]),
    .sum(sum_7[39]));
  AL_FADD comp7_4 (
    .a(i7[4]),
    .b(sum_6[4]),
    .c(cout_7[3]),
    .cout(cout_7[4]),
    .sum(sum_7[4]));
  AL_FADD comp7_40 (
    .a(i7[40]),
    .b(sum_6[40]),
    .c(cout_7[39]),
    .cout(cout_7[40]),
    .sum(sum_7[40]));
  AL_FADD comp7_41 (
    .a(i7[41]),
    .b(sum_6[41]),
    .c(cout_7[40]),
    .cout(cout_7[41]),
    .sum(sum_7[41]));
  AL_FADD comp7_42 (
    .a(i7[42]),
    .b(sum_6[42]),
    .c(cout_7[41]),
    .cout(cout_7[42]),
    .sum(sum_7[42]));
  AL_FADD comp7_43 (
    .a(i7[43]),
    .b(sum_6[43]),
    .c(cout_7[42]),
    .cout(cout_7[43]),
    .sum(sum_7[43]));
  AL_FADD comp7_44 (
    .a(i7[44]),
    .b(sum_6[44]),
    .c(cout_7[43]),
    .cout(cout_7[44]),
    .sum(sum_7[44]));
  AL_FADD comp7_45 (
    .a(i7[45]),
    .b(sum_6[45]),
    .c(cout_7[44]),
    .cout(cout_7[45]),
    .sum(sum_7[45]));
  AL_FADD comp7_46 (
    .a(i7[46]),
    .b(sum_6[46]),
    .c(cout_7[45]),
    .cout(cout_7[46]),
    .sum(sum_7[46]));
  AL_FADD comp7_47 (
    .a(i7[47]),
    .b(sum_6[47]),
    .c(cout_7[46]),
    .cout(cout_7[47]),
    .sum(sum_7[47]));
  AL_FADD comp7_48 (
    .a(i7[48]),
    .b(sum_6[48]),
    .c(cout_7[47]),
    .cout(cout_7[48]),
    .sum(sum_7[48]));
  AL_FADD comp7_49 (
    .a(i7[49]),
    .b(sum_6[49]),
    .c(cout_7[48]),
    .cout(cout_7[49]),
    .sum(sum_7[49]));
  AL_FADD comp7_5 (
    .a(i7[5]),
    .b(sum_6[5]),
    .c(cout_7[4]),
    .cout(cout_7[5]),
    .sum(sum_7[5]));
  AL_FADD comp7_50 (
    .a(i7[50]),
    .b(sum_6[50]),
    .c(cout_7[49]),
    .cout(cout_7[50]),
    .sum(sum_7[50]));
  AL_FADD comp7_51 (
    .a(i7[51]),
    .b(sum_6[51]),
    .c(cout_7[50]),
    .cout(cout_7[51]),
    .sum(sum_7[51]));
  AL_FADD comp7_52 (
    .a(i7[52]),
    .b(sum_6[52]),
    .c(cout_7[51]),
    .cout(cout_7[52]),
    .sum(sum_7[52]));
  AL_FADD comp7_53 (
    .a(i7[53]),
    .b(sum_6[53]),
    .c(cout_7[52]),
    .cout(cout_7[53]),
    .sum(sum_7[53]));
  AL_FADD comp7_54 (
    .a(1'b0),
    .b(sum_6[54]),
    .c(cout_7[53]),
    .cout(cout_7[54]),
    .sum(sum_7[54]));
  AL_FADD comp7_55 (
    .a(1'b0),
    .b(sum_6[55]),
    .c(cout_7[54]),
    .cout(cout_7[55]),
    .sum(sum_7[55]));
  AL_FADD comp7_56 (
    .a(1'b0),
    .b(sum_6[56]),
    .c(cout_7[55]),
    .cout(cout_7[56]),
    .sum(sum_7[56]));
  AL_FADD comp7_57 (
    .a(1'b0),
    .b(sum_6[57]),
    .c(cout_7[56]),
    .cout(cout_7[57]),
    .sum(sum_7[57]));
  AL_FADD comp7_58 (
    .a(1'b0),
    .b(sum_6[58]),
    .c(cout_7[57]),
    .cout(cout_7[58]),
    .sum(sum_7[58]));
  AL_FADD comp7_59 (
    .a(1'b0),
    .b(sum_6[59]),
    .c(cout_7[58]),
    .cout(cout_7[59]),
    .sum(sum_7[59]));
  AL_FADD comp7_6 (
    .a(i7[6]),
    .b(sum_6[6]),
    .c(cout_7[5]),
    .cout(cout_7[6]),
    .sum(sum_7[6]));
  AL_FADD comp7_60 (
    .a(1'b0),
    .b(sum_6[60]),
    .c(cout_7[59]),
    .cout(cout_7[60]),
    .sum(sum_7[60]));
  AL_FADD comp7_61 (
    .a(1'b0),
    .b(sum_6[61]),
    .c(cout_7[60]),
    .cout(cout_7[61]),
    .sum(sum_7[61]));
  AL_FADD comp7_62 (
    .a(1'b0),
    .b(sum_6[62]),
    .c(cout_7[61]),
    .cout(cout_7[62]),
    .sum(sum_7[62]));
  AL_FADD comp7_63 (
    .a(1'b0),
    .b(sum_6[63]),
    .c(cout_7[62]),
    .cout(cout_7[63]),
    .sum(sum_7[63]));
  AL_FADD comp7_7 (
    .a(i7[7]),
    .b(sum_6[7]),
    .c(cout_7[6]),
    .cout(cout_7[7]),
    .sum(sum_7[7]));
  AL_FADD comp7_8 (
    .a(i7[8]),
    .b(sum_6[8]),
    .c(cout_7[7]),
    .cout(cout_7[8]),
    .sum(sum_7[8]));
  AL_FADD comp7_9 (
    .a(i7[9]),
    .b(sum_6[9]),
    .c(cout_7[8]),
    .cout(cout_7[9]),
    .sum(sum_7[9]));
  AL_FADD comp8_0 (
    .a(i8[0]),
    .b(sum_7[0]),
    .c(1'b0),
    .cout(cout_8[0]),
    .sum(sum_8[0]));
  AL_FADD comp8_1 (
    .a(i8[1]),
    .b(sum_7[1]),
    .c(cout_8[0]),
    .cout(cout_8[1]),
    .sum(sum_8[1]));
  AL_FADD comp8_10 (
    .a(i8[10]),
    .b(sum_7[10]),
    .c(cout_8[9]),
    .cout(cout_8[10]),
    .sum(sum_8[10]));
  AL_FADD comp8_11 (
    .a(i8[11]),
    .b(sum_7[11]),
    .c(cout_8[10]),
    .cout(cout_8[11]),
    .sum(sum_8[11]));
  AL_FADD comp8_12 (
    .a(i8[12]),
    .b(sum_7[12]),
    .c(cout_8[11]),
    .cout(cout_8[12]),
    .sum(sum_8[12]));
  AL_FADD comp8_13 (
    .a(i8[13]),
    .b(sum_7[13]),
    .c(cout_8[12]),
    .cout(cout_8[13]),
    .sum(sum_8[13]));
  AL_FADD comp8_14 (
    .a(i8[14]),
    .b(sum_7[14]),
    .c(cout_8[13]),
    .cout(cout_8[14]),
    .sum(sum_8[14]));
  AL_FADD comp8_15 (
    .a(i8[15]),
    .b(sum_7[15]),
    .c(cout_8[14]),
    .cout(cout_8[15]),
    .sum(sum_8[15]));
  AL_FADD comp8_16 (
    .a(i8[16]),
    .b(sum_7[16]),
    .c(cout_8[15]),
    .cout(cout_8[16]),
    .sum(sum_8[16]));
  AL_FADD comp8_17 (
    .a(i8[17]),
    .b(sum_7[17]),
    .c(cout_8[16]),
    .cout(cout_8[17]),
    .sum(sum_8[17]));
  AL_FADD comp8_18 (
    .a(i8[18]),
    .b(sum_7[18]),
    .c(cout_8[17]),
    .cout(cout_8[18]),
    .sum(sum_8[18]));
  AL_FADD comp8_19 (
    .a(i8[19]),
    .b(sum_7[19]),
    .c(cout_8[18]),
    .cout(cout_8[19]),
    .sum(sum_8[19]));
  AL_FADD comp8_2 (
    .a(i8[2]),
    .b(sum_7[2]),
    .c(cout_8[1]),
    .cout(cout_8[2]),
    .sum(sum_8[2]));
  AL_FADD comp8_20 (
    .a(i8[20]),
    .b(sum_7[20]),
    .c(cout_8[19]),
    .cout(cout_8[20]),
    .sum(sum_8[20]));
  AL_FADD comp8_21 (
    .a(i8[21]),
    .b(sum_7[21]),
    .c(cout_8[20]),
    .cout(cout_8[21]),
    .sum(sum_8[21]));
  AL_FADD comp8_22 (
    .a(i8[22]),
    .b(sum_7[22]),
    .c(cout_8[21]),
    .cout(cout_8[22]),
    .sum(sum_8[22]));
  AL_FADD comp8_23 (
    .a(i8[23]),
    .b(sum_7[23]),
    .c(cout_8[22]),
    .cout(cout_8[23]),
    .sum(sum_8[23]));
  AL_FADD comp8_24 (
    .a(i8[24]),
    .b(sum_7[24]),
    .c(cout_8[23]),
    .cout(cout_8[24]),
    .sum(sum_8[24]));
  AL_FADD comp8_25 (
    .a(i8[25]),
    .b(sum_7[25]),
    .c(cout_8[24]),
    .cout(cout_8[25]),
    .sum(sum_8[25]));
  AL_FADD comp8_26 (
    .a(i8[26]),
    .b(sum_7[26]),
    .c(cout_8[25]),
    .cout(cout_8[26]),
    .sum(sum_8[26]));
  AL_FADD comp8_27 (
    .a(i8[27]),
    .b(sum_7[27]),
    .c(cout_8[26]),
    .cout(cout_8[27]),
    .sum(sum_8[27]));
  AL_FADD comp8_28 (
    .a(i8[28]),
    .b(sum_7[28]),
    .c(cout_8[27]),
    .cout(cout_8[28]),
    .sum(sum_8[28]));
  AL_FADD comp8_29 (
    .a(i8[29]),
    .b(sum_7[29]),
    .c(cout_8[28]),
    .cout(cout_8[29]),
    .sum(sum_8[29]));
  AL_FADD comp8_3 (
    .a(i8[3]),
    .b(sum_7[3]),
    .c(cout_8[2]),
    .cout(cout_8[3]),
    .sum(sum_8[3]));
  AL_FADD comp8_30 (
    .a(i8[30]),
    .b(sum_7[30]),
    .c(cout_8[29]),
    .cout(cout_8[30]),
    .sum(sum_8[30]));
  AL_FADD comp8_31 (
    .a(i8[31]),
    .b(sum_7[31]),
    .c(cout_8[30]),
    .cout(cout_8[31]),
    .sum(sum_8[31]));
  AL_FADD comp8_32 (
    .a(i8[32]),
    .b(sum_7[32]),
    .c(cout_8[31]),
    .cout(cout_8[32]),
    .sum(sum_8[32]));
  AL_FADD comp8_33 (
    .a(i8[33]),
    .b(sum_7[33]),
    .c(cout_8[32]),
    .cout(cout_8[33]),
    .sum(sum_8[33]));
  AL_FADD comp8_34 (
    .a(i8[34]),
    .b(sum_7[34]),
    .c(cout_8[33]),
    .cout(cout_8[34]),
    .sum(sum_8[34]));
  AL_FADD comp8_35 (
    .a(i8[35]),
    .b(sum_7[35]),
    .c(cout_8[34]),
    .cout(cout_8[35]),
    .sum(sum_8[35]));
  AL_FADD comp8_36 (
    .a(i8[36]),
    .b(sum_7[36]),
    .c(cout_8[35]),
    .cout(cout_8[36]),
    .sum(sum_8[36]));
  AL_FADD comp8_37 (
    .a(i8[37]),
    .b(sum_7[37]),
    .c(cout_8[36]),
    .cout(cout_8[37]),
    .sum(sum_8[37]));
  AL_FADD comp8_38 (
    .a(i8[38]),
    .b(sum_7[38]),
    .c(cout_8[37]),
    .cout(cout_8[38]),
    .sum(sum_8[38]));
  AL_FADD comp8_39 (
    .a(i8[39]),
    .b(sum_7[39]),
    .c(cout_8[38]),
    .cout(cout_8[39]),
    .sum(sum_8[39]));
  AL_FADD comp8_4 (
    .a(i8[4]),
    .b(sum_7[4]),
    .c(cout_8[3]),
    .cout(cout_8[4]),
    .sum(sum_8[4]));
  AL_FADD comp8_40 (
    .a(i8[40]),
    .b(sum_7[40]),
    .c(cout_8[39]),
    .cout(cout_8[40]),
    .sum(sum_8[40]));
  AL_FADD comp8_41 (
    .a(i8[41]),
    .b(sum_7[41]),
    .c(cout_8[40]),
    .cout(cout_8[41]),
    .sum(sum_8[41]));
  AL_FADD comp8_42 (
    .a(i8[42]),
    .b(sum_7[42]),
    .c(cout_8[41]),
    .cout(cout_8[42]),
    .sum(sum_8[42]));
  AL_FADD comp8_43 (
    .a(i8[43]),
    .b(sum_7[43]),
    .c(cout_8[42]),
    .cout(cout_8[43]),
    .sum(sum_8[43]));
  AL_FADD comp8_44 (
    .a(i8[44]),
    .b(sum_7[44]),
    .c(cout_8[43]),
    .cout(cout_8[44]),
    .sum(sum_8[44]));
  AL_FADD comp8_45 (
    .a(i8[45]),
    .b(sum_7[45]),
    .c(cout_8[44]),
    .cout(cout_8[45]),
    .sum(sum_8[45]));
  AL_FADD comp8_46 (
    .a(i8[46]),
    .b(sum_7[46]),
    .c(cout_8[45]),
    .cout(cout_8[46]),
    .sum(sum_8[46]));
  AL_FADD comp8_47 (
    .a(i8[47]),
    .b(sum_7[47]),
    .c(cout_8[46]),
    .cout(cout_8[47]),
    .sum(sum_8[47]));
  AL_FADD comp8_48 (
    .a(i8[48]),
    .b(sum_7[48]),
    .c(cout_8[47]),
    .cout(cout_8[48]),
    .sum(sum_8[48]));
  AL_FADD comp8_49 (
    .a(i8[49]),
    .b(sum_7[49]),
    .c(cout_8[48]),
    .cout(cout_8[49]),
    .sum(sum_8[49]));
  AL_FADD comp8_5 (
    .a(i8[5]),
    .b(sum_7[5]),
    .c(cout_8[4]),
    .cout(cout_8[5]),
    .sum(sum_8[5]));
  AL_FADD comp8_50 (
    .a(i8[50]),
    .b(sum_7[50]),
    .c(cout_8[49]),
    .cout(cout_8[50]),
    .sum(sum_8[50]));
  AL_FADD comp8_51 (
    .a(i8[51]),
    .b(sum_7[51]),
    .c(cout_8[50]),
    .cout(cout_8[51]),
    .sum(sum_8[51]));
  AL_FADD comp8_52 (
    .a(i8[52]),
    .b(sum_7[52]),
    .c(cout_8[51]),
    .cout(cout_8[52]),
    .sum(sum_8[52]));
  AL_FADD comp8_53 (
    .a(1'b0),
    .b(sum_7[53]),
    .c(cout_8[52]),
    .cout(cout_8[53]),
    .sum(sum_8[53]));
  AL_FADD comp8_54 (
    .a(1'b0),
    .b(sum_7[54]),
    .c(cout_8[53]),
    .cout(cout_8[54]),
    .sum(sum_8[54]));
  AL_FADD comp8_55 (
    .a(1'b0),
    .b(sum_7[55]),
    .c(cout_8[54]),
    .cout(cout_8[55]),
    .sum(sum_8[55]));
  AL_FADD comp8_56 (
    .a(1'b0),
    .b(sum_7[56]),
    .c(cout_8[55]),
    .cout(cout_8[56]),
    .sum(sum_8[56]));
  AL_FADD comp8_57 (
    .a(1'b0),
    .b(sum_7[57]),
    .c(cout_8[56]),
    .cout(cout_8[57]),
    .sum(sum_8[57]));
  AL_FADD comp8_58 (
    .a(1'b0),
    .b(sum_7[58]),
    .c(cout_8[57]),
    .cout(cout_8[58]),
    .sum(sum_8[58]));
  AL_FADD comp8_59 (
    .a(1'b0),
    .b(sum_7[59]),
    .c(cout_8[58]),
    .cout(cout_8[59]),
    .sum(sum_8[59]));
  AL_FADD comp8_6 (
    .a(i8[6]),
    .b(sum_7[6]),
    .c(cout_8[5]),
    .cout(cout_8[6]),
    .sum(sum_8[6]));
  AL_FADD comp8_60 (
    .a(1'b0),
    .b(sum_7[60]),
    .c(cout_8[59]),
    .cout(cout_8[60]),
    .sum(sum_8[60]));
  AL_FADD comp8_61 (
    .a(1'b0),
    .b(sum_7[61]),
    .c(cout_8[60]),
    .cout(cout_8[61]),
    .sum(sum_8[61]));
  AL_FADD comp8_62 (
    .a(1'b0),
    .b(sum_7[62]),
    .c(cout_8[61]),
    .cout(cout_8[62]),
    .sum(sum_8[62]));
  AL_FADD comp8_63 (
    .a(1'b0),
    .b(sum_7[63]),
    .c(cout_8[62]),
    .cout(cout_8[63]),
    .sum(sum_8[63]));
  AL_FADD comp8_7 (
    .a(i8[7]),
    .b(sum_7[7]),
    .c(cout_8[6]),
    .cout(cout_8[7]),
    .sum(sum_8[7]));
  AL_FADD comp8_8 (
    .a(i8[8]),
    .b(sum_7[8]),
    .c(cout_8[7]),
    .cout(cout_8[8]),
    .sum(sum_8[8]));
  AL_FADD comp8_9 (
    .a(i8[9]),
    .b(sum_7[9]),
    .c(cout_8[8]),
    .cout(cout_8[9]),
    .sum(sum_8[9]));
  AL_FADD comp9_0 (
    .a(i9[0]),
    .b(sum_8[0]),
    .c(1'b0),
    .cout(cout_9[0]),
    .sum(sum_9[0]));
  AL_FADD comp9_1 (
    .a(i9[1]),
    .b(sum_8[1]),
    .c(cout_9[0]),
    .cout(cout_9[1]),
    .sum(sum_9[1]));
  AL_FADD comp9_10 (
    .a(i9[10]),
    .b(sum_8[10]),
    .c(cout_9[9]),
    .cout(cout_9[10]),
    .sum(sum_9[10]));
  AL_FADD comp9_11 (
    .a(i9[11]),
    .b(sum_8[11]),
    .c(cout_9[10]),
    .cout(cout_9[11]),
    .sum(sum_9[11]));
  AL_FADD comp9_12 (
    .a(i9[12]),
    .b(sum_8[12]),
    .c(cout_9[11]),
    .cout(cout_9[12]),
    .sum(sum_9[12]));
  AL_FADD comp9_13 (
    .a(i9[13]),
    .b(sum_8[13]),
    .c(cout_9[12]),
    .cout(cout_9[13]),
    .sum(sum_9[13]));
  AL_FADD comp9_14 (
    .a(i9[14]),
    .b(sum_8[14]),
    .c(cout_9[13]),
    .cout(cout_9[14]),
    .sum(sum_9[14]));
  AL_FADD comp9_15 (
    .a(i9[15]),
    .b(sum_8[15]),
    .c(cout_9[14]),
    .cout(cout_9[15]),
    .sum(sum_9[15]));
  AL_FADD comp9_16 (
    .a(i9[16]),
    .b(sum_8[16]),
    .c(cout_9[15]),
    .cout(cout_9[16]),
    .sum(sum_9[16]));
  AL_FADD comp9_17 (
    .a(i9[17]),
    .b(sum_8[17]),
    .c(cout_9[16]),
    .cout(cout_9[17]),
    .sum(sum_9[17]));
  AL_FADD comp9_18 (
    .a(i9[18]),
    .b(sum_8[18]),
    .c(cout_9[17]),
    .cout(cout_9[18]),
    .sum(sum_9[18]));
  AL_FADD comp9_19 (
    .a(i9[19]),
    .b(sum_8[19]),
    .c(cout_9[18]),
    .cout(cout_9[19]),
    .sum(sum_9[19]));
  AL_FADD comp9_2 (
    .a(i9[2]),
    .b(sum_8[2]),
    .c(cout_9[1]),
    .cout(cout_9[2]),
    .sum(sum_9[2]));
  AL_FADD comp9_20 (
    .a(i9[20]),
    .b(sum_8[20]),
    .c(cout_9[19]),
    .cout(cout_9[20]),
    .sum(sum_9[20]));
  AL_FADD comp9_21 (
    .a(i9[21]),
    .b(sum_8[21]),
    .c(cout_9[20]),
    .cout(cout_9[21]),
    .sum(sum_9[21]));
  AL_FADD comp9_22 (
    .a(i9[22]),
    .b(sum_8[22]),
    .c(cout_9[21]),
    .cout(cout_9[22]),
    .sum(sum_9[22]));
  AL_FADD comp9_23 (
    .a(i9[23]),
    .b(sum_8[23]),
    .c(cout_9[22]),
    .cout(cout_9[23]),
    .sum(sum_9[23]));
  AL_FADD comp9_24 (
    .a(i9[24]),
    .b(sum_8[24]),
    .c(cout_9[23]),
    .cout(cout_9[24]),
    .sum(sum_9[24]));
  AL_FADD comp9_25 (
    .a(i9[25]),
    .b(sum_8[25]),
    .c(cout_9[24]),
    .cout(cout_9[25]),
    .sum(sum_9[25]));
  AL_FADD comp9_26 (
    .a(i9[26]),
    .b(sum_8[26]),
    .c(cout_9[25]),
    .cout(cout_9[26]),
    .sum(sum_9[26]));
  AL_FADD comp9_27 (
    .a(i9[27]),
    .b(sum_8[27]),
    .c(cout_9[26]),
    .cout(cout_9[27]),
    .sum(sum_9[27]));
  AL_FADD comp9_28 (
    .a(i9[28]),
    .b(sum_8[28]),
    .c(cout_9[27]),
    .cout(cout_9[28]),
    .sum(sum_9[28]));
  AL_FADD comp9_29 (
    .a(i9[29]),
    .b(sum_8[29]),
    .c(cout_9[28]),
    .cout(cout_9[29]),
    .sum(sum_9[29]));
  AL_FADD comp9_3 (
    .a(i9[3]),
    .b(sum_8[3]),
    .c(cout_9[2]),
    .cout(cout_9[3]),
    .sum(sum_9[3]));
  AL_FADD comp9_30 (
    .a(i9[30]),
    .b(sum_8[30]),
    .c(cout_9[29]),
    .cout(cout_9[30]),
    .sum(sum_9[30]));
  AL_FADD comp9_31 (
    .a(i9[31]),
    .b(sum_8[31]),
    .c(cout_9[30]),
    .cout(cout_9[31]),
    .sum(sum_9[31]));
  AL_FADD comp9_32 (
    .a(i9[32]),
    .b(sum_8[32]),
    .c(cout_9[31]),
    .cout(cout_9[32]),
    .sum(sum_9[32]));
  AL_FADD comp9_33 (
    .a(i9[33]),
    .b(sum_8[33]),
    .c(cout_9[32]),
    .cout(cout_9[33]),
    .sum(sum_9[33]));
  AL_FADD comp9_34 (
    .a(i9[34]),
    .b(sum_8[34]),
    .c(cout_9[33]),
    .cout(cout_9[34]),
    .sum(sum_9[34]));
  AL_FADD comp9_35 (
    .a(i9[35]),
    .b(sum_8[35]),
    .c(cout_9[34]),
    .cout(cout_9[35]),
    .sum(sum_9[35]));
  AL_FADD comp9_36 (
    .a(i9[36]),
    .b(sum_8[36]),
    .c(cout_9[35]),
    .cout(cout_9[36]),
    .sum(sum_9[36]));
  AL_FADD comp9_37 (
    .a(i9[37]),
    .b(sum_8[37]),
    .c(cout_9[36]),
    .cout(cout_9[37]),
    .sum(sum_9[37]));
  AL_FADD comp9_38 (
    .a(i9[38]),
    .b(sum_8[38]),
    .c(cout_9[37]),
    .cout(cout_9[38]),
    .sum(sum_9[38]));
  AL_FADD comp9_39 (
    .a(i9[39]),
    .b(sum_8[39]),
    .c(cout_9[38]),
    .cout(cout_9[39]),
    .sum(sum_9[39]));
  AL_FADD comp9_4 (
    .a(i9[4]),
    .b(sum_8[4]),
    .c(cout_9[3]),
    .cout(cout_9[4]),
    .sum(sum_9[4]));
  AL_FADD comp9_40 (
    .a(i9[40]),
    .b(sum_8[40]),
    .c(cout_9[39]),
    .cout(cout_9[40]),
    .sum(sum_9[40]));
  AL_FADD comp9_41 (
    .a(i9[41]),
    .b(sum_8[41]),
    .c(cout_9[40]),
    .cout(cout_9[41]),
    .sum(sum_9[41]));
  AL_FADD comp9_42 (
    .a(i9[42]),
    .b(sum_8[42]),
    .c(cout_9[41]),
    .cout(cout_9[42]),
    .sum(sum_9[42]));
  AL_FADD comp9_43 (
    .a(i9[43]),
    .b(sum_8[43]),
    .c(cout_9[42]),
    .cout(cout_9[43]),
    .sum(sum_9[43]));
  AL_FADD comp9_44 (
    .a(i9[44]),
    .b(sum_8[44]),
    .c(cout_9[43]),
    .cout(cout_9[44]),
    .sum(sum_9[44]));
  AL_FADD comp9_45 (
    .a(i9[45]),
    .b(sum_8[45]),
    .c(cout_9[44]),
    .cout(cout_9[45]),
    .sum(sum_9[45]));
  AL_FADD comp9_46 (
    .a(i9[46]),
    .b(sum_8[46]),
    .c(cout_9[45]),
    .cout(cout_9[46]),
    .sum(sum_9[46]));
  AL_FADD comp9_47 (
    .a(i9[47]),
    .b(sum_8[47]),
    .c(cout_9[46]),
    .cout(cout_9[47]),
    .sum(sum_9[47]));
  AL_FADD comp9_48 (
    .a(i9[48]),
    .b(sum_8[48]),
    .c(cout_9[47]),
    .cout(cout_9[48]),
    .sum(sum_9[48]));
  AL_FADD comp9_49 (
    .a(i9[49]),
    .b(sum_8[49]),
    .c(cout_9[48]),
    .cout(cout_9[49]),
    .sum(sum_9[49]));
  AL_FADD comp9_5 (
    .a(i9[5]),
    .b(sum_8[5]),
    .c(cout_9[4]),
    .cout(cout_9[5]),
    .sum(sum_9[5]));
  AL_FADD comp9_50 (
    .a(i9[50]),
    .b(sum_8[50]),
    .c(cout_9[49]),
    .cout(cout_9[50]),
    .sum(sum_9[50]));
  AL_FADD comp9_51 (
    .a(i9[51]),
    .b(sum_8[51]),
    .c(cout_9[50]),
    .cout(cout_9[51]),
    .sum(sum_9[51]));
  AL_FADD comp9_52 (
    .a(1'b0),
    .b(sum_8[52]),
    .c(cout_9[51]),
    .cout(cout_9[52]),
    .sum(sum_9[52]));
  AL_FADD comp9_53 (
    .a(1'b0),
    .b(sum_8[53]),
    .c(cout_9[52]),
    .cout(cout_9[53]),
    .sum(sum_9[53]));
  AL_FADD comp9_54 (
    .a(1'b0),
    .b(sum_8[54]),
    .c(cout_9[53]),
    .cout(cout_9[54]),
    .sum(sum_9[54]));
  AL_FADD comp9_55 (
    .a(1'b0),
    .b(sum_8[55]),
    .c(cout_9[54]),
    .cout(cout_9[55]),
    .sum(sum_9[55]));
  AL_FADD comp9_56 (
    .a(1'b0),
    .b(sum_8[56]),
    .c(cout_9[55]),
    .cout(cout_9[56]),
    .sum(sum_9[56]));
  AL_FADD comp9_57 (
    .a(1'b0),
    .b(sum_8[57]),
    .c(cout_9[56]),
    .cout(cout_9[57]),
    .sum(sum_9[57]));
  AL_FADD comp9_58 (
    .a(1'b0),
    .b(sum_8[58]),
    .c(cout_9[57]),
    .cout(cout_9[58]),
    .sum(sum_9[58]));
  AL_FADD comp9_59 (
    .a(1'b0),
    .b(sum_8[59]),
    .c(cout_9[58]),
    .cout(cout_9[59]),
    .sum(sum_9[59]));
  AL_FADD comp9_6 (
    .a(i9[6]),
    .b(sum_8[6]),
    .c(cout_9[5]),
    .cout(cout_9[6]),
    .sum(sum_9[6]));
  AL_FADD comp9_60 (
    .a(1'b0),
    .b(sum_8[60]),
    .c(cout_9[59]),
    .cout(cout_9[60]),
    .sum(sum_9[60]));
  AL_FADD comp9_61 (
    .a(1'b0),
    .b(sum_8[61]),
    .c(cout_9[60]),
    .cout(cout_9[61]),
    .sum(sum_9[61]));
  AL_FADD comp9_62 (
    .a(1'b0),
    .b(sum_8[62]),
    .c(cout_9[61]),
    .cout(cout_9[62]),
    .sum(sum_9[62]));
  AL_FADD comp9_63 (
    .a(1'b0),
    .b(sum_8[63]),
    .c(cout_9[62]),
    .cout(cout_9[63]),
    .sum(sum_9[63]));
  AL_FADD comp9_7 (
    .a(i9[7]),
    .b(sum_8[7]),
    .c(cout_9[6]),
    .cout(cout_9[7]),
    .sum(sum_9[7]));
  AL_FADD comp9_8 (
    .a(i9[8]),
    .b(sum_8[8]),
    .c(cout_9[7]),
    .cout(cout_9[8]),
    .sum(sum_9[8]));
  AL_FADD comp9_9 (
    .a(i9[9]),
    .b(sum_8[9]),
    .c(cout_9[8]),
    .cout(cout_9[9]),
    .sum(sum_9[9]));
  not inv_b31_0 (net_nb31_0, i31[0]);
  not inv_b31_1 (net_nb31_1, i31[1]);
  not inv_b31_10 (net_nb31_10, i31[10]);
  not inv_b31_11 (net_nb31_11, i31[11]);
  not inv_b31_12 (net_nb31_12, i31[12]);
  not inv_b31_13 (net_nb31_13, i31[13]);
  not inv_b31_14 (net_nb31_14, i31[14]);
  not inv_b31_15 (net_nb31_15, i31[15]);
  not inv_b31_16 (net_nb31_16, i31[16]);
  not inv_b31_17 (net_nb31_17, i31[17]);
  not inv_b31_18 (net_nb31_18, i31[18]);
  not inv_b31_19 (net_nb31_19, i31[19]);
  not inv_b31_2 (net_nb31_2, i31[2]);
  not inv_b31_20 (net_nb31_20, i31[20]);
  not inv_b31_21 (net_nb31_21, i31[21]);
  not inv_b31_22 (net_nb31_22, i31[22]);
  not inv_b31_23 (net_nb31_23, i31[23]);
  not inv_b31_24 (net_nb31_24, i31[24]);
  not inv_b31_25 (net_nb31_25, i31[25]);
  not inv_b31_26 (net_nb31_26, i31[26]);
  not inv_b31_27 (net_nb31_27, i31[27]);
  not inv_b31_28 (net_nb31_28, i31[28]);
  not inv_b31_29 (net_nb31_29, i31[29]);
  not inv_b31_3 (net_nb31_3, i31[3]);
  not inv_b31_30 (net_nb31_30, i31[30]);
  not inv_b31_31 (net_nb31_31, i31[31]);
  not inv_b31_32 (net_nb31_32, i31[32]);
  not inv_b31_33 (net_nb31_33, i31[33]);
  not inv_b31_34 (net_nb31_34, i31[34]);
  not inv_b31_35 (net_nb31_35, i31[35]);
  not inv_b31_36 (net_nb31_36, i31[36]);
  not inv_b31_37 (net_nb31_37, i31[37]);
  not inv_b31_38 (net_nb31_38, i31[38]);
  not inv_b31_39 (net_nb31_39, i31[39]);
  not inv_b31_4 (net_nb31_4, i31[4]);
  not inv_b31_40 (net_nb31_40, i31[40]);
  not inv_b31_41 (net_nb31_41, i31[41]);
  not inv_b31_42 (net_nb31_42, i31[42]);
  not inv_b31_43 (net_nb31_43, i31[43]);
  not inv_b31_44 (net_nb31_44, i31[44]);
  not inv_b31_45 (net_nb31_45, i31[45]);
  not inv_b31_46 (net_nb31_46, i31[46]);
  not inv_b31_47 (net_nb31_47, i31[47]);
  not inv_b31_48 (net_nb31_48, i31[48]);
  not inv_b31_49 (net_nb31_49, i31[49]);
  not inv_b31_5 (net_nb31_5, i31[5]);
  not inv_b31_50 (net_nb31_50, i31[50]);
  not inv_b31_51 (net_nb31_51, i31[51]);
  not inv_b31_52 (net_nb31_52, i31[52]);
  not inv_b31_53 (net_nb31_53, i31[53]);
  not inv_b31_54 (net_nb31_54, i31[54]);
  not inv_b31_55 (net_nb31_55, i31[55]);
  not inv_b31_56 (net_nb31_56, i31[56]);
  not inv_b31_57 (net_nb31_57, i31[57]);
  not inv_b31_58 (net_nb31_58, i31[58]);
  not inv_b31_59 (net_nb31_59, i31[59]);
  not inv_b31_6 (net_nb31_6, i31[6]);
  not inv_b31_60 (net_nb31_60, i31[60]);
  not inv_b31_61 (net_nb31_61, i31[61]);
  not inv_b31_62 (net_nb31_62, 1'b0);
  not inv_b31_63 (net_nb31_63, 1'b0);
  not inv_b31_7 (net_nb31_7, i31[7]);
  not inv_b31_8 (net_nb31_8, i31[8]);
  not inv_b31_9 (net_nb31_9, i31[9]);
  not inv_b32_0 (net_nb32_0, i32[0]);
  not inv_b32_1 (net_nb32_1, i32[1]);
  not inv_b32_10 (net_nb32_10, i32[10]);
  not inv_b32_11 (net_nb32_11, i32[11]);
  not inv_b32_12 (net_nb32_12, i32[12]);
  not inv_b32_13 (net_nb32_13, i32[13]);
  not inv_b32_14 (net_nb32_14, i32[14]);
  not inv_b32_15 (net_nb32_15, i32[15]);
  not inv_b32_16 (net_nb32_16, i32[16]);
  not inv_b32_17 (net_nb32_17, i32[17]);
  not inv_b32_18 (net_nb32_18, i32[18]);
  not inv_b32_19 (net_nb32_19, i32[19]);
  not inv_b32_2 (net_nb32_2, i32[2]);
  not inv_b32_20 (net_nb32_20, i32[20]);
  not inv_b32_21 (net_nb32_21, i32[21]);
  not inv_b32_22 (net_nb32_22, i32[22]);
  not inv_b32_23 (net_nb32_23, i32[23]);
  not inv_b32_24 (net_nb32_24, i32[24]);
  not inv_b32_25 (net_nb32_25, i32[25]);
  not inv_b32_26 (net_nb32_26, i32[26]);
  not inv_b32_27 (net_nb32_27, i32[27]);
  not inv_b32_28 (net_nb32_28, i32[28]);
  not inv_b32_29 (net_nb32_29, i32[29]);
  not inv_b32_3 (net_nb32_3, i32[3]);
  not inv_b32_30 (net_nb32_30, i32[30]);
  not inv_b32_31 (net_nb32_31, i32[31]);
  not inv_b32_32 (net_nb32_32, i32[32]);
  not inv_b32_33 (net_nb32_33, i32[33]);
  not inv_b32_34 (net_nb32_34, i32[34]);
  not inv_b32_35 (net_nb32_35, i32[35]);
  not inv_b32_36 (net_nb32_36, i32[36]);
  not inv_b32_37 (net_nb32_37, i32[37]);
  not inv_b32_38 (net_nb32_38, i32[38]);
  not inv_b32_39 (net_nb32_39, i32[39]);
  not inv_b32_4 (net_nb32_4, i32[4]);
  not inv_b32_40 (net_nb32_40, i32[40]);
  not inv_b32_41 (net_nb32_41, i32[41]);
  not inv_b32_42 (net_nb32_42, i32[42]);
  not inv_b32_43 (net_nb32_43, i32[43]);
  not inv_b32_44 (net_nb32_44, i32[44]);
  not inv_b32_45 (net_nb32_45, i32[45]);
  not inv_b32_46 (net_nb32_46, i32[46]);
  not inv_b32_47 (net_nb32_47, i32[47]);
  not inv_b32_48 (net_nb32_48, i32[48]);
  not inv_b32_49 (net_nb32_49, i32[49]);
  not inv_b32_5 (net_nb32_5, i32[5]);
  not inv_b32_50 (net_nb32_50, i32[50]);
  not inv_b32_51 (net_nb32_51, i32[51]);
  not inv_b32_52 (net_nb32_52, i32[52]);
  not inv_b32_53 (net_nb32_53, i32[53]);
  not inv_b32_54 (net_nb32_54, i32[54]);
  not inv_b32_55 (net_nb32_55, i32[55]);
  not inv_b32_56 (net_nb32_56, i32[56]);
  not inv_b32_57 (net_nb32_57, i32[57]);
  not inv_b32_58 (net_nb32_58, i32[58]);
  not inv_b32_59 (net_nb32_59, i32[59]);
  not inv_b32_6 (net_nb32_6, i32[6]);
  not inv_b32_60 (net_nb32_60, i32[60]);
  not inv_b32_61 (net_nb32_61, i32[61]);
  not inv_b32_62 (net_nb32_62, 1'b0);
  not inv_b32_63 (net_nb32_63, 1'b0);
  not inv_b32_7 (net_nb32_7, i32[7]);
  not inv_b32_8 (net_nb32_8, i32[8]);
  not inv_b32_9 (net_nb32_9, i32[9]);
  not inv_cout31_63 (net_ncout31_63, cout_31[63]);
  not inv_cout32_63 (net_ncout32_63, cout_32[63]);

endmodule 

module add_pu63_pu62_pu61_pu60_pu59_pu58_pu57_pu56_pu55_pu54_pu53_pu52_pu51_pu50_pu49_pu48_pu47_pu46_pu45_pu44_pu43_pu42_pu41_pu40_pu39_pu38_pu37_pu36_pu35_pu34_pu33_pu32_o64
  (
  i0,
  i1,
  i10,
  i11,
  i12,
  i13,
  i14,
  i15,
  i16,
  i17,
  i18,
  i19,
  i2,
  i20,
  i21,
  i22,
  i23,
  i24,
  i25,
  i26,
  i27,
  i28,
  i29,
  i3,
  i30,
  i31,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  o
  );

  input [62:0] i0;
  input [61:0] i1;
  input [52:0] i10;
  input [51:0] i11;
  input [50:0] i12;
  input [49:0] i13;
  input [48:0] i14;
  input [47:0] i15;
  input [46:0] i16;
  input [45:0] i17;
  input [44:0] i18;
  input [43:0] i19;
  input [60:0] i2;
  input [42:0] i20;
  input [41:0] i21;
  input [40:0] i22;
  input [39:0] i23;
  input [38:0] i24;
  input [37:0] i25;
  input [36:0] i26;
  input [35:0] i27;
  input [34:0] i28;
  input [33:0] i29;
  input [59:0] i3;
  input [32:0] i30;
  input [31:0] i31;
  input [58:0] i4;
  input [57:0] i5;
  input [56:0] i6;
  input [55:0] i7;
  input [54:0] i8;
  input [53:0] i9;
  output [63:0] o;

  wire [62:0] cout_1;
  wire [63:0] cout_10;
  wire [63:0] cout_11;
  wire [63:0] cout_12;
  wire [63:0] cout_13;
  wire [63:0] cout_14;
  wire [63:0] cout_15;
  wire [63:0] cout_16;
  wire [63:0] cout_17;
  wire [63:0] cout_18;
  wire [63:0] cout_19;
  wire [63:0] cout_2;
  wire [63:0] cout_20;
  wire [63:0] cout_21;
  wire [63:0] cout_22;
  wire [63:0] cout_23;
  wire [63:0] cout_24;
  wire [63:0] cout_25;
  wire [63:0] cout_26;
  wire [63:0] cout_27;
  wire [63:0] cout_28;
  wire [63:0] cout_29;
  wire [63:0] cout_3;
  wire [63:0] cout_30;
  wire [63:0] cout_31;
  wire [63:0] cout_4;
  wire [63:0] cout_5;
  wire [63:0] cout_6;
  wire [63:0] cout_7;
  wire [63:0] cout_8;
  wire [63:0] cout_9;
  wire [62:0] sum_1;
  wire [63:0] sum_10;
  wire [63:0] sum_11;
  wire [63:0] sum_12;
  wire [63:0] sum_13;
  wire [63:0] sum_14;
  wire [63:0] sum_15;
  wire [63:0] sum_16;
  wire [63:0] sum_17;
  wire [63:0] sum_18;
  wire [63:0] sum_19;
  wire [63:0] sum_2;
  wire [63:0] sum_20;
  wire [63:0] sum_21;
  wire [63:0] sum_22;
  wire [63:0] sum_23;
  wire [63:0] sum_24;
  wire [63:0] sum_25;
  wire [63:0] sum_26;
  wire [63:0] sum_27;
  wire [63:0] sum_28;
  wire [63:0] sum_29;
  wire [63:0] sum_3;
  wire [63:0] sum_30;
  wire [63:0] sum_31;
  wire [63:0] sum_4;
  wire [63:0] sum_5;
  wire [63:0] sum_6;
  wire [63:0] sum_7;
  wire [63:0] sum_8;
  wire [63:0] sum_9;

  assign o[63] = sum_31[63];
  assign o[62] = sum_31[62];
  assign o[61] = sum_31[61];
  assign o[60] = sum_31[60];
  assign o[59] = sum_31[59];
  assign o[58] = sum_31[58];
  assign o[57] = sum_31[57];
  assign o[56] = sum_31[56];
  assign o[55] = sum_31[55];
  assign o[54] = sum_31[54];
  assign o[53] = sum_31[53];
  assign o[52] = sum_31[52];
  assign o[51] = sum_31[51];
  assign o[50] = sum_31[50];
  assign o[49] = sum_31[49];
  assign o[48] = sum_31[48];
  assign o[47] = sum_31[47];
  assign o[46] = sum_31[46];
  assign o[45] = sum_31[45];
  assign o[44] = sum_31[44];
  assign o[43] = sum_31[43];
  assign o[42] = sum_31[42];
  assign o[41] = sum_31[41];
  assign o[40] = sum_31[40];
  assign o[39] = sum_31[39];
  assign o[38] = sum_31[38];
  assign o[37] = sum_31[37];
  assign o[36] = sum_31[36];
  assign o[35] = sum_31[35];
  assign o[34] = sum_31[34];
  assign o[33] = sum_31[33];
  assign o[32] = sum_31[32];
  assign o[31] = sum_31[31];
  assign o[30] = sum_31[30];
  assign o[29] = sum_31[29];
  assign o[28] = sum_31[28];
  assign o[27] = sum_31[27];
  assign o[26] = sum_31[26];
  assign o[25] = sum_31[25];
  assign o[24] = sum_31[24];
  assign o[23] = sum_31[23];
  assign o[22] = sum_31[22];
  assign o[21] = sum_31[21];
  assign o[20] = sum_31[20];
  assign o[19] = sum_31[19];
  assign o[18] = sum_31[18];
  assign o[17] = sum_31[17];
  assign o[16] = sum_31[16];
  assign o[15] = sum_31[15];
  assign o[14] = sum_31[14];
  assign o[13] = sum_31[13];
  assign o[12] = sum_31[12];
  assign o[11] = sum_31[11];
  assign o[10] = sum_31[10];
  assign o[9] = sum_31[9];
  assign o[8] = sum_31[8];
  assign o[7] = sum_31[7];
  assign o[6] = sum_31[6];
  assign o[5] = sum_31[5];
  assign o[4] = sum_31[4];
  assign o[3] = sum_31[3];
  assign o[2] = sum_31[2];
  assign o[1] = sum_31[1];
  assign o[0] = sum_31[0];
  AL_FADD comp10_0 (
    .a(i10[0]),
    .b(sum_9[0]),
    .c(1'b0),
    .cout(cout_10[0]),
    .sum(sum_10[0]));
  AL_FADD comp10_1 (
    .a(i10[1]),
    .b(sum_9[1]),
    .c(cout_10[0]),
    .cout(cout_10[1]),
    .sum(sum_10[1]));
  AL_FADD comp10_10 (
    .a(i10[10]),
    .b(sum_9[10]),
    .c(cout_10[9]),
    .cout(cout_10[10]),
    .sum(sum_10[10]));
  AL_FADD comp10_11 (
    .a(i10[11]),
    .b(sum_9[11]),
    .c(cout_10[10]),
    .cout(cout_10[11]),
    .sum(sum_10[11]));
  AL_FADD comp10_12 (
    .a(i10[12]),
    .b(sum_9[12]),
    .c(cout_10[11]),
    .cout(cout_10[12]),
    .sum(sum_10[12]));
  AL_FADD comp10_13 (
    .a(i10[13]),
    .b(sum_9[13]),
    .c(cout_10[12]),
    .cout(cout_10[13]),
    .sum(sum_10[13]));
  AL_FADD comp10_14 (
    .a(i10[14]),
    .b(sum_9[14]),
    .c(cout_10[13]),
    .cout(cout_10[14]),
    .sum(sum_10[14]));
  AL_FADD comp10_15 (
    .a(i10[15]),
    .b(sum_9[15]),
    .c(cout_10[14]),
    .cout(cout_10[15]),
    .sum(sum_10[15]));
  AL_FADD comp10_16 (
    .a(i10[16]),
    .b(sum_9[16]),
    .c(cout_10[15]),
    .cout(cout_10[16]),
    .sum(sum_10[16]));
  AL_FADD comp10_17 (
    .a(i10[17]),
    .b(sum_9[17]),
    .c(cout_10[16]),
    .cout(cout_10[17]),
    .sum(sum_10[17]));
  AL_FADD comp10_18 (
    .a(i10[18]),
    .b(sum_9[18]),
    .c(cout_10[17]),
    .cout(cout_10[18]),
    .sum(sum_10[18]));
  AL_FADD comp10_19 (
    .a(i10[19]),
    .b(sum_9[19]),
    .c(cout_10[18]),
    .cout(cout_10[19]),
    .sum(sum_10[19]));
  AL_FADD comp10_2 (
    .a(i10[2]),
    .b(sum_9[2]),
    .c(cout_10[1]),
    .cout(cout_10[2]),
    .sum(sum_10[2]));
  AL_FADD comp10_20 (
    .a(i10[20]),
    .b(sum_9[20]),
    .c(cout_10[19]),
    .cout(cout_10[20]),
    .sum(sum_10[20]));
  AL_FADD comp10_21 (
    .a(i10[21]),
    .b(sum_9[21]),
    .c(cout_10[20]),
    .cout(cout_10[21]),
    .sum(sum_10[21]));
  AL_FADD comp10_22 (
    .a(i10[22]),
    .b(sum_9[22]),
    .c(cout_10[21]),
    .cout(cout_10[22]),
    .sum(sum_10[22]));
  AL_FADD comp10_23 (
    .a(i10[23]),
    .b(sum_9[23]),
    .c(cout_10[22]),
    .cout(cout_10[23]),
    .sum(sum_10[23]));
  AL_FADD comp10_24 (
    .a(i10[24]),
    .b(sum_9[24]),
    .c(cout_10[23]),
    .cout(cout_10[24]),
    .sum(sum_10[24]));
  AL_FADD comp10_25 (
    .a(i10[25]),
    .b(sum_9[25]),
    .c(cout_10[24]),
    .cout(cout_10[25]),
    .sum(sum_10[25]));
  AL_FADD comp10_26 (
    .a(i10[26]),
    .b(sum_9[26]),
    .c(cout_10[25]),
    .cout(cout_10[26]),
    .sum(sum_10[26]));
  AL_FADD comp10_27 (
    .a(i10[27]),
    .b(sum_9[27]),
    .c(cout_10[26]),
    .cout(cout_10[27]),
    .sum(sum_10[27]));
  AL_FADD comp10_28 (
    .a(i10[28]),
    .b(sum_9[28]),
    .c(cout_10[27]),
    .cout(cout_10[28]),
    .sum(sum_10[28]));
  AL_FADD comp10_29 (
    .a(i10[29]),
    .b(sum_9[29]),
    .c(cout_10[28]),
    .cout(cout_10[29]),
    .sum(sum_10[29]));
  AL_FADD comp10_3 (
    .a(i10[3]),
    .b(sum_9[3]),
    .c(cout_10[2]),
    .cout(cout_10[3]),
    .sum(sum_10[3]));
  AL_FADD comp10_30 (
    .a(i10[30]),
    .b(sum_9[30]),
    .c(cout_10[29]),
    .cout(cout_10[30]),
    .sum(sum_10[30]));
  AL_FADD comp10_31 (
    .a(i10[31]),
    .b(sum_9[31]),
    .c(cout_10[30]),
    .cout(cout_10[31]),
    .sum(sum_10[31]));
  AL_FADD comp10_32 (
    .a(i10[32]),
    .b(sum_9[32]),
    .c(cout_10[31]),
    .cout(cout_10[32]),
    .sum(sum_10[32]));
  AL_FADD comp10_33 (
    .a(i10[33]),
    .b(sum_9[33]),
    .c(cout_10[32]),
    .cout(cout_10[33]),
    .sum(sum_10[33]));
  AL_FADD comp10_34 (
    .a(i10[34]),
    .b(sum_9[34]),
    .c(cout_10[33]),
    .cout(cout_10[34]),
    .sum(sum_10[34]));
  AL_FADD comp10_35 (
    .a(i10[35]),
    .b(sum_9[35]),
    .c(cout_10[34]),
    .cout(cout_10[35]),
    .sum(sum_10[35]));
  AL_FADD comp10_36 (
    .a(i10[36]),
    .b(sum_9[36]),
    .c(cout_10[35]),
    .cout(cout_10[36]),
    .sum(sum_10[36]));
  AL_FADD comp10_37 (
    .a(i10[37]),
    .b(sum_9[37]),
    .c(cout_10[36]),
    .cout(cout_10[37]),
    .sum(sum_10[37]));
  AL_FADD comp10_38 (
    .a(i10[38]),
    .b(sum_9[38]),
    .c(cout_10[37]),
    .cout(cout_10[38]),
    .sum(sum_10[38]));
  AL_FADD comp10_39 (
    .a(i10[39]),
    .b(sum_9[39]),
    .c(cout_10[38]),
    .cout(cout_10[39]),
    .sum(sum_10[39]));
  AL_FADD comp10_4 (
    .a(i10[4]),
    .b(sum_9[4]),
    .c(cout_10[3]),
    .cout(cout_10[4]),
    .sum(sum_10[4]));
  AL_FADD comp10_40 (
    .a(i10[40]),
    .b(sum_9[40]),
    .c(cout_10[39]),
    .cout(cout_10[40]),
    .sum(sum_10[40]));
  AL_FADD comp10_41 (
    .a(i10[41]),
    .b(sum_9[41]),
    .c(cout_10[40]),
    .cout(cout_10[41]),
    .sum(sum_10[41]));
  AL_FADD comp10_42 (
    .a(i10[42]),
    .b(sum_9[42]),
    .c(cout_10[41]),
    .cout(cout_10[42]),
    .sum(sum_10[42]));
  AL_FADD comp10_43 (
    .a(i10[43]),
    .b(sum_9[43]),
    .c(cout_10[42]),
    .cout(cout_10[43]),
    .sum(sum_10[43]));
  AL_FADD comp10_44 (
    .a(i10[44]),
    .b(sum_9[44]),
    .c(cout_10[43]),
    .cout(cout_10[44]),
    .sum(sum_10[44]));
  AL_FADD comp10_45 (
    .a(i10[45]),
    .b(sum_9[45]),
    .c(cout_10[44]),
    .cout(cout_10[45]),
    .sum(sum_10[45]));
  AL_FADD comp10_46 (
    .a(i10[46]),
    .b(sum_9[46]),
    .c(cout_10[45]),
    .cout(cout_10[46]),
    .sum(sum_10[46]));
  AL_FADD comp10_47 (
    .a(i10[47]),
    .b(sum_9[47]),
    .c(cout_10[46]),
    .cout(cout_10[47]),
    .sum(sum_10[47]));
  AL_FADD comp10_48 (
    .a(i10[48]),
    .b(sum_9[48]),
    .c(cout_10[47]),
    .cout(cout_10[48]),
    .sum(sum_10[48]));
  AL_FADD comp10_49 (
    .a(i10[49]),
    .b(sum_9[49]),
    .c(cout_10[48]),
    .cout(cout_10[49]),
    .sum(sum_10[49]));
  AL_FADD comp10_5 (
    .a(i10[5]),
    .b(sum_9[5]),
    .c(cout_10[4]),
    .cout(cout_10[5]),
    .sum(sum_10[5]));
  AL_FADD comp10_50 (
    .a(i10[50]),
    .b(sum_9[50]),
    .c(cout_10[49]),
    .cout(cout_10[50]),
    .sum(sum_10[50]));
  AL_FADD comp10_51 (
    .a(i10[51]),
    .b(sum_9[51]),
    .c(cout_10[50]),
    .cout(cout_10[51]),
    .sum(sum_10[51]));
  AL_FADD comp10_52 (
    .a(i10[52]),
    .b(sum_9[52]),
    .c(cout_10[51]),
    .cout(cout_10[52]),
    .sum(sum_10[52]));
  AL_FADD comp10_53 (
    .a(1'b0),
    .b(sum_9[53]),
    .c(cout_10[52]),
    .cout(cout_10[53]),
    .sum(sum_10[53]));
  AL_FADD comp10_54 (
    .a(1'b0),
    .b(sum_9[54]),
    .c(cout_10[53]),
    .cout(cout_10[54]),
    .sum(sum_10[54]));
  AL_FADD comp10_55 (
    .a(1'b0),
    .b(sum_9[55]),
    .c(cout_10[54]),
    .cout(cout_10[55]),
    .sum(sum_10[55]));
  AL_FADD comp10_56 (
    .a(1'b0),
    .b(sum_9[56]),
    .c(cout_10[55]),
    .cout(cout_10[56]),
    .sum(sum_10[56]));
  AL_FADD comp10_57 (
    .a(1'b0),
    .b(sum_9[57]),
    .c(cout_10[56]),
    .cout(cout_10[57]),
    .sum(sum_10[57]));
  AL_FADD comp10_58 (
    .a(1'b0),
    .b(sum_9[58]),
    .c(cout_10[57]),
    .cout(cout_10[58]),
    .sum(sum_10[58]));
  AL_FADD comp10_59 (
    .a(1'b0),
    .b(sum_9[59]),
    .c(cout_10[58]),
    .cout(cout_10[59]),
    .sum(sum_10[59]));
  AL_FADD comp10_6 (
    .a(i10[6]),
    .b(sum_9[6]),
    .c(cout_10[5]),
    .cout(cout_10[6]),
    .sum(sum_10[6]));
  AL_FADD comp10_60 (
    .a(1'b0),
    .b(sum_9[60]),
    .c(cout_10[59]),
    .cout(cout_10[60]),
    .sum(sum_10[60]));
  AL_FADD comp10_61 (
    .a(1'b0),
    .b(sum_9[61]),
    .c(cout_10[60]),
    .cout(cout_10[61]),
    .sum(sum_10[61]));
  AL_FADD comp10_62 (
    .a(1'b0),
    .b(sum_9[62]),
    .c(cout_10[61]),
    .cout(cout_10[62]),
    .sum(sum_10[62]));
  AL_FADD comp10_63 (
    .a(1'b0),
    .b(sum_9[63]),
    .c(cout_10[62]),
    .cout(cout_10[63]),
    .sum(sum_10[63]));
  AL_FADD comp10_7 (
    .a(i10[7]),
    .b(sum_9[7]),
    .c(cout_10[6]),
    .cout(cout_10[7]),
    .sum(sum_10[7]));
  AL_FADD comp10_8 (
    .a(i10[8]),
    .b(sum_9[8]),
    .c(cout_10[7]),
    .cout(cout_10[8]),
    .sum(sum_10[8]));
  AL_FADD comp10_9 (
    .a(i10[9]),
    .b(sum_9[9]),
    .c(cout_10[8]),
    .cout(cout_10[9]),
    .sum(sum_10[9]));
  AL_FADD comp11_0 (
    .a(i11[0]),
    .b(sum_10[0]),
    .c(1'b0),
    .cout(cout_11[0]),
    .sum(sum_11[0]));
  AL_FADD comp11_1 (
    .a(i11[1]),
    .b(sum_10[1]),
    .c(cout_11[0]),
    .cout(cout_11[1]),
    .sum(sum_11[1]));
  AL_FADD comp11_10 (
    .a(i11[10]),
    .b(sum_10[10]),
    .c(cout_11[9]),
    .cout(cout_11[10]),
    .sum(sum_11[10]));
  AL_FADD comp11_11 (
    .a(i11[11]),
    .b(sum_10[11]),
    .c(cout_11[10]),
    .cout(cout_11[11]),
    .sum(sum_11[11]));
  AL_FADD comp11_12 (
    .a(i11[12]),
    .b(sum_10[12]),
    .c(cout_11[11]),
    .cout(cout_11[12]),
    .sum(sum_11[12]));
  AL_FADD comp11_13 (
    .a(i11[13]),
    .b(sum_10[13]),
    .c(cout_11[12]),
    .cout(cout_11[13]),
    .sum(sum_11[13]));
  AL_FADD comp11_14 (
    .a(i11[14]),
    .b(sum_10[14]),
    .c(cout_11[13]),
    .cout(cout_11[14]),
    .sum(sum_11[14]));
  AL_FADD comp11_15 (
    .a(i11[15]),
    .b(sum_10[15]),
    .c(cout_11[14]),
    .cout(cout_11[15]),
    .sum(sum_11[15]));
  AL_FADD comp11_16 (
    .a(i11[16]),
    .b(sum_10[16]),
    .c(cout_11[15]),
    .cout(cout_11[16]),
    .sum(sum_11[16]));
  AL_FADD comp11_17 (
    .a(i11[17]),
    .b(sum_10[17]),
    .c(cout_11[16]),
    .cout(cout_11[17]),
    .sum(sum_11[17]));
  AL_FADD comp11_18 (
    .a(i11[18]),
    .b(sum_10[18]),
    .c(cout_11[17]),
    .cout(cout_11[18]),
    .sum(sum_11[18]));
  AL_FADD comp11_19 (
    .a(i11[19]),
    .b(sum_10[19]),
    .c(cout_11[18]),
    .cout(cout_11[19]),
    .sum(sum_11[19]));
  AL_FADD comp11_2 (
    .a(i11[2]),
    .b(sum_10[2]),
    .c(cout_11[1]),
    .cout(cout_11[2]),
    .sum(sum_11[2]));
  AL_FADD comp11_20 (
    .a(i11[20]),
    .b(sum_10[20]),
    .c(cout_11[19]),
    .cout(cout_11[20]),
    .sum(sum_11[20]));
  AL_FADD comp11_21 (
    .a(i11[21]),
    .b(sum_10[21]),
    .c(cout_11[20]),
    .cout(cout_11[21]),
    .sum(sum_11[21]));
  AL_FADD comp11_22 (
    .a(i11[22]),
    .b(sum_10[22]),
    .c(cout_11[21]),
    .cout(cout_11[22]),
    .sum(sum_11[22]));
  AL_FADD comp11_23 (
    .a(i11[23]),
    .b(sum_10[23]),
    .c(cout_11[22]),
    .cout(cout_11[23]),
    .sum(sum_11[23]));
  AL_FADD comp11_24 (
    .a(i11[24]),
    .b(sum_10[24]),
    .c(cout_11[23]),
    .cout(cout_11[24]),
    .sum(sum_11[24]));
  AL_FADD comp11_25 (
    .a(i11[25]),
    .b(sum_10[25]),
    .c(cout_11[24]),
    .cout(cout_11[25]),
    .sum(sum_11[25]));
  AL_FADD comp11_26 (
    .a(i11[26]),
    .b(sum_10[26]),
    .c(cout_11[25]),
    .cout(cout_11[26]),
    .sum(sum_11[26]));
  AL_FADD comp11_27 (
    .a(i11[27]),
    .b(sum_10[27]),
    .c(cout_11[26]),
    .cout(cout_11[27]),
    .sum(sum_11[27]));
  AL_FADD comp11_28 (
    .a(i11[28]),
    .b(sum_10[28]),
    .c(cout_11[27]),
    .cout(cout_11[28]),
    .sum(sum_11[28]));
  AL_FADD comp11_29 (
    .a(i11[29]),
    .b(sum_10[29]),
    .c(cout_11[28]),
    .cout(cout_11[29]),
    .sum(sum_11[29]));
  AL_FADD comp11_3 (
    .a(i11[3]),
    .b(sum_10[3]),
    .c(cout_11[2]),
    .cout(cout_11[3]),
    .sum(sum_11[3]));
  AL_FADD comp11_30 (
    .a(i11[30]),
    .b(sum_10[30]),
    .c(cout_11[29]),
    .cout(cout_11[30]),
    .sum(sum_11[30]));
  AL_FADD comp11_31 (
    .a(i11[31]),
    .b(sum_10[31]),
    .c(cout_11[30]),
    .cout(cout_11[31]),
    .sum(sum_11[31]));
  AL_FADD comp11_32 (
    .a(i11[32]),
    .b(sum_10[32]),
    .c(cout_11[31]),
    .cout(cout_11[32]),
    .sum(sum_11[32]));
  AL_FADD comp11_33 (
    .a(i11[33]),
    .b(sum_10[33]),
    .c(cout_11[32]),
    .cout(cout_11[33]),
    .sum(sum_11[33]));
  AL_FADD comp11_34 (
    .a(i11[34]),
    .b(sum_10[34]),
    .c(cout_11[33]),
    .cout(cout_11[34]),
    .sum(sum_11[34]));
  AL_FADD comp11_35 (
    .a(i11[35]),
    .b(sum_10[35]),
    .c(cout_11[34]),
    .cout(cout_11[35]),
    .sum(sum_11[35]));
  AL_FADD comp11_36 (
    .a(i11[36]),
    .b(sum_10[36]),
    .c(cout_11[35]),
    .cout(cout_11[36]),
    .sum(sum_11[36]));
  AL_FADD comp11_37 (
    .a(i11[37]),
    .b(sum_10[37]),
    .c(cout_11[36]),
    .cout(cout_11[37]),
    .sum(sum_11[37]));
  AL_FADD comp11_38 (
    .a(i11[38]),
    .b(sum_10[38]),
    .c(cout_11[37]),
    .cout(cout_11[38]),
    .sum(sum_11[38]));
  AL_FADD comp11_39 (
    .a(i11[39]),
    .b(sum_10[39]),
    .c(cout_11[38]),
    .cout(cout_11[39]),
    .sum(sum_11[39]));
  AL_FADD comp11_4 (
    .a(i11[4]),
    .b(sum_10[4]),
    .c(cout_11[3]),
    .cout(cout_11[4]),
    .sum(sum_11[4]));
  AL_FADD comp11_40 (
    .a(i11[40]),
    .b(sum_10[40]),
    .c(cout_11[39]),
    .cout(cout_11[40]),
    .sum(sum_11[40]));
  AL_FADD comp11_41 (
    .a(i11[41]),
    .b(sum_10[41]),
    .c(cout_11[40]),
    .cout(cout_11[41]),
    .sum(sum_11[41]));
  AL_FADD comp11_42 (
    .a(i11[42]),
    .b(sum_10[42]),
    .c(cout_11[41]),
    .cout(cout_11[42]),
    .sum(sum_11[42]));
  AL_FADD comp11_43 (
    .a(i11[43]),
    .b(sum_10[43]),
    .c(cout_11[42]),
    .cout(cout_11[43]),
    .sum(sum_11[43]));
  AL_FADD comp11_44 (
    .a(i11[44]),
    .b(sum_10[44]),
    .c(cout_11[43]),
    .cout(cout_11[44]),
    .sum(sum_11[44]));
  AL_FADD comp11_45 (
    .a(i11[45]),
    .b(sum_10[45]),
    .c(cout_11[44]),
    .cout(cout_11[45]),
    .sum(sum_11[45]));
  AL_FADD comp11_46 (
    .a(i11[46]),
    .b(sum_10[46]),
    .c(cout_11[45]),
    .cout(cout_11[46]),
    .sum(sum_11[46]));
  AL_FADD comp11_47 (
    .a(i11[47]),
    .b(sum_10[47]),
    .c(cout_11[46]),
    .cout(cout_11[47]),
    .sum(sum_11[47]));
  AL_FADD comp11_48 (
    .a(i11[48]),
    .b(sum_10[48]),
    .c(cout_11[47]),
    .cout(cout_11[48]),
    .sum(sum_11[48]));
  AL_FADD comp11_49 (
    .a(i11[49]),
    .b(sum_10[49]),
    .c(cout_11[48]),
    .cout(cout_11[49]),
    .sum(sum_11[49]));
  AL_FADD comp11_5 (
    .a(i11[5]),
    .b(sum_10[5]),
    .c(cout_11[4]),
    .cout(cout_11[5]),
    .sum(sum_11[5]));
  AL_FADD comp11_50 (
    .a(i11[50]),
    .b(sum_10[50]),
    .c(cout_11[49]),
    .cout(cout_11[50]),
    .sum(sum_11[50]));
  AL_FADD comp11_51 (
    .a(i11[51]),
    .b(sum_10[51]),
    .c(cout_11[50]),
    .cout(cout_11[51]),
    .sum(sum_11[51]));
  AL_FADD comp11_52 (
    .a(1'b0),
    .b(sum_10[52]),
    .c(cout_11[51]),
    .cout(cout_11[52]),
    .sum(sum_11[52]));
  AL_FADD comp11_53 (
    .a(1'b0),
    .b(sum_10[53]),
    .c(cout_11[52]),
    .cout(cout_11[53]),
    .sum(sum_11[53]));
  AL_FADD comp11_54 (
    .a(1'b0),
    .b(sum_10[54]),
    .c(cout_11[53]),
    .cout(cout_11[54]),
    .sum(sum_11[54]));
  AL_FADD comp11_55 (
    .a(1'b0),
    .b(sum_10[55]),
    .c(cout_11[54]),
    .cout(cout_11[55]),
    .sum(sum_11[55]));
  AL_FADD comp11_56 (
    .a(1'b0),
    .b(sum_10[56]),
    .c(cout_11[55]),
    .cout(cout_11[56]),
    .sum(sum_11[56]));
  AL_FADD comp11_57 (
    .a(1'b0),
    .b(sum_10[57]),
    .c(cout_11[56]),
    .cout(cout_11[57]),
    .sum(sum_11[57]));
  AL_FADD comp11_58 (
    .a(1'b0),
    .b(sum_10[58]),
    .c(cout_11[57]),
    .cout(cout_11[58]),
    .sum(sum_11[58]));
  AL_FADD comp11_59 (
    .a(1'b0),
    .b(sum_10[59]),
    .c(cout_11[58]),
    .cout(cout_11[59]),
    .sum(sum_11[59]));
  AL_FADD comp11_6 (
    .a(i11[6]),
    .b(sum_10[6]),
    .c(cout_11[5]),
    .cout(cout_11[6]),
    .sum(sum_11[6]));
  AL_FADD comp11_60 (
    .a(1'b0),
    .b(sum_10[60]),
    .c(cout_11[59]),
    .cout(cout_11[60]),
    .sum(sum_11[60]));
  AL_FADD comp11_61 (
    .a(1'b0),
    .b(sum_10[61]),
    .c(cout_11[60]),
    .cout(cout_11[61]),
    .sum(sum_11[61]));
  AL_FADD comp11_62 (
    .a(1'b0),
    .b(sum_10[62]),
    .c(cout_11[61]),
    .cout(cout_11[62]),
    .sum(sum_11[62]));
  AL_FADD comp11_63 (
    .a(1'b0),
    .b(sum_10[63]),
    .c(cout_11[62]),
    .cout(cout_11[63]),
    .sum(sum_11[63]));
  AL_FADD comp11_7 (
    .a(i11[7]),
    .b(sum_10[7]),
    .c(cout_11[6]),
    .cout(cout_11[7]),
    .sum(sum_11[7]));
  AL_FADD comp11_8 (
    .a(i11[8]),
    .b(sum_10[8]),
    .c(cout_11[7]),
    .cout(cout_11[8]),
    .sum(sum_11[8]));
  AL_FADD comp11_9 (
    .a(i11[9]),
    .b(sum_10[9]),
    .c(cout_11[8]),
    .cout(cout_11[9]),
    .sum(sum_11[9]));
  AL_FADD comp12_0 (
    .a(i12[0]),
    .b(sum_11[0]),
    .c(1'b0),
    .cout(cout_12[0]),
    .sum(sum_12[0]));
  AL_FADD comp12_1 (
    .a(i12[1]),
    .b(sum_11[1]),
    .c(cout_12[0]),
    .cout(cout_12[1]),
    .sum(sum_12[1]));
  AL_FADD comp12_10 (
    .a(i12[10]),
    .b(sum_11[10]),
    .c(cout_12[9]),
    .cout(cout_12[10]),
    .sum(sum_12[10]));
  AL_FADD comp12_11 (
    .a(i12[11]),
    .b(sum_11[11]),
    .c(cout_12[10]),
    .cout(cout_12[11]),
    .sum(sum_12[11]));
  AL_FADD comp12_12 (
    .a(i12[12]),
    .b(sum_11[12]),
    .c(cout_12[11]),
    .cout(cout_12[12]),
    .sum(sum_12[12]));
  AL_FADD comp12_13 (
    .a(i12[13]),
    .b(sum_11[13]),
    .c(cout_12[12]),
    .cout(cout_12[13]),
    .sum(sum_12[13]));
  AL_FADD comp12_14 (
    .a(i12[14]),
    .b(sum_11[14]),
    .c(cout_12[13]),
    .cout(cout_12[14]),
    .sum(sum_12[14]));
  AL_FADD comp12_15 (
    .a(i12[15]),
    .b(sum_11[15]),
    .c(cout_12[14]),
    .cout(cout_12[15]),
    .sum(sum_12[15]));
  AL_FADD comp12_16 (
    .a(i12[16]),
    .b(sum_11[16]),
    .c(cout_12[15]),
    .cout(cout_12[16]),
    .sum(sum_12[16]));
  AL_FADD comp12_17 (
    .a(i12[17]),
    .b(sum_11[17]),
    .c(cout_12[16]),
    .cout(cout_12[17]),
    .sum(sum_12[17]));
  AL_FADD comp12_18 (
    .a(i12[18]),
    .b(sum_11[18]),
    .c(cout_12[17]),
    .cout(cout_12[18]),
    .sum(sum_12[18]));
  AL_FADD comp12_19 (
    .a(i12[19]),
    .b(sum_11[19]),
    .c(cout_12[18]),
    .cout(cout_12[19]),
    .sum(sum_12[19]));
  AL_FADD comp12_2 (
    .a(i12[2]),
    .b(sum_11[2]),
    .c(cout_12[1]),
    .cout(cout_12[2]),
    .sum(sum_12[2]));
  AL_FADD comp12_20 (
    .a(i12[20]),
    .b(sum_11[20]),
    .c(cout_12[19]),
    .cout(cout_12[20]),
    .sum(sum_12[20]));
  AL_FADD comp12_21 (
    .a(i12[21]),
    .b(sum_11[21]),
    .c(cout_12[20]),
    .cout(cout_12[21]),
    .sum(sum_12[21]));
  AL_FADD comp12_22 (
    .a(i12[22]),
    .b(sum_11[22]),
    .c(cout_12[21]),
    .cout(cout_12[22]),
    .sum(sum_12[22]));
  AL_FADD comp12_23 (
    .a(i12[23]),
    .b(sum_11[23]),
    .c(cout_12[22]),
    .cout(cout_12[23]),
    .sum(sum_12[23]));
  AL_FADD comp12_24 (
    .a(i12[24]),
    .b(sum_11[24]),
    .c(cout_12[23]),
    .cout(cout_12[24]),
    .sum(sum_12[24]));
  AL_FADD comp12_25 (
    .a(i12[25]),
    .b(sum_11[25]),
    .c(cout_12[24]),
    .cout(cout_12[25]),
    .sum(sum_12[25]));
  AL_FADD comp12_26 (
    .a(i12[26]),
    .b(sum_11[26]),
    .c(cout_12[25]),
    .cout(cout_12[26]),
    .sum(sum_12[26]));
  AL_FADD comp12_27 (
    .a(i12[27]),
    .b(sum_11[27]),
    .c(cout_12[26]),
    .cout(cout_12[27]),
    .sum(sum_12[27]));
  AL_FADD comp12_28 (
    .a(i12[28]),
    .b(sum_11[28]),
    .c(cout_12[27]),
    .cout(cout_12[28]),
    .sum(sum_12[28]));
  AL_FADD comp12_29 (
    .a(i12[29]),
    .b(sum_11[29]),
    .c(cout_12[28]),
    .cout(cout_12[29]),
    .sum(sum_12[29]));
  AL_FADD comp12_3 (
    .a(i12[3]),
    .b(sum_11[3]),
    .c(cout_12[2]),
    .cout(cout_12[3]),
    .sum(sum_12[3]));
  AL_FADD comp12_30 (
    .a(i12[30]),
    .b(sum_11[30]),
    .c(cout_12[29]),
    .cout(cout_12[30]),
    .sum(sum_12[30]));
  AL_FADD comp12_31 (
    .a(i12[31]),
    .b(sum_11[31]),
    .c(cout_12[30]),
    .cout(cout_12[31]),
    .sum(sum_12[31]));
  AL_FADD comp12_32 (
    .a(i12[32]),
    .b(sum_11[32]),
    .c(cout_12[31]),
    .cout(cout_12[32]),
    .sum(sum_12[32]));
  AL_FADD comp12_33 (
    .a(i12[33]),
    .b(sum_11[33]),
    .c(cout_12[32]),
    .cout(cout_12[33]),
    .sum(sum_12[33]));
  AL_FADD comp12_34 (
    .a(i12[34]),
    .b(sum_11[34]),
    .c(cout_12[33]),
    .cout(cout_12[34]),
    .sum(sum_12[34]));
  AL_FADD comp12_35 (
    .a(i12[35]),
    .b(sum_11[35]),
    .c(cout_12[34]),
    .cout(cout_12[35]),
    .sum(sum_12[35]));
  AL_FADD comp12_36 (
    .a(i12[36]),
    .b(sum_11[36]),
    .c(cout_12[35]),
    .cout(cout_12[36]),
    .sum(sum_12[36]));
  AL_FADD comp12_37 (
    .a(i12[37]),
    .b(sum_11[37]),
    .c(cout_12[36]),
    .cout(cout_12[37]),
    .sum(sum_12[37]));
  AL_FADD comp12_38 (
    .a(i12[38]),
    .b(sum_11[38]),
    .c(cout_12[37]),
    .cout(cout_12[38]),
    .sum(sum_12[38]));
  AL_FADD comp12_39 (
    .a(i12[39]),
    .b(sum_11[39]),
    .c(cout_12[38]),
    .cout(cout_12[39]),
    .sum(sum_12[39]));
  AL_FADD comp12_4 (
    .a(i12[4]),
    .b(sum_11[4]),
    .c(cout_12[3]),
    .cout(cout_12[4]),
    .sum(sum_12[4]));
  AL_FADD comp12_40 (
    .a(i12[40]),
    .b(sum_11[40]),
    .c(cout_12[39]),
    .cout(cout_12[40]),
    .sum(sum_12[40]));
  AL_FADD comp12_41 (
    .a(i12[41]),
    .b(sum_11[41]),
    .c(cout_12[40]),
    .cout(cout_12[41]),
    .sum(sum_12[41]));
  AL_FADD comp12_42 (
    .a(i12[42]),
    .b(sum_11[42]),
    .c(cout_12[41]),
    .cout(cout_12[42]),
    .sum(sum_12[42]));
  AL_FADD comp12_43 (
    .a(i12[43]),
    .b(sum_11[43]),
    .c(cout_12[42]),
    .cout(cout_12[43]),
    .sum(sum_12[43]));
  AL_FADD comp12_44 (
    .a(i12[44]),
    .b(sum_11[44]),
    .c(cout_12[43]),
    .cout(cout_12[44]),
    .sum(sum_12[44]));
  AL_FADD comp12_45 (
    .a(i12[45]),
    .b(sum_11[45]),
    .c(cout_12[44]),
    .cout(cout_12[45]),
    .sum(sum_12[45]));
  AL_FADD comp12_46 (
    .a(i12[46]),
    .b(sum_11[46]),
    .c(cout_12[45]),
    .cout(cout_12[46]),
    .sum(sum_12[46]));
  AL_FADD comp12_47 (
    .a(i12[47]),
    .b(sum_11[47]),
    .c(cout_12[46]),
    .cout(cout_12[47]),
    .sum(sum_12[47]));
  AL_FADD comp12_48 (
    .a(i12[48]),
    .b(sum_11[48]),
    .c(cout_12[47]),
    .cout(cout_12[48]),
    .sum(sum_12[48]));
  AL_FADD comp12_49 (
    .a(i12[49]),
    .b(sum_11[49]),
    .c(cout_12[48]),
    .cout(cout_12[49]),
    .sum(sum_12[49]));
  AL_FADD comp12_5 (
    .a(i12[5]),
    .b(sum_11[5]),
    .c(cout_12[4]),
    .cout(cout_12[5]),
    .sum(sum_12[5]));
  AL_FADD comp12_50 (
    .a(i12[50]),
    .b(sum_11[50]),
    .c(cout_12[49]),
    .cout(cout_12[50]),
    .sum(sum_12[50]));
  AL_FADD comp12_51 (
    .a(1'b0),
    .b(sum_11[51]),
    .c(cout_12[50]),
    .cout(cout_12[51]),
    .sum(sum_12[51]));
  AL_FADD comp12_52 (
    .a(1'b0),
    .b(sum_11[52]),
    .c(cout_12[51]),
    .cout(cout_12[52]),
    .sum(sum_12[52]));
  AL_FADD comp12_53 (
    .a(1'b0),
    .b(sum_11[53]),
    .c(cout_12[52]),
    .cout(cout_12[53]),
    .sum(sum_12[53]));
  AL_FADD comp12_54 (
    .a(1'b0),
    .b(sum_11[54]),
    .c(cout_12[53]),
    .cout(cout_12[54]),
    .sum(sum_12[54]));
  AL_FADD comp12_55 (
    .a(1'b0),
    .b(sum_11[55]),
    .c(cout_12[54]),
    .cout(cout_12[55]),
    .sum(sum_12[55]));
  AL_FADD comp12_56 (
    .a(1'b0),
    .b(sum_11[56]),
    .c(cout_12[55]),
    .cout(cout_12[56]),
    .sum(sum_12[56]));
  AL_FADD comp12_57 (
    .a(1'b0),
    .b(sum_11[57]),
    .c(cout_12[56]),
    .cout(cout_12[57]),
    .sum(sum_12[57]));
  AL_FADD comp12_58 (
    .a(1'b0),
    .b(sum_11[58]),
    .c(cout_12[57]),
    .cout(cout_12[58]),
    .sum(sum_12[58]));
  AL_FADD comp12_59 (
    .a(1'b0),
    .b(sum_11[59]),
    .c(cout_12[58]),
    .cout(cout_12[59]),
    .sum(sum_12[59]));
  AL_FADD comp12_6 (
    .a(i12[6]),
    .b(sum_11[6]),
    .c(cout_12[5]),
    .cout(cout_12[6]),
    .sum(sum_12[6]));
  AL_FADD comp12_60 (
    .a(1'b0),
    .b(sum_11[60]),
    .c(cout_12[59]),
    .cout(cout_12[60]),
    .sum(sum_12[60]));
  AL_FADD comp12_61 (
    .a(1'b0),
    .b(sum_11[61]),
    .c(cout_12[60]),
    .cout(cout_12[61]),
    .sum(sum_12[61]));
  AL_FADD comp12_62 (
    .a(1'b0),
    .b(sum_11[62]),
    .c(cout_12[61]),
    .cout(cout_12[62]),
    .sum(sum_12[62]));
  AL_FADD comp12_63 (
    .a(1'b0),
    .b(sum_11[63]),
    .c(cout_12[62]),
    .cout(cout_12[63]),
    .sum(sum_12[63]));
  AL_FADD comp12_7 (
    .a(i12[7]),
    .b(sum_11[7]),
    .c(cout_12[6]),
    .cout(cout_12[7]),
    .sum(sum_12[7]));
  AL_FADD comp12_8 (
    .a(i12[8]),
    .b(sum_11[8]),
    .c(cout_12[7]),
    .cout(cout_12[8]),
    .sum(sum_12[8]));
  AL_FADD comp12_9 (
    .a(i12[9]),
    .b(sum_11[9]),
    .c(cout_12[8]),
    .cout(cout_12[9]),
    .sum(sum_12[9]));
  AL_FADD comp13_0 (
    .a(i13[0]),
    .b(sum_12[0]),
    .c(1'b0),
    .cout(cout_13[0]),
    .sum(sum_13[0]));
  AL_FADD comp13_1 (
    .a(i13[1]),
    .b(sum_12[1]),
    .c(cout_13[0]),
    .cout(cout_13[1]),
    .sum(sum_13[1]));
  AL_FADD comp13_10 (
    .a(i13[10]),
    .b(sum_12[10]),
    .c(cout_13[9]),
    .cout(cout_13[10]),
    .sum(sum_13[10]));
  AL_FADD comp13_11 (
    .a(i13[11]),
    .b(sum_12[11]),
    .c(cout_13[10]),
    .cout(cout_13[11]),
    .sum(sum_13[11]));
  AL_FADD comp13_12 (
    .a(i13[12]),
    .b(sum_12[12]),
    .c(cout_13[11]),
    .cout(cout_13[12]),
    .sum(sum_13[12]));
  AL_FADD comp13_13 (
    .a(i13[13]),
    .b(sum_12[13]),
    .c(cout_13[12]),
    .cout(cout_13[13]),
    .sum(sum_13[13]));
  AL_FADD comp13_14 (
    .a(i13[14]),
    .b(sum_12[14]),
    .c(cout_13[13]),
    .cout(cout_13[14]),
    .sum(sum_13[14]));
  AL_FADD comp13_15 (
    .a(i13[15]),
    .b(sum_12[15]),
    .c(cout_13[14]),
    .cout(cout_13[15]),
    .sum(sum_13[15]));
  AL_FADD comp13_16 (
    .a(i13[16]),
    .b(sum_12[16]),
    .c(cout_13[15]),
    .cout(cout_13[16]),
    .sum(sum_13[16]));
  AL_FADD comp13_17 (
    .a(i13[17]),
    .b(sum_12[17]),
    .c(cout_13[16]),
    .cout(cout_13[17]),
    .sum(sum_13[17]));
  AL_FADD comp13_18 (
    .a(i13[18]),
    .b(sum_12[18]),
    .c(cout_13[17]),
    .cout(cout_13[18]),
    .sum(sum_13[18]));
  AL_FADD comp13_19 (
    .a(i13[19]),
    .b(sum_12[19]),
    .c(cout_13[18]),
    .cout(cout_13[19]),
    .sum(sum_13[19]));
  AL_FADD comp13_2 (
    .a(i13[2]),
    .b(sum_12[2]),
    .c(cout_13[1]),
    .cout(cout_13[2]),
    .sum(sum_13[2]));
  AL_FADD comp13_20 (
    .a(i13[20]),
    .b(sum_12[20]),
    .c(cout_13[19]),
    .cout(cout_13[20]),
    .sum(sum_13[20]));
  AL_FADD comp13_21 (
    .a(i13[21]),
    .b(sum_12[21]),
    .c(cout_13[20]),
    .cout(cout_13[21]),
    .sum(sum_13[21]));
  AL_FADD comp13_22 (
    .a(i13[22]),
    .b(sum_12[22]),
    .c(cout_13[21]),
    .cout(cout_13[22]),
    .sum(sum_13[22]));
  AL_FADD comp13_23 (
    .a(i13[23]),
    .b(sum_12[23]),
    .c(cout_13[22]),
    .cout(cout_13[23]),
    .sum(sum_13[23]));
  AL_FADD comp13_24 (
    .a(i13[24]),
    .b(sum_12[24]),
    .c(cout_13[23]),
    .cout(cout_13[24]),
    .sum(sum_13[24]));
  AL_FADD comp13_25 (
    .a(i13[25]),
    .b(sum_12[25]),
    .c(cout_13[24]),
    .cout(cout_13[25]),
    .sum(sum_13[25]));
  AL_FADD comp13_26 (
    .a(i13[26]),
    .b(sum_12[26]),
    .c(cout_13[25]),
    .cout(cout_13[26]),
    .sum(sum_13[26]));
  AL_FADD comp13_27 (
    .a(i13[27]),
    .b(sum_12[27]),
    .c(cout_13[26]),
    .cout(cout_13[27]),
    .sum(sum_13[27]));
  AL_FADD comp13_28 (
    .a(i13[28]),
    .b(sum_12[28]),
    .c(cout_13[27]),
    .cout(cout_13[28]),
    .sum(sum_13[28]));
  AL_FADD comp13_29 (
    .a(i13[29]),
    .b(sum_12[29]),
    .c(cout_13[28]),
    .cout(cout_13[29]),
    .sum(sum_13[29]));
  AL_FADD comp13_3 (
    .a(i13[3]),
    .b(sum_12[3]),
    .c(cout_13[2]),
    .cout(cout_13[3]),
    .sum(sum_13[3]));
  AL_FADD comp13_30 (
    .a(i13[30]),
    .b(sum_12[30]),
    .c(cout_13[29]),
    .cout(cout_13[30]),
    .sum(sum_13[30]));
  AL_FADD comp13_31 (
    .a(i13[31]),
    .b(sum_12[31]),
    .c(cout_13[30]),
    .cout(cout_13[31]),
    .sum(sum_13[31]));
  AL_FADD comp13_32 (
    .a(i13[32]),
    .b(sum_12[32]),
    .c(cout_13[31]),
    .cout(cout_13[32]),
    .sum(sum_13[32]));
  AL_FADD comp13_33 (
    .a(i13[33]),
    .b(sum_12[33]),
    .c(cout_13[32]),
    .cout(cout_13[33]),
    .sum(sum_13[33]));
  AL_FADD comp13_34 (
    .a(i13[34]),
    .b(sum_12[34]),
    .c(cout_13[33]),
    .cout(cout_13[34]),
    .sum(sum_13[34]));
  AL_FADD comp13_35 (
    .a(i13[35]),
    .b(sum_12[35]),
    .c(cout_13[34]),
    .cout(cout_13[35]),
    .sum(sum_13[35]));
  AL_FADD comp13_36 (
    .a(i13[36]),
    .b(sum_12[36]),
    .c(cout_13[35]),
    .cout(cout_13[36]),
    .sum(sum_13[36]));
  AL_FADD comp13_37 (
    .a(i13[37]),
    .b(sum_12[37]),
    .c(cout_13[36]),
    .cout(cout_13[37]),
    .sum(sum_13[37]));
  AL_FADD comp13_38 (
    .a(i13[38]),
    .b(sum_12[38]),
    .c(cout_13[37]),
    .cout(cout_13[38]),
    .sum(sum_13[38]));
  AL_FADD comp13_39 (
    .a(i13[39]),
    .b(sum_12[39]),
    .c(cout_13[38]),
    .cout(cout_13[39]),
    .sum(sum_13[39]));
  AL_FADD comp13_4 (
    .a(i13[4]),
    .b(sum_12[4]),
    .c(cout_13[3]),
    .cout(cout_13[4]),
    .sum(sum_13[4]));
  AL_FADD comp13_40 (
    .a(i13[40]),
    .b(sum_12[40]),
    .c(cout_13[39]),
    .cout(cout_13[40]),
    .sum(sum_13[40]));
  AL_FADD comp13_41 (
    .a(i13[41]),
    .b(sum_12[41]),
    .c(cout_13[40]),
    .cout(cout_13[41]),
    .sum(sum_13[41]));
  AL_FADD comp13_42 (
    .a(i13[42]),
    .b(sum_12[42]),
    .c(cout_13[41]),
    .cout(cout_13[42]),
    .sum(sum_13[42]));
  AL_FADD comp13_43 (
    .a(i13[43]),
    .b(sum_12[43]),
    .c(cout_13[42]),
    .cout(cout_13[43]),
    .sum(sum_13[43]));
  AL_FADD comp13_44 (
    .a(i13[44]),
    .b(sum_12[44]),
    .c(cout_13[43]),
    .cout(cout_13[44]),
    .sum(sum_13[44]));
  AL_FADD comp13_45 (
    .a(i13[45]),
    .b(sum_12[45]),
    .c(cout_13[44]),
    .cout(cout_13[45]),
    .sum(sum_13[45]));
  AL_FADD comp13_46 (
    .a(i13[46]),
    .b(sum_12[46]),
    .c(cout_13[45]),
    .cout(cout_13[46]),
    .sum(sum_13[46]));
  AL_FADD comp13_47 (
    .a(i13[47]),
    .b(sum_12[47]),
    .c(cout_13[46]),
    .cout(cout_13[47]),
    .sum(sum_13[47]));
  AL_FADD comp13_48 (
    .a(i13[48]),
    .b(sum_12[48]),
    .c(cout_13[47]),
    .cout(cout_13[48]),
    .sum(sum_13[48]));
  AL_FADD comp13_49 (
    .a(i13[49]),
    .b(sum_12[49]),
    .c(cout_13[48]),
    .cout(cout_13[49]),
    .sum(sum_13[49]));
  AL_FADD comp13_5 (
    .a(i13[5]),
    .b(sum_12[5]),
    .c(cout_13[4]),
    .cout(cout_13[5]),
    .sum(sum_13[5]));
  AL_FADD comp13_50 (
    .a(1'b0),
    .b(sum_12[50]),
    .c(cout_13[49]),
    .cout(cout_13[50]),
    .sum(sum_13[50]));
  AL_FADD comp13_51 (
    .a(1'b0),
    .b(sum_12[51]),
    .c(cout_13[50]),
    .cout(cout_13[51]),
    .sum(sum_13[51]));
  AL_FADD comp13_52 (
    .a(1'b0),
    .b(sum_12[52]),
    .c(cout_13[51]),
    .cout(cout_13[52]),
    .sum(sum_13[52]));
  AL_FADD comp13_53 (
    .a(1'b0),
    .b(sum_12[53]),
    .c(cout_13[52]),
    .cout(cout_13[53]),
    .sum(sum_13[53]));
  AL_FADD comp13_54 (
    .a(1'b0),
    .b(sum_12[54]),
    .c(cout_13[53]),
    .cout(cout_13[54]),
    .sum(sum_13[54]));
  AL_FADD comp13_55 (
    .a(1'b0),
    .b(sum_12[55]),
    .c(cout_13[54]),
    .cout(cout_13[55]),
    .sum(sum_13[55]));
  AL_FADD comp13_56 (
    .a(1'b0),
    .b(sum_12[56]),
    .c(cout_13[55]),
    .cout(cout_13[56]),
    .sum(sum_13[56]));
  AL_FADD comp13_57 (
    .a(1'b0),
    .b(sum_12[57]),
    .c(cout_13[56]),
    .cout(cout_13[57]),
    .sum(sum_13[57]));
  AL_FADD comp13_58 (
    .a(1'b0),
    .b(sum_12[58]),
    .c(cout_13[57]),
    .cout(cout_13[58]),
    .sum(sum_13[58]));
  AL_FADD comp13_59 (
    .a(1'b0),
    .b(sum_12[59]),
    .c(cout_13[58]),
    .cout(cout_13[59]),
    .sum(sum_13[59]));
  AL_FADD comp13_6 (
    .a(i13[6]),
    .b(sum_12[6]),
    .c(cout_13[5]),
    .cout(cout_13[6]),
    .sum(sum_13[6]));
  AL_FADD comp13_60 (
    .a(1'b0),
    .b(sum_12[60]),
    .c(cout_13[59]),
    .cout(cout_13[60]),
    .sum(sum_13[60]));
  AL_FADD comp13_61 (
    .a(1'b0),
    .b(sum_12[61]),
    .c(cout_13[60]),
    .cout(cout_13[61]),
    .sum(sum_13[61]));
  AL_FADD comp13_62 (
    .a(1'b0),
    .b(sum_12[62]),
    .c(cout_13[61]),
    .cout(cout_13[62]),
    .sum(sum_13[62]));
  AL_FADD comp13_63 (
    .a(1'b0),
    .b(sum_12[63]),
    .c(cout_13[62]),
    .cout(cout_13[63]),
    .sum(sum_13[63]));
  AL_FADD comp13_7 (
    .a(i13[7]),
    .b(sum_12[7]),
    .c(cout_13[6]),
    .cout(cout_13[7]),
    .sum(sum_13[7]));
  AL_FADD comp13_8 (
    .a(i13[8]),
    .b(sum_12[8]),
    .c(cout_13[7]),
    .cout(cout_13[8]),
    .sum(sum_13[8]));
  AL_FADD comp13_9 (
    .a(i13[9]),
    .b(sum_12[9]),
    .c(cout_13[8]),
    .cout(cout_13[9]),
    .sum(sum_13[9]));
  AL_FADD comp14_0 (
    .a(i14[0]),
    .b(sum_13[0]),
    .c(1'b0),
    .cout(cout_14[0]),
    .sum(sum_14[0]));
  AL_FADD comp14_1 (
    .a(i14[1]),
    .b(sum_13[1]),
    .c(cout_14[0]),
    .cout(cout_14[1]),
    .sum(sum_14[1]));
  AL_FADD comp14_10 (
    .a(i14[10]),
    .b(sum_13[10]),
    .c(cout_14[9]),
    .cout(cout_14[10]),
    .sum(sum_14[10]));
  AL_FADD comp14_11 (
    .a(i14[11]),
    .b(sum_13[11]),
    .c(cout_14[10]),
    .cout(cout_14[11]),
    .sum(sum_14[11]));
  AL_FADD comp14_12 (
    .a(i14[12]),
    .b(sum_13[12]),
    .c(cout_14[11]),
    .cout(cout_14[12]),
    .sum(sum_14[12]));
  AL_FADD comp14_13 (
    .a(i14[13]),
    .b(sum_13[13]),
    .c(cout_14[12]),
    .cout(cout_14[13]),
    .sum(sum_14[13]));
  AL_FADD comp14_14 (
    .a(i14[14]),
    .b(sum_13[14]),
    .c(cout_14[13]),
    .cout(cout_14[14]),
    .sum(sum_14[14]));
  AL_FADD comp14_15 (
    .a(i14[15]),
    .b(sum_13[15]),
    .c(cout_14[14]),
    .cout(cout_14[15]),
    .sum(sum_14[15]));
  AL_FADD comp14_16 (
    .a(i14[16]),
    .b(sum_13[16]),
    .c(cout_14[15]),
    .cout(cout_14[16]),
    .sum(sum_14[16]));
  AL_FADD comp14_17 (
    .a(i14[17]),
    .b(sum_13[17]),
    .c(cout_14[16]),
    .cout(cout_14[17]),
    .sum(sum_14[17]));
  AL_FADD comp14_18 (
    .a(i14[18]),
    .b(sum_13[18]),
    .c(cout_14[17]),
    .cout(cout_14[18]),
    .sum(sum_14[18]));
  AL_FADD comp14_19 (
    .a(i14[19]),
    .b(sum_13[19]),
    .c(cout_14[18]),
    .cout(cout_14[19]),
    .sum(sum_14[19]));
  AL_FADD comp14_2 (
    .a(i14[2]),
    .b(sum_13[2]),
    .c(cout_14[1]),
    .cout(cout_14[2]),
    .sum(sum_14[2]));
  AL_FADD comp14_20 (
    .a(i14[20]),
    .b(sum_13[20]),
    .c(cout_14[19]),
    .cout(cout_14[20]),
    .sum(sum_14[20]));
  AL_FADD comp14_21 (
    .a(i14[21]),
    .b(sum_13[21]),
    .c(cout_14[20]),
    .cout(cout_14[21]),
    .sum(sum_14[21]));
  AL_FADD comp14_22 (
    .a(i14[22]),
    .b(sum_13[22]),
    .c(cout_14[21]),
    .cout(cout_14[22]),
    .sum(sum_14[22]));
  AL_FADD comp14_23 (
    .a(i14[23]),
    .b(sum_13[23]),
    .c(cout_14[22]),
    .cout(cout_14[23]),
    .sum(sum_14[23]));
  AL_FADD comp14_24 (
    .a(i14[24]),
    .b(sum_13[24]),
    .c(cout_14[23]),
    .cout(cout_14[24]),
    .sum(sum_14[24]));
  AL_FADD comp14_25 (
    .a(i14[25]),
    .b(sum_13[25]),
    .c(cout_14[24]),
    .cout(cout_14[25]),
    .sum(sum_14[25]));
  AL_FADD comp14_26 (
    .a(i14[26]),
    .b(sum_13[26]),
    .c(cout_14[25]),
    .cout(cout_14[26]),
    .sum(sum_14[26]));
  AL_FADD comp14_27 (
    .a(i14[27]),
    .b(sum_13[27]),
    .c(cout_14[26]),
    .cout(cout_14[27]),
    .sum(sum_14[27]));
  AL_FADD comp14_28 (
    .a(i14[28]),
    .b(sum_13[28]),
    .c(cout_14[27]),
    .cout(cout_14[28]),
    .sum(sum_14[28]));
  AL_FADD comp14_29 (
    .a(i14[29]),
    .b(sum_13[29]),
    .c(cout_14[28]),
    .cout(cout_14[29]),
    .sum(sum_14[29]));
  AL_FADD comp14_3 (
    .a(i14[3]),
    .b(sum_13[3]),
    .c(cout_14[2]),
    .cout(cout_14[3]),
    .sum(sum_14[3]));
  AL_FADD comp14_30 (
    .a(i14[30]),
    .b(sum_13[30]),
    .c(cout_14[29]),
    .cout(cout_14[30]),
    .sum(sum_14[30]));
  AL_FADD comp14_31 (
    .a(i14[31]),
    .b(sum_13[31]),
    .c(cout_14[30]),
    .cout(cout_14[31]),
    .sum(sum_14[31]));
  AL_FADD comp14_32 (
    .a(i14[32]),
    .b(sum_13[32]),
    .c(cout_14[31]),
    .cout(cout_14[32]),
    .sum(sum_14[32]));
  AL_FADD comp14_33 (
    .a(i14[33]),
    .b(sum_13[33]),
    .c(cout_14[32]),
    .cout(cout_14[33]),
    .sum(sum_14[33]));
  AL_FADD comp14_34 (
    .a(i14[34]),
    .b(sum_13[34]),
    .c(cout_14[33]),
    .cout(cout_14[34]),
    .sum(sum_14[34]));
  AL_FADD comp14_35 (
    .a(i14[35]),
    .b(sum_13[35]),
    .c(cout_14[34]),
    .cout(cout_14[35]),
    .sum(sum_14[35]));
  AL_FADD comp14_36 (
    .a(i14[36]),
    .b(sum_13[36]),
    .c(cout_14[35]),
    .cout(cout_14[36]),
    .sum(sum_14[36]));
  AL_FADD comp14_37 (
    .a(i14[37]),
    .b(sum_13[37]),
    .c(cout_14[36]),
    .cout(cout_14[37]),
    .sum(sum_14[37]));
  AL_FADD comp14_38 (
    .a(i14[38]),
    .b(sum_13[38]),
    .c(cout_14[37]),
    .cout(cout_14[38]),
    .sum(sum_14[38]));
  AL_FADD comp14_39 (
    .a(i14[39]),
    .b(sum_13[39]),
    .c(cout_14[38]),
    .cout(cout_14[39]),
    .sum(sum_14[39]));
  AL_FADD comp14_4 (
    .a(i14[4]),
    .b(sum_13[4]),
    .c(cout_14[3]),
    .cout(cout_14[4]),
    .sum(sum_14[4]));
  AL_FADD comp14_40 (
    .a(i14[40]),
    .b(sum_13[40]),
    .c(cout_14[39]),
    .cout(cout_14[40]),
    .sum(sum_14[40]));
  AL_FADD comp14_41 (
    .a(i14[41]),
    .b(sum_13[41]),
    .c(cout_14[40]),
    .cout(cout_14[41]),
    .sum(sum_14[41]));
  AL_FADD comp14_42 (
    .a(i14[42]),
    .b(sum_13[42]),
    .c(cout_14[41]),
    .cout(cout_14[42]),
    .sum(sum_14[42]));
  AL_FADD comp14_43 (
    .a(i14[43]),
    .b(sum_13[43]),
    .c(cout_14[42]),
    .cout(cout_14[43]),
    .sum(sum_14[43]));
  AL_FADD comp14_44 (
    .a(i14[44]),
    .b(sum_13[44]),
    .c(cout_14[43]),
    .cout(cout_14[44]),
    .sum(sum_14[44]));
  AL_FADD comp14_45 (
    .a(i14[45]),
    .b(sum_13[45]),
    .c(cout_14[44]),
    .cout(cout_14[45]),
    .sum(sum_14[45]));
  AL_FADD comp14_46 (
    .a(i14[46]),
    .b(sum_13[46]),
    .c(cout_14[45]),
    .cout(cout_14[46]),
    .sum(sum_14[46]));
  AL_FADD comp14_47 (
    .a(i14[47]),
    .b(sum_13[47]),
    .c(cout_14[46]),
    .cout(cout_14[47]),
    .sum(sum_14[47]));
  AL_FADD comp14_48 (
    .a(i14[48]),
    .b(sum_13[48]),
    .c(cout_14[47]),
    .cout(cout_14[48]),
    .sum(sum_14[48]));
  AL_FADD comp14_49 (
    .a(1'b0),
    .b(sum_13[49]),
    .c(cout_14[48]),
    .cout(cout_14[49]),
    .sum(sum_14[49]));
  AL_FADD comp14_5 (
    .a(i14[5]),
    .b(sum_13[5]),
    .c(cout_14[4]),
    .cout(cout_14[5]),
    .sum(sum_14[5]));
  AL_FADD comp14_50 (
    .a(1'b0),
    .b(sum_13[50]),
    .c(cout_14[49]),
    .cout(cout_14[50]),
    .sum(sum_14[50]));
  AL_FADD comp14_51 (
    .a(1'b0),
    .b(sum_13[51]),
    .c(cout_14[50]),
    .cout(cout_14[51]),
    .sum(sum_14[51]));
  AL_FADD comp14_52 (
    .a(1'b0),
    .b(sum_13[52]),
    .c(cout_14[51]),
    .cout(cout_14[52]),
    .sum(sum_14[52]));
  AL_FADD comp14_53 (
    .a(1'b0),
    .b(sum_13[53]),
    .c(cout_14[52]),
    .cout(cout_14[53]),
    .sum(sum_14[53]));
  AL_FADD comp14_54 (
    .a(1'b0),
    .b(sum_13[54]),
    .c(cout_14[53]),
    .cout(cout_14[54]),
    .sum(sum_14[54]));
  AL_FADD comp14_55 (
    .a(1'b0),
    .b(sum_13[55]),
    .c(cout_14[54]),
    .cout(cout_14[55]),
    .sum(sum_14[55]));
  AL_FADD comp14_56 (
    .a(1'b0),
    .b(sum_13[56]),
    .c(cout_14[55]),
    .cout(cout_14[56]),
    .sum(sum_14[56]));
  AL_FADD comp14_57 (
    .a(1'b0),
    .b(sum_13[57]),
    .c(cout_14[56]),
    .cout(cout_14[57]),
    .sum(sum_14[57]));
  AL_FADD comp14_58 (
    .a(1'b0),
    .b(sum_13[58]),
    .c(cout_14[57]),
    .cout(cout_14[58]),
    .sum(sum_14[58]));
  AL_FADD comp14_59 (
    .a(1'b0),
    .b(sum_13[59]),
    .c(cout_14[58]),
    .cout(cout_14[59]),
    .sum(sum_14[59]));
  AL_FADD comp14_6 (
    .a(i14[6]),
    .b(sum_13[6]),
    .c(cout_14[5]),
    .cout(cout_14[6]),
    .sum(sum_14[6]));
  AL_FADD comp14_60 (
    .a(1'b0),
    .b(sum_13[60]),
    .c(cout_14[59]),
    .cout(cout_14[60]),
    .sum(sum_14[60]));
  AL_FADD comp14_61 (
    .a(1'b0),
    .b(sum_13[61]),
    .c(cout_14[60]),
    .cout(cout_14[61]),
    .sum(sum_14[61]));
  AL_FADD comp14_62 (
    .a(1'b0),
    .b(sum_13[62]),
    .c(cout_14[61]),
    .cout(cout_14[62]),
    .sum(sum_14[62]));
  AL_FADD comp14_63 (
    .a(1'b0),
    .b(sum_13[63]),
    .c(cout_14[62]),
    .cout(cout_14[63]),
    .sum(sum_14[63]));
  AL_FADD comp14_7 (
    .a(i14[7]),
    .b(sum_13[7]),
    .c(cout_14[6]),
    .cout(cout_14[7]),
    .sum(sum_14[7]));
  AL_FADD comp14_8 (
    .a(i14[8]),
    .b(sum_13[8]),
    .c(cout_14[7]),
    .cout(cout_14[8]),
    .sum(sum_14[8]));
  AL_FADD comp14_9 (
    .a(i14[9]),
    .b(sum_13[9]),
    .c(cout_14[8]),
    .cout(cout_14[9]),
    .sum(sum_14[9]));
  AL_FADD comp15_0 (
    .a(i15[0]),
    .b(sum_14[0]),
    .c(1'b0),
    .cout(cout_15[0]),
    .sum(sum_15[0]));
  AL_FADD comp15_1 (
    .a(i15[1]),
    .b(sum_14[1]),
    .c(cout_15[0]),
    .cout(cout_15[1]),
    .sum(sum_15[1]));
  AL_FADD comp15_10 (
    .a(i15[10]),
    .b(sum_14[10]),
    .c(cout_15[9]),
    .cout(cout_15[10]),
    .sum(sum_15[10]));
  AL_FADD comp15_11 (
    .a(i15[11]),
    .b(sum_14[11]),
    .c(cout_15[10]),
    .cout(cout_15[11]),
    .sum(sum_15[11]));
  AL_FADD comp15_12 (
    .a(i15[12]),
    .b(sum_14[12]),
    .c(cout_15[11]),
    .cout(cout_15[12]),
    .sum(sum_15[12]));
  AL_FADD comp15_13 (
    .a(i15[13]),
    .b(sum_14[13]),
    .c(cout_15[12]),
    .cout(cout_15[13]),
    .sum(sum_15[13]));
  AL_FADD comp15_14 (
    .a(i15[14]),
    .b(sum_14[14]),
    .c(cout_15[13]),
    .cout(cout_15[14]),
    .sum(sum_15[14]));
  AL_FADD comp15_15 (
    .a(i15[15]),
    .b(sum_14[15]),
    .c(cout_15[14]),
    .cout(cout_15[15]),
    .sum(sum_15[15]));
  AL_FADD comp15_16 (
    .a(i15[16]),
    .b(sum_14[16]),
    .c(cout_15[15]),
    .cout(cout_15[16]),
    .sum(sum_15[16]));
  AL_FADD comp15_17 (
    .a(i15[17]),
    .b(sum_14[17]),
    .c(cout_15[16]),
    .cout(cout_15[17]),
    .sum(sum_15[17]));
  AL_FADD comp15_18 (
    .a(i15[18]),
    .b(sum_14[18]),
    .c(cout_15[17]),
    .cout(cout_15[18]),
    .sum(sum_15[18]));
  AL_FADD comp15_19 (
    .a(i15[19]),
    .b(sum_14[19]),
    .c(cout_15[18]),
    .cout(cout_15[19]),
    .sum(sum_15[19]));
  AL_FADD comp15_2 (
    .a(i15[2]),
    .b(sum_14[2]),
    .c(cout_15[1]),
    .cout(cout_15[2]),
    .sum(sum_15[2]));
  AL_FADD comp15_20 (
    .a(i15[20]),
    .b(sum_14[20]),
    .c(cout_15[19]),
    .cout(cout_15[20]),
    .sum(sum_15[20]));
  AL_FADD comp15_21 (
    .a(i15[21]),
    .b(sum_14[21]),
    .c(cout_15[20]),
    .cout(cout_15[21]),
    .sum(sum_15[21]));
  AL_FADD comp15_22 (
    .a(i15[22]),
    .b(sum_14[22]),
    .c(cout_15[21]),
    .cout(cout_15[22]),
    .sum(sum_15[22]));
  AL_FADD comp15_23 (
    .a(i15[23]),
    .b(sum_14[23]),
    .c(cout_15[22]),
    .cout(cout_15[23]),
    .sum(sum_15[23]));
  AL_FADD comp15_24 (
    .a(i15[24]),
    .b(sum_14[24]),
    .c(cout_15[23]),
    .cout(cout_15[24]),
    .sum(sum_15[24]));
  AL_FADD comp15_25 (
    .a(i15[25]),
    .b(sum_14[25]),
    .c(cout_15[24]),
    .cout(cout_15[25]),
    .sum(sum_15[25]));
  AL_FADD comp15_26 (
    .a(i15[26]),
    .b(sum_14[26]),
    .c(cout_15[25]),
    .cout(cout_15[26]),
    .sum(sum_15[26]));
  AL_FADD comp15_27 (
    .a(i15[27]),
    .b(sum_14[27]),
    .c(cout_15[26]),
    .cout(cout_15[27]),
    .sum(sum_15[27]));
  AL_FADD comp15_28 (
    .a(i15[28]),
    .b(sum_14[28]),
    .c(cout_15[27]),
    .cout(cout_15[28]),
    .sum(sum_15[28]));
  AL_FADD comp15_29 (
    .a(i15[29]),
    .b(sum_14[29]),
    .c(cout_15[28]),
    .cout(cout_15[29]),
    .sum(sum_15[29]));
  AL_FADD comp15_3 (
    .a(i15[3]),
    .b(sum_14[3]),
    .c(cout_15[2]),
    .cout(cout_15[3]),
    .sum(sum_15[3]));
  AL_FADD comp15_30 (
    .a(i15[30]),
    .b(sum_14[30]),
    .c(cout_15[29]),
    .cout(cout_15[30]),
    .sum(sum_15[30]));
  AL_FADD comp15_31 (
    .a(i15[31]),
    .b(sum_14[31]),
    .c(cout_15[30]),
    .cout(cout_15[31]),
    .sum(sum_15[31]));
  AL_FADD comp15_32 (
    .a(i15[32]),
    .b(sum_14[32]),
    .c(cout_15[31]),
    .cout(cout_15[32]),
    .sum(sum_15[32]));
  AL_FADD comp15_33 (
    .a(i15[33]),
    .b(sum_14[33]),
    .c(cout_15[32]),
    .cout(cout_15[33]),
    .sum(sum_15[33]));
  AL_FADD comp15_34 (
    .a(i15[34]),
    .b(sum_14[34]),
    .c(cout_15[33]),
    .cout(cout_15[34]),
    .sum(sum_15[34]));
  AL_FADD comp15_35 (
    .a(i15[35]),
    .b(sum_14[35]),
    .c(cout_15[34]),
    .cout(cout_15[35]),
    .sum(sum_15[35]));
  AL_FADD comp15_36 (
    .a(i15[36]),
    .b(sum_14[36]),
    .c(cout_15[35]),
    .cout(cout_15[36]),
    .sum(sum_15[36]));
  AL_FADD comp15_37 (
    .a(i15[37]),
    .b(sum_14[37]),
    .c(cout_15[36]),
    .cout(cout_15[37]),
    .sum(sum_15[37]));
  AL_FADD comp15_38 (
    .a(i15[38]),
    .b(sum_14[38]),
    .c(cout_15[37]),
    .cout(cout_15[38]),
    .sum(sum_15[38]));
  AL_FADD comp15_39 (
    .a(i15[39]),
    .b(sum_14[39]),
    .c(cout_15[38]),
    .cout(cout_15[39]),
    .sum(sum_15[39]));
  AL_FADD comp15_4 (
    .a(i15[4]),
    .b(sum_14[4]),
    .c(cout_15[3]),
    .cout(cout_15[4]),
    .sum(sum_15[4]));
  AL_FADD comp15_40 (
    .a(i15[40]),
    .b(sum_14[40]),
    .c(cout_15[39]),
    .cout(cout_15[40]),
    .sum(sum_15[40]));
  AL_FADD comp15_41 (
    .a(i15[41]),
    .b(sum_14[41]),
    .c(cout_15[40]),
    .cout(cout_15[41]),
    .sum(sum_15[41]));
  AL_FADD comp15_42 (
    .a(i15[42]),
    .b(sum_14[42]),
    .c(cout_15[41]),
    .cout(cout_15[42]),
    .sum(sum_15[42]));
  AL_FADD comp15_43 (
    .a(i15[43]),
    .b(sum_14[43]),
    .c(cout_15[42]),
    .cout(cout_15[43]),
    .sum(sum_15[43]));
  AL_FADD comp15_44 (
    .a(i15[44]),
    .b(sum_14[44]),
    .c(cout_15[43]),
    .cout(cout_15[44]),
    .sum(sum_15[44]));
  AL_FADD comp15_45 (
    .a(i15[45]),
    .b(sum_14[45]),
    .c(cout_15[44]),
    .cout(cout_15[45]),
    .sum(sum_15[45]));
  AL_FADD comp15_46 (
    .a(i15[46]),
    .b(sum_14[46]),
    .c(cout_15[45]),
    .cout(cout_15[46]),
    .sum(sum_15[46]));
  AL_FADD comp15_47 (
    .a(i15[47]),
    .b(sum_14[47]),
    .c(cout_15[46]),
    .cout(cout_15[47]),
    .sum(sum_15[47]));
  AL_FADD comp15_48 (
    .a(1'b0),
    .b(sum_14[48]),
    .c(cout_15[47]),
    .cout(cout_15[48]),
    .sum(sum_15[48]));
  AL_FADD comp15_49 (
    .a(1'b0),
    .b(sum_14[49]),
    .c(cout_15[48]),
    .cout(cout_15[49]),
    .sum(sum_15[49]));
  AL_FADD comp15_5 (
    .a(i15[5]),
    .b(sum_14[5]),
    .c(cout_15[4]),
    .cout(cout_15[5]),
    .sum(sum_15[5]));
  AL_FADD comp15_50 (
    .a(1'b0),
    .b(sum_14[50]),
    .c(cout_15[49]),
    .cout(cout_15[50]),
    .sum(sum_15[50]));
  AL_FADD comp15_51 (
    .a(1'b0),
    .b(sum_14[51]),
    .c(cout_15[50]),
    .cout(cout_15[51]),
    .sum(sum_15[51]));
  AL_FADD comp15_52 (
    .a(1'b0),
    .b(sum_14[52]),
    .c(cout_15[51]),
    .cout(cout_15[52]),
    .sum(sum_15[52]));
  AL_FADD comp15_53 (
    .a(1'b0),
    .b(sum_14[53]),
    .c(cout_15[52]),
    .cout(cout_15[53]),
    .sum(sum_15[53]));
  AL_FADD comp15_54 (
    .a(1'b0),
    .b(sum_14[54]),
    .c(cout_15[53]),
    .cout(cout_15[54]),
    .sum(sum_15[54]));
  AL_FADD comp15_55 (
    .a(1'b0),
    .b(sum_14[55]),
    .c(cout_15[54]),
    .cout(cout_15[55]),
    .sum(sum_15[55]));
  AL_FADD comp15_56 (
    .a(1'b0),
    .b(sum_14[56]),
    .c(cout_15[55]),
    .cout(cout_15[56]),
    .sum(sum_15[56]));
  AL_FADD comp15_57 (
    .a(1'b0),
    .b(sum_14[57]),
    .c(cout_15[56]),
    .cout(cout_15[57]),
    .sum(sum_15[57]));
  AL_FADD comp15_58 (
    .a(1'b0),
    .b(sum_14[58]),
    .c(cout_15[57]),
    .cout(cout_15[58]),
    .sum(sum_15[58]));
  AL_FADD comp15_59 (
    .a(1'b0),
    .b(sum_14[59]),
    .c(cout_15[58]),
    .cout(cout_15[59]),
    .sum(sum_15[59]));
  AL_FADD comp15_6 (
    .a(i15[6]),
    .b(sum_14[6]),
    .c(cout_15[5]),
    .cout(cout_15[6]),
    .sum(sum_15[6]));
  AL_FADD comp15_60 (
    .a(1'b0),
    .b(sum_14[60]),
    .c(cout_15[59]),
    .cout(cout_15[60]),
    .sum(sum_15[60]));
  AL_FADD comp15_61 (
    .a(1'b0),
    .b(sum_14[61]),
    .c(cout_15[60]),
    .cout(cout_15[61]),
    .sum(sum_15[61]));
  AL_FADD comp15_62 (
    .a(1'b0),
    .b(sum_14[62]),
    .c(cout_15[61]),
    .cout(cout_15[62]),
    .sum(sum_15[62]));
  AL_FADD comp15_63 (
    .a(1'b0),
    .b(sum_14[63]),
    .c(cout_15[62]),
    .cout(cout_15[63]),
    .sum(sum_15[63]));
  AL_FADD comp15_7 (
    .a(i15[7]),
    .b(sum_14[7]),
    .c(cout_15[6]),
    .cout(cout_15[7]),
    .sum(sum_15[7]));
  AL_FADD comp15_8 (
    .a(i15[8]),
    .b(sum_14[8]),
    .c(cout_15[7]),
    .cout(cout_15[8]),
    .sum(sum_15[8]));
  AL_FADD comp15_9 (
    .a(i15[9]),
    .b(sum_14[9]),
    .c(cout_15[8]),
    .cout(cout_15[9]),
    .sum(sum_15[9]));
  AL_FADD comp16_0 (
    .a(i16[0]),
    .b(sum_15[0]),
    .c(1'b0),
    .cout(cout_16[0]),
    .sum(sum_16[0]));
  AL_FADD comp16_1 (
    .a(i16[1]),
    .b(sum_15[1]),
    .c(cout_16[0]),
    .cout(cout_16[1]),
    .sum(sum_16[1]));
  AL_FADD comp16_10 (
    .a(i16[10]),
    .b(sum_15[10]),
    .c(cout_16[9]),
    .cout(cout_16[10]),
    .sum(sum_16[10]));
  AL_FADD comp16_11 (
    .a(i16[11]),
    .b(sum_15[11]),
    .c(cout_16[10]),
    .cout(cout_16[11]),
    .sum(sum_16[11]));
  AL_FADD comp16_12 (
    .a(i16[12]),
    .b(sum_15[12]),
    .c(cout_16[11]),
    .cout(cout_16[12]),
    .sum(sum_16[12]));
  AL_FADD comp16_13 (
    .a(i16[13]),
    .b(sum_15[13]),
    .c(cout_16[12]),
    .cout(cout_16[13]),
    .sum(sum_16[13]));
  AL_FADD comp16_14 (
    .a(i16[14]),
    .b(sum_15[14]),
    .c(cout_16[13]),
    .cout(cout_16[14]),
    .sum(sum_16[14]));
  AL_FADD comp16_15 (
    .a(i16[15]),
    .b(sum_15[15]),
    .c(cout_16[14]),
    .cout(cout_16[15]),
    .sum(sum_16[15]));
  AL_FADD comp16_16 (
    .a(i16[16]),
    .b(sum_15[16]),
    .c(cout_16[15]),
    .cout(cout_16[16]),
    .sum(sum_16[16]));
  AL_FADD comp16_17 (
    .a(i16[17]),
    .b(sum_15[17]),
    .c(cout_16[16]),
    .cout(cout_16[17]),
    .sum(sum_16[17]));
  AL_FADD comp16_18 (
    .a(i16[18]),
    .b(sum_15[18]),
    .c(cout_16[17]),
    .cout(cout_16[18]),
    .sum(sum_16[18]));
  AL_FADD comp16_19 (
    .a(i16[19]),
    .b(sum_15[19]),
    .c(cout_16[18]),
    .cout(cout_16[19]),
    .sum(sum_16[19]));
  AL_FADD comp16_2 (
    .a(i16[2]),
    .b(sum_15[2]),
    .c(cout_16[1]),
    .cout(cout_16[2]),
    .sum(sum_16[2]));
  AL_FADD comp16_20 (
    .a(i16[20]),
    .b(sum_15[20]),
    .c(cout_16[19]),
    .cout(cout_16[20]),
    .sum(sum_16[20]));
  AL_FADD comp16_21 (
    .a(i16[21]),
    .b(sum_15[21]),
    .c(cout_16[20]),
    .cout(cout_16[21]),
    .sum(sum_16[21]));
  AL_FADD comp16_22 (
    .a(i16[22]),
    .b(sum_15[22]),
    .c(cout_16[21]),
    .cout(cout_16[22]),
    .sum(sum_16[22]));
  AL_FADD comp16_23 (
    .a(i16[23]),
    .b(sum_15[23]),
    .c(cout_16[22]),
    .cout(cout_16[23]),
    .sum(sum_16[23]));
  AL_FADD comp16_24 (
    .a(i16[24]),
    .b(sum_15[24]),
    .c(cout_16[23]),
    .cout(cout_16[24]),
    .sum(sum_16[24]));
  AL_FADD comp16_25 (
    .a(i16[25]),
    .b(sum_15[25]),
    .c(cout_16[24]),
    .cout(cout_16[25]),
    .sum(sum_16[25]));
  AL_FADD comp16_26 (
    .a(i16[26]),
    .b(sum_15[26]),
    .c(cout_16[25]),
    .cout(cout_16[26]),
    .sum(sum_16[26]));
  AL_FADD comp16_27 (
    .a(i16[27]),
    .b(sum_15[27]),
    .c(cout_16[26]),
    .cout(cout_16[27]),
    .sum(sum_16[27]));
  AL_FADD comp16_28 (
    .a(i16[28]),
    .b(sum_15[28]),
    .c(cout_16[27]),
    .cout(cout_16[28]),
    .sum(sum_16[28]));
  AL_FADD comp16_29 (
    .a(i16[29]),
    .b(sum_15[29]),
    .c(cout_16[28]),
    .cout(cout_16[29]),
    .sum(sum_16[29]));
  AL_FADD comp16_3 (
    .a(i16[3]),
    .b(sum_15[3]),
    .c(cout_16[2]),
    .cout(cout_16[3]),
    .sum(sum_16[3]));
  AL_FADD comp16_30 (
    .a(i16[30]),
    .b(sum_15[30]),
    .c(cout_16[29]),
    .cout(cout_16[30]),
    .sum(sum_16[30]));
  AL_FADD comp16_31 (
    .a(i16[31]),
    .b(sum_15[31]),
    .c(cout_16[30]),
    .cout(cout_16[31]),
    .sum(sum_16[31]));
  AL_FADD comp16_32 (
    .a(i16[32]),
    .b(sum_15[32]),
    .c(cout_16[31]),
    .cout(cout_16[32]),
    .sum(sum_16[32]));
  AL_FADD comp16_33 (
    .a(i16[33]),
    .b(sum_15[33]),
    .c(cout_16[32]),
    .cout(cout_16[33]),
    .sum(sum_16[33]));
  AL_FADD comp16_34 (
    .a(i16[34]),
    .b(sum_15[34]),
    .c(cout_16[33]),
    .cout(cout_16[34]),
    .sum(sum_16[34]));
  AL_FADD comp16_35 (
    .a(i16[35]),
    .b(sum_15[35]),
    .c(cout_16[34]),
    .cout(cout_16[35]),
    .sum(sum_16[35]));
  AL_FADD comp16_36 (
    .a(i16[36]),
    .b(sum_15[36]),
    .c(cout_16[35]),
    .cout(cout_16[36]),
    .sum(sum_16[36]));
  AL_FADD comp16_37 (
    .a(i16[37]),
    .b(sum_15[37]),
    .c(cout_16[36]),
    .cout(cout_16[37]),
    .sum(sum_16[37]));
  AL_FADD comp16_38 (
    .a(i16[38]),
    .b(sum_15[38]),
    .c(cout_16[37]),
    .cout(cout_16[38]),
    .sum(sum_16[38]));
  AL_FADD comp16_39 (
    .a(i16[39]),
    .b(sum_15[39]),
    .c(cout_16[38]),
    .cout(cout_16[39]),
    .sum(sum_16[39]));
  AL_FADD comp16_4 (
    .a(i16[4]),
    .b(sum_15[4]),
    .c(cout_16[3]),
    .cout(cout_16[4]),
    .sum(sum_16[4]));
  AL_FADD comp16_40 (
    .a(i16[40]),
    .b(sum_15[40]),
    .c(cout_16[39]),
    .cout(cout_16[40]),
    .sum(sum_16[40]));
  AL_FADD comp16_41 (
    .a(i16[41]),
    .b(sum_15[41]),
    .c(cout_16[40]),
    .cout(cout_16[41]),
    .sum(sum_16[41]));
  AL_FADD comp16_42 (
    .a(i16[42]),
    .b(sum_15[42]),
    .c(cout_16[41]),
    .cout(cout_16[42]),
    .sum(sum_16[42]));
  AL_FADD comp16_43 (
    .a(i16[43]),
    .b(sum_15[43]),
    .c(cout_16[42]),
    .cout(cout_16[43]),
    .sum(sum_16[43]));
  AL_FADD comp16_44 (
    .a(i16[44]),
    .b(sum_15[44]),
    .c(cout_16[43]),
    .cout(cout_16[44]),
    .sum(sum_16[44]));
  AL_FADD comp16_45 (
    .a(i16[45]),
    .b(sum_15[45]),
    .c(cout_16[44]),
    .cout(cout_16[45]),
    .sum(sum_16[45]));
  AL_FADD comp16_46 (
    .a(i16[46]),
    .b(sum_15[46]),
    .c(cout_16[45]),
    .cout(cout_16[46]),
    .sum(sum_16[46]));
  AL_FADD comp16_47 (
    .a(1'b0),
    .b(sum_15[47]),
    .c(cout_16[46]),
    .cout(cout_16[47]),
    .sum(sum_16[47]));
  AL_FADD comp16_48 (
    .a(1'b0),
    .b(sum_15[48]),
    .c(cout_16[47]),
    .cout(cout_16[48]),
    .sum(sum_16[48]));
  AL_FADD comp16_49 (
    .a(1'b0),
    .b(sum_15[49]),
    .c(cout_16[48]),
    .cout(cout_16[49]),
    .sum(sum_16[49]));
  AL_FADD comp16_5 (
    .a(i16[5]),
    .b(sum_15[5]),
    .c(cout_16[4]),
    .cout(cout_16[5]),
    .sum(sum_16[5]));
  AL_FADD comp16_50 (
    .a(1'b0),
    .b(sum_15[50]),
    .c(cout_16[49]),
    .cout(cout_16[50]),
    .sum(sum_16[50]));
  AL_FADD comp16_51 (
    .a(1'b0),
    .b(sum_15[51]),
    .c(cout_16[50]),
    .cout(cout_16[51]),
    .sum(sum_16[51]));
  AL_FADD comp16_52 (
    .a(1'b0),
    .b(sum_15[52]),
    .c(cout_16[51]),
    .cout(cout_16[52]),
    .sum(sum_16[52]));
  AL_FADD comp16_53 (
    .a(1'b0),
    .b(sum_15[53]),
    .c(cout_16[52]),
    .cout(cout_16[53]),
    .sum(sum_16[53]));
  AL_FADD comp16_54 (
    .a(1'b0),
    .b(sum_15[54]),
    .c(cout_16[53]),
    .cout(cout_16[54]),
    .sum(sum_16[54]));
  AL_FADD comp16_55 (
    .a(1'b0),
    .b(sum_15[55]),
    .c(cout_16[54]),
    .cout(cout_16[55]),
    .sum(sum_16[55]));
  AL_FADD comp16_56 (
    .a(1'b0),
    .b(sum_15[56]),
    .c(cout_16[55]),
    .cout(cout_16[56]),
    .sum(sum_16[56]));
  AL_FADD comp16_57 (
    .a(1'b0),
    .b(sum_15[57]),
    .c(cout_16[56]),
    .cout(cout_16[57]),
    .sum(sum_16[57]));
  AL_FADD comp16_58 (
    .a(1'b0),
    .b(sum_15[58]),
    .c(cout_16[57]),
    .cout(cout_16[58]),
    .sum(sum_16[58]));
  AL_FADD comp16_59 (
    .a(1'b0),
    .b(sum_15[59]),
    .c(cout_16[58]),
    .cout(cout_16[59]),
    .sum(sum_16[59]));
  AL_FADD comp16_6 (
    .a(i16[6]),
    .b(sum_15[6]),
    .c(cout_16[5]),
    .cout(cout_16[6]),
    .sum(sum_16[6]));
  AL_FADD comp16_60 (
    .a(1'b0),
    .b(sum_15[60]),
    .c(cout_16[59]),
    .cout(cout_16[60]),
    .sum(sum_16[60]));
  AL_FADD comp16_61 (
    .a(1'b0),
    .b(sum_15[61]),
    .c(cout_16[60]),
    .cout(cout_16[61]),
    .sum(sum_16[61]));
  AL_FADD comp16_62 (
    .a(1'b0),
    .b(sum_15[62]),
    .c(cout_16[61]),
    .cout(cout_16[62]),
    .sum(sum_16[62]));
  AL_FADD comp16_63 (
    .a(1'b0),
    .b(sum_15[63]),
    .c(cout_16[62]),
    .cout(cout_16[63]),
    .sum(sum_16[63]));
  AL_FADD comp16_7 (
    .a(i16[7]),
    .b(sum_15[7]),
    .c(cout_16[6]),
    .cout(cout_16[7]),
    .sum(sum_16[7]));
  AL_FADD comp16_8 (
    .a(i16[8]),
    .b(sum_15[8]),
    .c(cout_16[7]),
    .cout(cout_16[8]),
    .sum(sum_16[8]));
  AL_FADD comp16_9 (
    .a(i16[9]),
    .b(sum_15[9]),
    .c(cout_16[8]),
    .cout(cout_16[9]),
    .sum(sum_16[9]));
  AL_FADD comp17_0 (
    .a(i17[0]),
    .b(sum_16[0]),
    .c(1'b0),
    .cout(cout_17[0]),
    .sum(sum_17[0]));
  AL_FADD comp17_1 (
    .a(i17[1]),
    .b(sum_16[1]),
    .c(cout_17[0]),
    .cout(cout_17[1]),
    .sum(sum_17[1]));
  AL_FADD comp17_10 (
    .a(i17[10]),
    .b(sum_16[10]),
    .c(cout_17[9]),
    .cout(cout_17[10]),
    .sum(sum_17[10]));
  AL_FADD comp17_11 (
    .a(i17[11]),
    .b(sum_16[11]),
    .c(cout_17[10]),
    .cout(cout_17[11]),
    .sum(sum_17[11]));
  AL_FADD comp17_12 (
    .a(i17[12]),
    .b(sum_16[12]),
    .c(cout_17[11]),
    .cout(cout_17[12]),
    .sum(sum_17[12]));
  AL_FADD comp17_13 (
    .a(i17[13]),
    .b(sum_16[13]),
    .c(cout_17[12]),
    .cout(cout_17[13]),
    .sum(sum_17[13]));
  AL_FADD comp17_14 (
    .a(i17[14]),
    .b(sum_16[14]),
    .c(cout_17[13]),
    .cout(cout_17[14]),
    .sum(sum_17[14]));
  AL_FADD comp17_15 (
    .a(i17[15]),
    .b(sum_16[15]),
    .c(cout_17[14]),
    .cout(cout_17[15]),
    .sum(sum_17[15]));
  AL_FADD comp17_16 (
    .a(i17[16]),
    .b(sum_16[16]),
    .c(cout_17[15]),
    .cout(cout_17[16]),
    .sum(sum_17[16]));
  AL_FADD comp17_17 (
    .a(i17[17]),
    .b(sum_16[17]),
    .c(cout_17[16]),
    .cout(cout_17[17]),
    .sum(sum_17[17]));
  AL_FADD comp17_18 (
    .a(i17[18]),
    .b(sum_16[18]),
    .c(cout_17[17]),
    .cout(cout_17[18]),
    .sum(sum_17[18]));
  AL_FADD comp17_19 (
    .a(i17[19]),
    .b(sum_16[19]),
    .c(cout_17[18]),
    .cout(cout_17[19]),
    .sum(sum_17[19]));
  AL_FADD comp17_2 (
    .a(i17[2]),
    .b(sum_16[2]),
    .c(cout_17[1]),
    .cout(cout_17[2]),
    .sum(sum_17[2]));
  AL_FADD comp17_20 (
    .a(i17[20]),
    .b(sum_16[20]),
    .c(cout_17[19]),
    .cout(cout_17[20]),
    .sum(sum_17[20]));
  AL_FADD comp17_21 (
    .a(i17[21]),
    .b(sum_16[21]),
    .c(cout_17[20]),
    .cout(cout_17[21]),
    .sum(sum_17[21]));
  AL_FADD comp17_22 (
    .a(i17[22]),
    .b(sum_16[22]),
    .c(cout_17[21]),
    .cout(cout_17[22]),
    .sum(sum_17[22]));
  AL_FADD comp17_23 (
    .a(i17[23]),
    .b(sum_16[23]),
    .c(cout_17[22]),
    .cout(cout_17[23]),
    .sum(sum_17[23]));
  AL_FADD comp17_24 (
    .a(i17[24]),
    .b(sum_16[24]),
    .c(cout_17[23]),
    .cout(cout_17[24]),
    .sum(sum_17[24]));
  AL_FADD comp17_25 (
    .a(i17[25]),
    .b(sum_16[25]),
    .c(cout_17[24]),
    .cout(cout_17[25]),
    .sum(sum_17[25]));
  AL_FADD comp17_26 (
    .a(i17[26]),
    .b(sum_16[26]),
    .c(cout_17[25]),
    .cout(cout_17[26]),
    .sum(sum_17[26]));
  AL_FADD comp17_27 (
    .a(i17[27]),
    .b(sum_16[27]),
    .c(cout_17[26]),
    .cout(cout_17[27]),
    .sum(sum_17[27]));
  AL_FADD comp17_28 (
    .a(i17[28]),
    .b(sum_16[28]),
    .c(cout_17[27]),
    .cout(cout_17[28]),
    .sum(sum_17[28]));
  AL_FADD comp17_29 (
    .a(i17[29]),
    .b(sum_16[29]),
    .c(cout_17[28]),
    .cout(cout_17[29]),
    .sum(sum_17[29]));
  AL_FADD comp17_3 (
    .a(i17[3]),
    .b(sum_16[3]),
    .c(cout_17[2]),
    .cout(cout_17[3]),
    .sum(sum_17[3]));
  AL_FADD comp17_30 (
    .a(i17[30]),
    .b(sum_16[30]),
    .c(cout_17[29]),
    .cout(cout_17[30]),
    .sum(sum_17[30]));
  AL_FADD comp17_31 (
    .a(i17[31]),
    .b(sum_16[31]),
    .c(cout_17[30]),
    .cout(cout_17[31]),
    .sum(sum_17[31]));
  AL_FADD comp17_32 (
    .a(i17[32]),
    .b(sum_16[32]),
    .c(cout_17[31]),
    .cout(cout_17[32]),
    .sum(sum_17[32]));
  AL_FADD comp17_33 (
    .a(i17[33]),
    .b(sum_16[33]),
    .c(cout_17[32]),
    .cout(cout_17[33]),
    .sum(sum_17[33]));
  AL_FADD comp17_34 (
    .a(i17[34]),
    .b(sum_16[34]),
    .c(cout_17[33]),
    .cout(cout_17[34]),
    .sum(sum_17[34]));
  AL_FADD comp17_35 (
    .a(i17[35]),
    .b(sum_16[35]),
    .c(cout_17[34]),
    .cout(cout_17[35]),
    .sum(sum_17[35]));
  AL_FADD comp17_36 (
    .a(i17[36]),
    .b(sum_16[36]),
    .c(cout_17[35]),
    .cout(cout_17[36]),
    .sum(sum_17[36]));
  AL_FADD comp17_37 (
    .a(i17[37]),
    .b(sum_16[37]),
    .c(cout_17[36]),
    .cout(cout_17[37]),
    .sum(sum_17[37]));
  AL_FADD comp17_38 (
    .a(i17[38]),
    .b(sum_16[38]),
    .c(cout_17[37]),
    .cout(cout_17[38]),
    .sum(sum_17[38]));
  AL_FADD comp17_39 (
    .a(i17[39]),
    .b(sum_16[39]),
    .c(cout_17[38]),
    .cout(cout_17[39]),
    .sum(sum_17[39]));
  AL_FADD comp17_4 (
    .a(i17[4]),
    .b(sum_16[4]),
    .c(cout_17[3]),
    .cout(cout_17[4]),
    .sum(sum_17[4]));
  AL_FADD comp17_40 (
    .a(i17[40]),
    .b(sum_16[40]),
    .c(cout_17[39]),
    .cout(cout_17[40]),
    .sum(sum_17[40]));
  AL_FADD comp17_41 (
    .a(i17[41]),
    .b(sum_16[41]),
    .c(cout_17[40]),
    .cout(cout_17[41]),
    .sum(sum_17[41]));
  AL_FADD comp17_42 (
    .a(i17[42]),
    .b(sum_16[42]),
    .c(cout_17[41]),
    .cout(cout_17[42]),
    .sum(sum_17[42]));
  AL_FADD comp17_43 (
    .a(i17[43]),
    .b(sum_16[43]),
    .c(cout_17[42]),
    .cout(cout_17[43]),
    .sum(sum_17[43]));
  AL_FADD comp17_44 (
    .a(i17[44]),
    .b(sum_16[44]),
    .c(cout_17[43]),
    .cout(cout_17[44]),
    .sum(sum_17[44]));
  AL_FADD comp17_45 (
    .a(i17[45]),
    .b(sum_16[45]),
    .c(cout_17[44]),
    .cout(cout_17[45]),
    .sum(sum_17[45]));
  AL_FADD comp17_46 (
    .a(1'b0),
    .b(sum_16[46]),
    .c(cout_17[45]),
    .cout(cout_17[46]),
    .sum(sum_17[46]));
  AL_FADD comp17_47 (
    .a(1'b0),
    .b(sum_16[47]),
    .c(cout_17[46]),
    .cout(cout_17[47]),
    .sum(sum_17[47]));
  AL_FADD comp17_48 (
    .a(1'b0),
    .b(sum_16[48]),
    .c(cout_17[47]),
    .cout(cout_17[48]),
    .sum(sum_17[48]));
  AL_FADD comp17_49 (
    .a(1'b0),
    .b(sum_16[49]),
    .c(cout_17[48]),
    .cout(cout_17[49]),
    .sum(sum_17[49]));
  AL_FADD comp17_5 (
    .a(i17[5]),
    .b(sum_16[5]),
    .c(cout_17[4]),
    .cout(cout_17[5]),
    .sum(sum_17[5]));
  AL_FADD comp17_50 (
    .a(1'b0),
    .b(sum_16[50]),
    .c(cout_17[49]),
    .cout(cout_17[50]),
    .sum(sum_17[50]));
  AL_FADD comp17_51 (
    .a(1'b0),
    .b(sum_16[51]),
    .c(cout_17[50]),
    .cout(cout_17[51]),
    .sum(sum_17[51]));
  AL_FADD comp17_52 (
    .a(1'b0),
    .b(sum_16[52]),
    .c(cout_17[51]),
    .cout(cout_17[52]),
    .sum(sum_17[52]));
  AL_FADD comp17_53 (
    .a(1'b0),
    .b(sum_16[53]),
    .c(cout_17[52]),
    .cout(cout_17[53]),
    .sum(sum_17[53]));
  AL_FADD comp17_54 (
    .a(1'b0),
    .b(sum_16[54]),
    .c(cout_17[53]),
    .cout(cout_17[54]),
    .sum(sum_17[54]));
  AL_FADD comp17_55 (
    .a(1'b0),
    .b(sum_16[55]),
    .c(cout_17[54]),
    .cout(cout_17[55]),
    .sum(sum_17[55]));
  AL_FADD comp17_56 (
    .a(1'b0),
    .b(sum_16[56]),
    .c(cout_17[55]),
    .cout(cout_17[56]),
    .sum(sum_17[56]));
  AL_FADD comp17_57 (
    .a(1'b0),
    .b(sum_16[57]),
    .c(cout_17[56]),
    .cout(cout_17[57]),
    .sum(sum_17[57]));
  AL_FADD comp17_58 (
    .a(1'b0),
    .b(sum_16[58]),
    .c(cout_17[57]),
    .cout(cout_17[58]),
    .sum(sum_17[58]));
  AL_FADD comp17_59 (
    .a(1'b0),
    .b(sum_16[59]),
    .c(cout_17[58]),
    .cout(cout_17[59]),
    .sum(sum_17[59]));
  AL_FADD comp17_6 (
    .a(i17[6]),
    .b(sum_16[6]),
    .c(cout_17[5]),
    .cout(cout_17[6]),
    .sum(sum_17[6]));
  AL_FADD comp17_60 (
    .a(1'b0),
    .b(sum_16[60]),
    .c(cout_17[59]),
    .cout(cout_17[60]),
    .sum(sum_17[60]));
  AL_FADD comp17_61 (
    .a(1'b0),
    .b(sum_16[61]),
    .c(cout_17[60]),
    .cout(cout_17[61]),
    .sum(sum_17[61]));
  AL_FADD comp17_62 (
    .a(1'b0),
    .b(sum_16[62]),
    .c(cout_17[61]),
    .cout(cout_17[62]),
    .sum(sum_17[62]));
  AL_FADD comp17_63 (
    .a(1'b0),
    .b(sum_16[63]),
    .c(cout_17[62]),
    .cout(cout_17[63]),
    .sum(sum_17[63]));
  AL_FADD comp17_7 (
    .a(i17[7]),
    .b(sum_16[7]),
    .c(cout_17[6]),
    .cout(cout_17[7]),
    .sum(sum_17[7]));
  AL_FADD comp17_8 (
    .a(i17[8]),
    .b(sum_16[8]),
    .c(cout_17[7]),
    .cout(cout_17[8]),
    .sum(sum_17[8]));
  AL_FADD comp17_9 (
    .a(i17[9]),
    .b(sum_16[9]),
    .c(cout_17[8]),
    .cout(cout_17[9]),
    .sum(sum_17[9]));
  AL_FADD comp18_0 (
    .a(i18[0]),
    .b(sum_17[0]),
    .c(1'b0),
    .cout(cout_18[0]),
    .sum(sum_18[0]));
  AL_FADD comp18_1 (
    .a(i18[1]),
    .b(sum_17[1]),
    .c(cout_18[0]),
    .cout(cout_18[1]),
    .sum(sum_18[1]));
  AL_FADD comp18_10 (
    .a(i18[10]),
    .b(sum_17[10]),
    .c(cout_18[9]),
    .cout(cout_18[10]),
    .sum(sum_18[10]));
  AL_FADD comp18_11 (
    .a(i18[11]),
    .b(sum_17[11]),
    .c(cout_18[10]),
    .cout(cout_18[11]),
    .sum(sum_18[11]));
  AL_FADD comp18_12 (
    .a(i18[12]),
    .b(sum_17[12]),
    .c(cout_18[11]),
    .cout(cout_18[12]),
    .sum(sum_18[12]));
  AL_FADD comp18_13 (
    .a(i18[13]),
    .b(sum_17[13]),
    .c(cout_18[12]),
    .cout(cout_18[13]),
    .sum(sum_18[13]));
  AL_FADD comp18_14 (
    .a(i18[14]),
    .b(sum_17[14]),
    .c(cout_18[13]),
    .cout(cout_18[14]),
    .sum(sum_18[14]));
  AL_FADD comp18_15 (
    .a(i18[15]),
    .b(sum_17[15]),
    .c(cout_18[14]),
    .cout(cout_18[15]),
    .sum(sum_18[15]));
  AL_FADD comp18_16 (
    .a(i18[16]),
    .b(sum_17[16]),
    .c(cout_18[15]),
    .cout(cout_18[16]),
    .sum(sum_18[16]));
  AL_FADD comp18_17 (
    .a(i18[17]),
    .b(sum_17[17]),
    .c(cout_18[16]),
    .cout(cout_18[17]),
    .sum(sum_18[17]));
  AL_FADD comp18_18 (
    .a(i18[18]),
    .b(sum_17[18]),
    .c(cout_18[17]),
    .cout(cout_18[18]),
    .sum(sum_18[18]));
  AL_FADD comp18_19 (
    .a(i18[19]),
    .b(sum_17[19]),
    .c(cout_18[18]),
    .cout(cout_18[19]),
    .sum(sum_18[19]));
  AL_FADD comp18_2 (
    .a(i18[2]),
    .b(sum_17[2]),
    .c(cout_18[1]),
    .cout(cout_18[2]),
    .sum(sum_18[2]));
  AL_FADD comp18_20 (
    .a(i18[20]),
    .b(sum_17[20]),
    .c(cout_18[19]),
    .cout(cout_18[20]),
    .sum(sum_18[20]));
  AL_FADD comp18_21 (
    .a(i18[21]),
    .b(sum_17[21]),
    .c(cout_18[20]),
    .cout(cout_18[21]),
    .sum(sum_18[21]));
  AL_FADD comp18_22 (
    .a(i18[22]),
    .b(sum_17[22]),
    .c(cout_18[21]),
    .cout(cout_18[22]),
    .sum(sum_18[22]));
  AL_FADD comp18_23 (
    .a(i18[23]),
    .b(sum_17[23]),
    .c(cout_18[22]),
    .cout(cout_18[23]),
    .sum(sum_18[23]));
  AL_FADD comp18_24 (
    .a(i18[24]),
    .b(sum_17[24]),
    .c(cout_18[23]),
    .cout(cout_18[24]),
    .sum(sum_18[24]));
  AL_FADD comp18_25 (
    .a(i18[25]),
    .b(sum_17[25]),
    .c(cout_18[24]),
    .cout(cout_18[25]),
    .sum(sum_18[25]));
  AL_FADD comp18_26 (
    .a(i18[26]),
    .b(sum_17[26]),
    .c(cout_18[25]),
    .cout(cout_18[26]),
    .sum(sum_18[26]));
  AL_FADD comp18_27 (
    .a(i18[27]),
    .b(sum_17[27]),
    .c(cout_18[26]),
    .cout(cout_18[27]),
    .sum(sum_18[27]));
  AL_FADD comp18_28 (
    .a(i18[28]),
    .b(sum_17[28]),
    .c(cout_18[27]),
    .cout(cout_18[28]),
    .sum(sum_18[28]));
  AL_FADD comp18_29 (
    .a(i18[29]),
    .b(sum_17[29]),
    .c(cout_18[28]),
    .cout(cout_18[29]),
    .sum(sum_18[29]));
  AL_FADD comp18_3 (
    .a(i18[3]),
    .b(sum_17[3]),
    .c(cout_18[2]),
    .cout(cout_18[3]),
    .sum(sum_18[3]));
  AL_FADD comp18_30 (
    .a(i18[30]),
    .b(sum_17[30]),
    .c(cout_18[29]),
    .cout(cout_18[30]),
    .sum(sum_18[30]));
  AL_FADD comp18_31 (
    .a(i18[31]),
    .b(sum_17[31]),
    .c(cout_18[30]),
    .cout(cout_18[31]),
    .sum(sum_18[31]));
  AL_FADD comp18_32 (
    .a(i18[32]),
    .b(sum_17[32]),
    .c(cout_18[31]),
    .cout(cout_18[32]),
    .sum(sum_18[32]));
  AL_FADD comp18_33 (
    .a(i18[33]),
    .b(sum_17[33]),
    .c(cout_18[32]),
    .cout(cout_18[33]),
    .sum(sum_18[33]));
  AL_FADD comp18_34 (
    .a(i18[34]),
    .b(sum_17[34]),
    .c(cout_18[33]),
    .cout(cout_18[34]),
    .sum(sum_18[34]));
  AL_FADD comp18_35 (
    .a(i18[35]),
    .b(sum_17[35]),
    .c(cout_18[34]),
    .cout(cout_18[35]),
    .sum(sum_18[35]));
  AL_FADD comp18_36 (
    .a(i18[36]),
    .b(sum_17[36]),
    .c(cout_18[35]),
    .cout(cout_18[36]),
    .sum(sum_18[36]));
  AL_FADD comp18_37 (
    .a(i18[37]),
    .b(sum_17[37]),
    .c(cout_18[36]),
    .cout(cout_18[37]),
    .sum(sum_18[37]));
  AL_FADD comp18_38 (
    .a(i18[38]),
    .b(sum_17[38]),
    .c(cout_18[37]),
    .cout(cout_18[38]),
    .sum(sum_18[38]));
  AL_FADD comp18_39 (
    .a(i18[39]),
    .b(sum_17[39]),
    .c(cout_18[38]),
    .cout(cout_18[39]),
    .sum(sum_18[39]));
  AL_FADD comp18_4 (
    .a(i18[4]),
    .b(sum_17[4]),
    .c(cout_18[3]),
    .cout(cout_18[4]),
    .sum(sum_18[4]));
  AL_FADD comp18_40 (
    .a(i18[40]),
    .b(sum_17[40]),
    .c(cout_18[39]),
    .cout(cout_18[40]),
    .sum(sum_18[40]));
  AL_FADD comp18_41 (
    .a(i18[41]),
    .b(sum_17[41]),
    .c(cout_18[40]),
    .cout(cout_18[41]),
    .sum(sum_18[41]));
  AL_FADD comp18_42 (
    .a(i18[42]),
    .b(sum_17[42]),
    .c(cout_18[41]),
    .cout(cout_18[42]),
    .sum(sum_18[42]));
  AL_FADD comp18_43 (
    .a(i18[43]),
    .b(sum_17[43]),
    .c(cout_18[42]),
    .cout(cout_18[43]),
    .sum(sum_18[43]));
  AL_FADD comp18_44 (
    .a(i18[44]),
    .b(sum_17[44]),
    .c(cout_18[43]),
    .cout(cout_18[44]),
    .sum(sum_18[44]));
  AL_FADD comp18_45 (
    .a(1'b0),
    .b(sum_17[45]),
    .c(cout_18[44]),
    .cout(cout_18[45]),
    .sum(sum_18[45]));
  AL_FADD comp18_46 (
    .a(1'b0),
    .b(sum_17[46]),
    .c(cout_18[45]),
    .cout(cout_18[46]),
    .sum(sum_18[46]));
  AL_FADD comp18_47 (
    .a(1'b0),
    .b(sum_17[47]),
    .c(cout_18[46]),
    .cout(cout_18[47]),
    .sum(sum_18[47]));
  AL_FADD comp18_48 (
    .a(1'b0),
    .b(sum_17[48]),
    .c(cout_18[47]),
    .cout(cout_18[48]),
    .sum(sum_18[48]));
  AL_FADD comp18_49 (
    .a(1'b0),
    .b(sum_17[49]),
    .c(cout_18[48]),
    .cout(cout_18[49]),
    .sum(sum_18[49]));
  AL_FADD comp18_5 (
    .a(i18[5]),
    .b(sum_17[5]),
    .c(cout_18[4]),
    .cout(cout_18[5]),
    .sum(sum_18[5]));
  AL_FADD comp18_50 (
    .a(1'b0),
    .b(sum_17[50]),
    .c(cout_18[49]),
    .cout(cout_18[50]),
    .sum(sum_18[50]));
  AL_FADD comp18_51 (
    .a(1'b0),
    .b(sum_17[51]),
    .c(cout_18[50]),
    .cout(cout_18[51]),
    .sum(sum_18[51]));
  AL_FADD comp18_52 (
    .a(1'b0),
    .b(sum_17[52]),
    .c(cout_18[51]),
    .cout(cout_18[52]),
    .sum(sum_18[52]));
  AL_FADD comp18_53 (
    .a(1'b0),
    .b(sum_17[53]),
    .c(cout_18[52]),
    .cout(cout_18[53]),
    .sum(sum_18[53]));
  AL_FADD comp18_54 (
    .a(1'b0),
    .b(sum_17[54]),
    .c(cout_18[53]),
    .cout(cout_18[54]),
    .sum(sum_18[54]));
  AL_FADD comp18_55 (
    .a(1'b0),
    .b(sum_17[55]),
    .c(cout_18[54]),
    .cout(cout_18[55]),
    .sum(sum_18[55]));
  AL_FADD comp18_56 (
    .a(1'b0),
    .b(sum_17[56]),
    .c(cout_18[55]),
    .cout(cout_18[56]),
    .sum(sum_18[56]));
  AL_FADD comp18_57 (
    .a(1'b0),
    .b(sum_17[57]),
    .c(cout_18[56]),
    .cout(cout_18[57]),
    .sum(sum_18[57]));
  AL_FADD comp18_58 (
    .a(1'b0),
    .b(sum_17[58]),
    .c(cout_18[57]),
    .cout(cout_18[58]),
    .sum(sum_18[58]));
  AL_FADD comp18_59 (
    .a(1'b0),
    .b(sum_17[59]),
    .c(cout_18[58]),
    .cout(cout_18[59]),
    .sum(sum_18[59]));
  AL_FADD comp18_6 (
    .a(i18[6]),
    .b(sum_17[6]),
    .c(cout_18[5]),
    .cout(cout_18[6]),
    .sum(sum_18[6]));
  AL_FADD comp18_60 (
    .a(1'b0),
    .b(sum_17[60]),
    .c(cout_18[59]),
    .cout(cout_18[60]),
    .sum(sum_18[60]));
  AL_FADD comp18_61 (
    .a(1'b0),
    .b(sum_17[61]),
    .c(cout_18[60]),
    .cout(cout_18[61]),
    .sum(sum_18[61]));
  AL_FADD comp18_62 (
    .a(1'b0),
    .b(sum_17[62]),
    .c(cout_18[61]),
    .cout(cout_18[62]),
    .sum(sum_18[62]));
  AL_FADD comp18_63 (
    .a(1'b0),
    .b(sum_17[63]),
    .c(cout_18[62]),
    .cout(cout_18[63]),
    .sum(sum_18[63]));
  AL_FADD comp18_7 (
    .a(i18[7]),
    .b(sum_17[7]),
    .c(cout_18[6]),
    .cout(cout_18[7]),
    .sum(sum_18[7]));
  AL_FADD comp18_8 (
    .a(i18[8]),
    .b(sum_17[8]),
    .c(cout_18[7]),
    .cout(cout_18[8]),
    .sum(sum_18[8]));
  AL_FADD comp18_9 (
    .a(i18[9]),
    .b(sum_17[9]),
    .c(cout_18[8]),
    .cout(cout_18[9]),
    .sum(sum_18[9]));
  AL_FADD comp19_0 (
    .a(i19[0]),
    .b(sum_18[0]),
    .c(1'b0),
    .cout(cout_19[0]),
    .sum(sum_19[0]));
  AL_FADD comp19_1 (
    .a(i19[1]),
    .b(sum_18[1]),
    .c(cout_19[0]),
    .cout(cout_19[1]),
    .sum(sum_19[1]));
  AL_FADD comp19_10 (
    .a(i19[10]),
    .b(sum_18[10]),
    .c(cout_19[9]),
    .cout(cout_19[10]),
    .sum(sum_19[10]));
  AL_FADD comp19_11 (
    .a(i19[11]),
    .b(sum_18[11]),
    .c(cout_19[10]),
    .cout(cout_19[11]),
    .sum(sum_19[11]));
  AL_FADD comp19_12 (
    .a(i19[12]),
    .b(sum_18[12]),
    .c(cout_19[11]),
    .cout(cout_19[12]),
    .sum(sum_19[12]));
  AL_FADD comp19_13 (
    .a(i19[13]),
    .b(sum_18[13]),
    .c(cout_19[12]),
    .cout(cout_19[13]),
    .sum(sum_19[13]));
  AL_FADD comp19_14 (
    .a(i19[14]),
    .b(sum_18[14]),
    .c(cout_19[13]),
    .cout(cout_19[14]),
    .sum(sum_19[14]));
  AL_FADD comp19_15 (
    .a(i19[15]),
    .b(sum_18[15]),
    .c(cout_19[14]),
    .cout(cout_19[15]),
    .sum(sum_19[15]));
  AL_FADD comp19_16 (
    .a(i19[16]),
    .b(sum_18[16]),
    .c(cout_19[15]),
    .cout(cout_19[16]),
    .sum(sum_19[16]));
  AL_FADD comp19_17 (
    .a(i19[17]),
    .b(sum_18[17]),
    .c(cout_19[16]),
    .cout(cout_19[17]),
    .sum(sum_19[17]));
  AL_FADD comp19_18 (
    .a(i19[18]),
    .b(sum_18[18]),
    .c(cout_19[17]),
    .cout(cout_19[18]),
    .sum(sum_19[18]));
  AL_FADD comp19_19 (
    .a(i19[19]),
    .b(sum_18[19]),
    .c(cout_19[18]),
    .cout(cout_19[19]),
    .sum(sum_19[19]));
  AL_FADD comp19_2 (
    .a(i19[2]),
    .b(sum_18[2]),
    .c(cout_19[1]),
    .cout(cout_19[2]),
    .sum(sum_19[2]));
  AL_FADD comp19_20 (
    .a(i19[20]),
    .b(sum_18[20]),
    .c(cout_19[19]),
    .cout(cout_19[20]),
    .sum(sum_19[20]));
  AL_FADD comp19_21 (
    .a(i19[21]),
    .b(sum_18[21]),
    .c(cout_19[20]),
    .cout(cout_19[21]),
    .sum(sum_19[21]));
  AL_FADD comp19_22 (
    .a(i19[22]),
    .b(sum_18[22]),
    .c(cout_19[21]),
    .cout(cout_19[22]),
    .sum(sum_19[22]));
  AL_FADD comp19_23 (
    .a(i19[23]),
    .b(sum_18[23]),
    .c(cout_19[22]),
    .cout(cout_19[23]),
    .sum(sum_19[23]));
  AL_FADD comp19_24 (
    .a(i19[24]),
    .b(sum_18[24]),
    .c(cout_19[23]),
    .cout(cout_19[24]),
    .sum(sum_19[24]));
  AL_FADD comp19_25 (
    .a(i19[25]),
    .b(sum_18[25]),
    .c(cout_19[24]),
    .cout(cout_19[25]),
    .sum(sum_19[25]));
  AL_FADD comp19_26 (
    .a(i19[26]),
    .b(sum_18[26]),
    .c(cout_19[25]),
    .cout(cout_19[26]),
    .sum(sum_19[26]));
  AL_FADD comp19_27 (
    .a(i19[27]),
    .b(sum_18[27]),
    .c(cout_19[26]),
    .cout(cout_19[27]),
    .sum(sum_19[27]));
  AL_FADD comp19_28 (
    .a(i19[28]),
    .b(sum_18[28]),
    .c(cout_19[27]),
    .cout(cout_19[28]),
    .sum(sum_19[28]));
  AL_FADD comp19_29 (
    .a(i19[29]),
    .b(sum_18[29]),
    .c(cout_19[28]),
    .cout(cout_19[29]),
    .sum(sum_19[29]));
  AL_FADD comp19_3 (
    .a(i19[3]),
    .b(sum_18[3]),
    .c(cout_19[2]),
    .cout(cout_19[3]),
    .sum(sum_19[3]));
  AL_FADD comp19_30 (
    .a(i19[30]),
    .b(sum_18[30]),
    .c(cout_19[29]),
    .cout(cout_19[30]),
    .sum(sum_19[30]));
  AL_FADD comp19_31 (
    .a(i19[31]),
    .b(sum_18[31]),
    .c(cout_19[30]),
    .cout(cout_19[31]),
    .sum(sum_19[31]));
  AL_FADD comp19_32 (
    .a(i19[32]),
    .b(sum_18[32]),
    .c(cout_19[31]),
    .cout(cout_19[32]),
    .sum(sum_19[32]));
  AL_FADD comp19_33 (
    .a(i19[33]),
    .b(sum_18[33]),
    .c(cout_19[32]),
    .cout(cout_19[33]),
    .sum(sum_19[33]));
  AL_FADD comp19_34 (
    .a(i19[34]),
    .b(sum_18[34]),
    .c(cout_19[33]),
    .cout(cout_19[34]),
    .sum(sum_19[34]));
  AL_FADD comp19_35 (
    .a(i19[35]),
    .b(sum_18[35]),
    .c(cout_19[34]),
    .cout(cout_19[35]),
    .sum(sum_19[35]));
  AL_FADD comp19_36 (
    .a(i19[36]),
    .b(sum_18[36]),
    .c(cout_19[35]),
    .cout(cout_19[36]),
    .sum(sum_19[36]));
  AL_FADD comp19_37 (
    .a(i19[37]),
    .b(sum_18[37]),
    .c(cout_19[36]),
    .cout(cout_19[37]),
    .sum(sum_19[37]));
  AL_FADD comp19_38 (
    .a(i19[38]),
    .b(sum_18[38]),
    .c(cout_19[37]),
    .cout(cout_19[38]),
    .sum(sum_19[38]));
  AL_FADD comp19_39 (
    .a(i19[39]),
    .b(sum_18[39]),
    .c(cout_19[38]),
    .cout(cout_19[39]),
    .sum(sum_19[39]));
  AL_FADD comp19_4 (
    .a(i19[4]),
    .b(sum_18[4]),
    .c(cout_19[3]),
    .cout(cout_19[4]),
    .sum(sum_19[4]));
  AL_FADD comp19_40 (
    .a(i19[40]),
    .b(sum_18[40]),
    .c(cout_19[39]),
    .cout(cout_19[40]),
    .sum(sum_19[40]));
  AL_FADD comp19_41 (
    .a(i19[41]),
    .b(sum_18[41]),
    .c(cout_19[40]),
    .cout(cout_19[41]),
    .sum(sum_19[41]));
  AL_FADD comp19_42 (
    .a(i19[42]),
    .b(sum_18[42]),
    .c(cout_19[41]),
    .cout(cout_19[42]),
    .sum(sum_19[42]));
  AL_FADD comp19_43 (
    .a(i19[43]),
    .b(sum_18[43]),
    .c(cout_19[42]),
    .cout(cout_19[43]),
    .sum(sum_19[43]));
  AL_FADD comp19_44 (
    .a(1'b0),
    .b(sum_18[44]),
    .c(cout_19[43]),
    .cout(cout_19[44]),
    .sum(sum_19[44]));
  AL_FADD comp19_45 (
    .a(1'b0),
    .b(sum_18[45]),
    .c(cout_19[44]),
    .cout(cout_19[45]),
    .sum(sum_19[45]));
  AL_FADD comp19_46 (
    .a(1'b0),
    .b(sum_18[46]),
    .c(cout_19[45]),
    .cout(cout_19[46]),
    .sum(sum_19[46]));
  AL_FADD comp19_47 (
    .a(1'b0),
    .b(sum_18[47]),
    .c(cout_19[46]),
    .cout(cout_19[47]),
    .sum(sum_19[47]));
  AL_FADD comp19_48 (
    .a(1'b0),
    .b(sum_18[48]),
    .c(cout_19[47]),
    .cout(cout_19[48]),
    .sum(sum_19[48]));
  AL_FADD comp19_49 (
    .a(1'b0),
    .b(sum_18[49]),
    .c(cout_19[48]),
    .cout(cout_19[49]),
    .sum(sum_19[49]));
  AL_FADD comp19_5 (
    .a(i19[5]),
    .b(sum_18[5]),
    .c(cout_19[4]),
    .cout(cout_19[5]),
    .sum(sum_19[5]));
  AL_FADD comp19_50 (
    .a(1'b0),
    .b(sum_18[50]),
    .c(cout_19[49]),
    .cout(cout_19[50]),
    .sum(sum_19[50]));
  AL_FADD comp19_51 (
    .a(1'b0),
    .b(sum_18[51]),
    .c(cout_19[50]),
    .cout(cout_19[51]),
    .sum(sum_19[51]));
  AL_FADD comp19_52 (
    .a(1'b0),
    .b(sum_18[52]),
    .c(cout_19[51]),
    .cout(cout_19[52]),
    .sum(sum_19[52]));
  AL_FADD comp19_53 (
    .a(1'b0),
    .b(sum_18[53]),
    .c(cout_19[52]),
    .cout(cout_19[53]),
    .sum(sum_19[53]));
  AL_FADD comp19_54 (
    .a(1'b0),
    .b(sum_18[54]),
    .c(cout_19[53]),
    .cout(cout_19[54]),
    .sum(sum_19[54]));
  AL_FADD comp19_55 (
    .a(1'b0),
    .b(sum_18[55]),
    .c(cout_19[54]),
    .cout(cout_19[55]),
    .sum(sum_19[55]));
  AL_FADD comp19_56 (
    .a(1'b0),
    .b(sum_18[56]),
    .c(cout_19[55]),
    .cout(cout_19[56]),
    .sum(sum_19[56]));
  AL_FADD comp19_57 (
    .a(1'b0),
    .b(sum_18[57]),
    .c(cout_19[56]),
    .cout(cout_19[57]),
    .sum(sum_19[57]));
  AL_FADD comp19_58 (
    .a(1'b0),
    .b(sum_18[58]),
    .c(cout_19[57]),
    .cout(cout_19[58]),
    .sum(sum_19[58]));
  AL_FADD comp19_59 (
    .a(1'b0),
    .b(sum_18[59]),
    .c(cout_19[58]),
    .cout(cout_19[59]),
    .sum(sum_19[59]));
  AL_FADD comp19_6 (
    .a(i19[6]),
    .b(sum_18[6]),
    .c(cout_19[5]),
    .cout(cout_19[6]),
    .sum(sum_19[6]));
  AL_FADD comp19_60 (
    .a(1'b0),
    .b(sum_18[60]),
    .c(cout_19[59]),
    .cout(cout_19[60]),
    .sum(sum_19[60]));
  AL_FADD comp19_61 (
    .a(1'b0),
    .b(sum_18[61]),
    .c(cout_19[60]),
    .cout(cout_19[61]),
    .sum(sum_19[61]));
  AL_FADD comp19_62 (
    .a(1'b0),
    .b(sum_18[62]),
    .c(cout_19[61]),
    .cout(cout_19[62]),
    .sum(sum_19[62]));
  AL_FADD comp19_63 (
    .a(1'b0),
    .b(sum_18[63]),
    .c(cout_19[62]),
    .cout(cout_19[63]),
    .sum(sum_19[63]));
  AL_FADD comp19_7 (
    .a(i19[7]),
    .b(sum_18[7]),
    .c(cout_19[6]),
    .cout(cout_19[7]),
    .sum(sum_19[7]));
  AL_FADD comp19_8 (
    .a(i19[8]),
    .b(sum_18[8]),
    .c(cout_19[7]),
    .cout(cout_19[8]),
    .sum(sum_19[8]));
  AL_FADD comp19_9 (
    .a(i19[9]),
    .b(sum_18[9]),
    .c(cout_19[8]),
    .cout(cout_19[9]),
    .sum(sum_19[9]));
  AL_FADD comp1_0 (
    .a(i1[0]),
    .b(i0[0]),
    .c(1'b0),
    .cout(cout_1[0]),
    .sum(sum_1[0]));
  AL_FADD comp1_1 (
    .a(i1[1]),
    .b(i0[1]),
    .c(cout_1[0]),
    .cout(cout_1[1]),
    .sum(sum_1[1]));
  AL_FADD comp1_10 (
    .a(i1[10]),
    .b(i0[10]),
    .c(cout_1[9]),
    .cout(cout_1[10]),
    .sum(sum_1[10]));
  AL_FADD comp1_11 (
    .a(i1[11]),
    .b(i0[11]),
    .c(cout_1[10]),
    .cout(cout_1[11]),
    .sum(sum_1[11]));
  AL_FADD comp1_12 (
    .a(i1[12]),
    .b(i0[12]),
    .c(cout_1[11]),
    .cout(cout_1[12]),
    .sum(sum_1[12]));
  AL_FADD comp1_13 (
    .a(i1[13]),
    .b(i0[13]),
    .c(cout_1[12]),
    .cout(cout_1[13]),
    .sum(sum_1[13]));
  AL_FADD comp1_14 (
    .a(i1[14]),
    .b(i0[14]),
    .c(cout_1[13]),
    .cout(cout_1[14]),
    .sum(sum_1[14]));
  AL_FADD comp1_15 (
    .a(i1[15]),
    .b(i0[15]),
    .c(cout_1[14]),
    .cout(cout_1[15]),
    .sum(sum_1[15]));
  AL_FADD comp1_16 (
    .a(i1[16]),
    .b(i0[16]),
    .c(cout_1[15]),
    .cout(cout_1[16]),
    .sum(sum_1[16]));
  AL_FADD comp1_17 (
    .a(i1[17]),
    .b(i0[17]),
    .c(cout_1[16]),
    .cout(cout_1[17]),
    .sum(sum_1[17]));
  AL_FADD comp1_18 (
    .a(i1[18]),
    .b(i0[18]),
    .c(cout_1[17]),
    .cout(cout_1[18]),
    .sum(sum_1[18]));
  AL_FADD comp1_19 (
    .a(i1[19]),
    .b(i0[19]),
    .c(cout_1[18]),
    .cout(cout_1[19]),
    .sum(sum_1[19]));
  AL_FADD comp1_2 (
    .a(i1[2]),
    .b(i0[2]),
    .c(cout_1[1]),
    .cout(cout_1[2]),
    .sum(sum_1[2]));
  AL_FADD comp1_20 (
    .a(i1[20]),
    .b(i0[20]),
    .c(cout_1[19]),
    .cout(cout_1[20]),
    .sum(sum_1[20]));
  AL_FADD comp1_21 (
    .a(i1[21]),
    .b(i0[21]),
    .c(cout_1[20]),
    .cout(cout_1[21]),
    .sum(sum_1[21]));
  AL_FADD comp1_22 (
    .a(i1[22]),
    .b(i0[22]),
    .c(cout_1[21]),
    .cout(cout_1[22]),
    .sum(sum_1[22]));
  AL_FADD comp1_23 (
    .a(i1[23]),
    .b(i0[23]),
    .c(cout_1[22]),
    .cout(cout_1[23]),
    .sum(sum_1[23]));
  AL_FADD comp1_24 (
    .a(i1[24]),
    .b(i0[24]),
    .c(cout_1[23]),
    .cout(cout_1[24]),
    .sum(sum_1[24]));
  AL_FADD comp1_25 (
    .a(i1[25]),
    .b(i0[25]),
    .c(cout_1[24]),
    .cout(cout_1[25]),
    .sum(sum_1[25]));
  AL_FADD comp1_26 (
    .a(i1[26]),
    .b(i0[26]),
    .c(cout_1[25]),
    .cout(cout_1[26]),
    .sum(sum_1[26]));
  AL_FADD comp1_27 (
    .a(i1[27]),
    .b(i0[27]),
    .c(cout_1[26]),
    .cout(cout_1[27]),
    .sum(sum_1[27]));
  AL_FADD comp1_28 (
    .a(i1[28]),
    .b(i0[28]),
    .c(cout_1[27]),
    .cout(cout_1[28]),
    .sum(sum_1[28]));
  AL_FADD comp1_29 (
    .a(i1[29]),
    .b(i0[29]),
    .c(cout_1[28]),
    .cout(cout_1[29]),
    .sum(sum_1[29]));
  AL_FADD comp1_3 (
    .a(i1[3]),
    .b(i0[3]),
    .c(cout_1[2]),
    .cout(cout_1[3]),
    .sum(sum_1[3]));
  AL_FADD comp1_30 (
    .a(i1[30]),
    .b(i0[30]),
    .c(cout_1[29]),
    .cout(cout_1[30]),
    .sum(sum_1[30]));
  AL_FADD comp1_31 (
    .a(i1[31]),
    .b(i0[31]),
    .c(cout_1[30]),
    .cout(cout_1[31]),
    .sum(sum_1[31]));
  AL_FADD comp1_32 (
    .a(i1[32]),
    .b(i0[32]),
    .c(cout_1[31]),
    .cout(cout_1[32]),
    .sum(sum_1[32]));
  AL_FADD comp1_33 (
    .a(i1[33]),
    .b(i0[33]),
    .c(cout_1[32]),
    .cout(cout_1[33]),
    .sum(sum_1[33]));
  AL_FADD comp1_34 (
    .a(i1[34]),
    .b(i0[34]),
    .c(cout_1[33]),
    .cout(cout_1[34]),
    .sum(sum_1[34]));
  AL_FADD comp1_35 (
    .a(i1[35]),
    .b(i0[35]),
    .c(cout_1[34]),
    .cout(cout_1[35]),
    .sum(sum_1[35]));
  AL_FADD comp1_36 (
    .a(i1[36]),
    .b(i0[36]),
    .c(cout_1[35]),
    .cout(cout_1[36]),
    .sum(sum_1[36]));
  AL_FADD comp1_37 (
    .a(i1[37]),
    .b(i0[37]),
    .c(cout_1[36]),
    .cout(cout_1[37]),
    .sum(sum_1[37]));
  AL_FADD comp1_38 (
    .a(i1[38]),
    .b(i0[38]),
    .c(cout_1[37]),
    .cout(cout_1[38]),
    .sum(sum_1[38]));
  AL_FADD comp1_39 (
    .a(i1[39]),
    .b(i0[39]),
    .c(cout_1[38]),
    .cout(cout_1[39]),
    .sum(sum_1[39]));
  AL_FADD comp1_4 (
    .a(i1[4]),
    .b(i0[4]),
    .c(cout_1[3]),
    .cout(cout_1[4]),
    .sum(sum_1[4]));
  AL_FADD comp1_40 (
    .a(i1[40]),
    .b(i0[40]),
    .c(cout_1[39]),
    .cout(cout_1[40]),
    .sum(sum_1[40]));
  AL_FADD comp1_41 (
    .a(i1[41]),
    .b(i0[41]),
    .c(cout_1[40]),
    .cout(cout_1[41]),
    .sum(sum_1[41]));
  AL_FADD comp1_42 (
    .a(i1[42]),
    .b(i0[42]),
    .c(cout_1[41]),
    .cout(cout_1[42]),
    .sum(sum_1[42]));
  AL_FADD comp1_43 (
    .a(i1[43]),
    .b(i0[43]),
    .c(cout_1[42]),
    .cout(cout_1[43]),
    .sum(sum_1[43]));
  AL_FADD comp1_44 (
    .a(i1[44]),
    .b(i0[44]),
    .c(cout_1[43]),
    .cout(cout_1[44]),
    .sum(sum_1[44]));
  AL_FADD comp1_45 (
    .a(i1[45]),
    .b(i0[45]),
    .c(cout_1[44]),
    .cout(cout_1[45]),
    .sum(sum_1[45]));
  AL_FADD comp1_46 (
    .a(i1[46]),
    .b(i0[46]),
    .c(cout_1[45]),
    .cout(cout_1[46]),
    .sum(sum_1[46]));
  AL_FADD comp1_47 (
    .a(i1[47]),
    .b(i0[47]),
    .c(cout_1[46]),
    .cout(cout_1[47]),
    .sum(sum_1[47]));
  AL_FADD comp1_48 (
    .a(i1[48]),
    .b(i0[48]),
    .c(cout_1[47]),
    .cout(cout_1[48]),
    .sum(sum_1[48]));
  AL_FADD comp1_49 (
    .a(i1[49]),
    .b(i0[49]),
    .c(cout_1[48]),
    .cout(cout_1[49]),
    .sum(sum_1[49]));
  AL_FADD comp1_5 (
    .a(i1[5]),
    .b(i0[5]),
    .c(cout_1[4]),
    .cout(cout_1[5]),
    .sum(sum_1[5]));
  AL_FADD comp1_50 (
    .a(i1[50]),
    .b(i0[50]),
    .c(cout_1[49]),
    .cout(cout_1[50]),
    .sum(sum_1[50]));
  AL_FADD comp1_51 (
    .a(i1[51]),
    .b(i0[51]),
    .c(cout_1[50]),
    .cout(cout_1[51]),
    .sum(sum_1[51]));
  AL_FADD comp1_52 (
    .a(i1[52]),
    .b(i0[52]),
    .c(cout_1[51]),
    .cout(cout_1[52]),
    .sum(sum_1[52]));
  AL_FADD comp1_53 (
    .a(i1[53]),
    .b(i0[53]),
    .c(cout_1[52]),
    .cout(cout_1[53]),
    .sum(sum_1[53]));
  AL_FADD comp1_54 (
    .a(i1[54]),
    .b(i0[54]),
    .c(cout_1[53]),
    .cout(cout_1[54]),
    .sum(sum_1[54]));
  AL_FADD comp1_55 (
    .a(i1[55]),
    .b(i0[55]),
    .c(cout_1[54]),
    .cout(cout_1[55]),
    .sum(sum_1[55]));
  AL_FADD comp1_56 (
    .a(i1[56]),
    .b(i0[56]),
    .c(cout_1[55]),
    .cout(cout_1[56]),
    .sum(sum_1[56]));
  AL_FADD comp1_57 (
    .a(i1[57]),
    .b(i0[57]),
    .c(cout_1[56]),
    .cout(cout_1[57]),
    .sum(sum_1[57]));
  AL_FADD comp1_58 (
    .a(i1[58]),
    .b(i0[58]),
    .c(cout_1[57]),
    .cout(cout_1[58]),
    .sum(sum_1[58]));
  AL_FADD comp1_59 (
    .a(i1[59]),
    .b(i0[59]),
    .c(cout_1[58]),
    .cout(cout_1[59]),
    .sum(sum_1[59]));
  AL_FADD comp1_6 (
    .a(i1[6]),
    .b(i0[6]),
    .c(cout_1[5]),
    .cout(cout_1[6]),
    .sum(sum_1[6]));
  AL_FADD comp1_60 (
    .a(i1[60]),
    .b(i0[60]),
    .c(cout_1[59]),
    .cout(cout_1[60]),
    .sum(sum_1[60]));
  AL_FADD comp1_61 (
    .a(i1[61]),
    .b(i0[61]),
    .c(cout_1[60]),
    .cout(cout_1[61]),
    .sum(sum_1[61]));
  AL_FADD comp1_62 (
    .a(1'b0),
    .b(i0[62]),
    .c(cout_1[61]),
    .cout(cout_1[62]),
    .sum(sum_1[62]));
  AL_FADD comp1_7 (
    .a(i1[7]),
    .b(i0[7]),
    .c(cout_1[6]),
    .cout(cout_1[7]),
    .sum(sum_1[7]));
  AL_FADD comp1_8 (
    .a(i1[8]),
    .b(i0[8]),
    .c(cout_1[7]),
    .cout(cout_1[8]),
    .sum(sum_1[8]));
  AL_FADD comp1_9 (
    .a(i1[9]),
    .b(i0[9]),
    .c(cout_1[8]),
    .cout(cout_1[9]),
    .sum(sum_1[9]));
  AL_FADD comp20_0 (
    .a(i20[0]),
    .b(sum_19[0]),
    .c(1'b0),
    .cout(cout_20[0]),
    .sum(sum_20[0]));
  AL_FADD comp20_1 (
    .a(i20[1]),
    .b(sum_19[1]),
    .c(cout_20[0]),
    .cout(cout_20[1]),
    .sum(sum_20[1]));
  AL_FADD comp20_10 (
    .a(i20[10]),
    .b(sum_19[10]),
    .c(cout_20[9]),
    .cout(cout_20[10]),
    .sum(sum_20[10]));
  AL_FADD comp20_11 (
    .a(i20[11]),
    .b(sum_19[11]),
    .c(cout_20[10]),
    .cout(cout_20[11]),
    .sum(sum_20[11]));
  AL_FADD comp20_12 (
    .a(i20[12]),
    .b(sum_19[12]),
    .c(cout_20[11]),
    .cout(cout_20[12]),
    .sum(sum_20[12]));
  AL_FADD comp20_13 (
    .a(i20[13]),
    .b(sum_19[13]),
    .c(cout_20[12]),
    .cout(cout_20[13]),
    .sum(sum_20[13]));
  AL_FADD comp20_14 (
    .a(i20[14]),
    .b(sum_19[14]),
    .c(cout_20[13]),
    .cout(cout_20[14]),
    .sum(sum_20[14]));
  AL_FADD comp20_15 (
    .a(i20[15]),
    .b(sum_19[15]),
    .c(cout_20[14]),
    .cout(cout_20[15]),
    .sum(sum_20[15]));
  AL_FADD comp20_16 (
    .a(i20[16]),
    .b(sum_19[16]),
    .c(cout_20[15]),
    .cout(cout_20[16]),
    .sum(sum_20[16]));
  AL_FADD comp20_17 (
    .a(i20[17]),
    .b(sum_19[17]),
    .c(cout_20[16]),
    .cout(cout_20[17]),
    .sum(sum_20[17]));
  AL_FADD comp20_18 (
    .a(i20[18]),
    .b(sum_19[18]),
    .c(cout_20[17]),
    .cout(cout_20[18]),
    .sum(sum_20[18]));
  AL_FADD comp20_19 (
    .a(i20[19]),
    .b(sum_19[19]),
    .c(cout_20[18]),
    .cout(cout_20[19]),
    .sum(sum_20[19]));
  AL_FADD comp20_2 (
    .a(i20[2]),
    .b(sum_19[2]),
    .c(cout_20[1]),
    .cout(cout_20[2]),
    .sum(sum_20[2]));
  AL_FADD comp20_20 (
    .a(i20[20]),
    .b(sum_19[20]),
    .c(cout_20[19]),
    .cout(cout_20[20]),
    .sum(sum_20[20]));
  AL_FADD comp20_21 (
    .a(i20[21]),
    .b(sum_19[21]),
    .c(cout_20[20]),
    .cout(cout_20[21]),
    .sum(sum_20[21]));
  AL_FADD comp20_22 (
    .a(i20[22]),
    .b(sum_19[22]),
    .c(cout_20[21]),
    .cout(cout_20[22]),
    .sum(sum_20[22]));
  AL_FADD comp20_23 (
    .a(i20[23]),
    .b(sum_19[23]),
    .c(cout_20[22]),
    .cout(cout_20[23]),
    .sum(sum_20[23]));
  AL_FADD comp20_24 (
    .a(i20[24]),
    .b(sum_19[24]),
    .c(cout_20[23]),
    .cout(cout_20[24]),
    .sum(sum_20[24]));
  AL_FADD comp20_25 (
    .a(i20[25]),
    .b(sum_19[25]),
    .c(cout_20[24]),
    .cout(cout_20[25]),
    .sum(sum_20[25]));
  AL_FADD comp20_26 (
    .a(i20[26]),
    .b(sum_19[26]),
    .c(cout_20[25]),
    .cout(cout_20[26]),
    .sum(sum_20[26]));
  AL_FADD comp20_27 (
    .a(i20[27]),
    .b(sum_19[27]),
    .c(cout_20[26]),
    .cout(cout_20[27]),
    .sum(sum_20[27]));
  AL_FADD comp20_28 (
    .a(i20[28]),
    .b(sum_19[28]),
    .c(cout_20[27]),
    .cout(cout_20[28]),
    .sum(sum_20[28]));
  AL_FADD comp20_29 (
    .a(i20[29]),
    .b(sum_19[29]),
    .c(cout_20[28]),
    .cout(cout_20[29]),
    .sum(sum_20[29]));
  AL_FADD comp20_3 (
    .a(i20[3]),
    .b(sum_19[3]),
    .c(cout_20[2]),
    .cout(cout_20[3]),
    .sum(sum_20[3]));
  AL_FADD comp20_30 (
    .a(i20[30]),
    .b(sum_19[30]),
    .c(cout_20[29]),
    .cout(cout_20[30]),
    .sum(sum_20[30]));
  AL_FADD comp20_31 (
    .a(i20[31]),
    .b(sum_19[31]),
    .c(cout_20[30]),
    .cout(cout_20[31]),
    .sum(sum_20[31]));
  AL_FADD comp20_32 (
    .a(i20[32]),
    .b(sum_19[32]),
    .c(cout_20[31]),
    .cout(cout_20[32]),
    .sum(sum_20[32]));
  AL_FADD comp20_33 (
    .a(i20[33]),
    .b(sum_19[33]),
    .c(cout_20[32]),
    .cout(cout_20[33]),
    .sum(sum_20[33]));
  AL_FADD comp20_34 (
    .a(i20[34]),
    .b(sum_19[34]),
    .c(cout_20[33]),
    .cout(cout_20[34]),
    .sum(sum_20[34]));
  AL_FADD comp20_35 (
    .a(i20[35]),
    .b(sum_19[35]),
    .c(cout_20[34]),
    .cout(cout_20[35]),
    .sum(sum_20[35]));
  AL_FADD comp20_36 (
    .a(i20[36]),
    .b(sum_19[36]),
    .c(cout_20[35]),
    .cout(cout_20[36]),
    .sum(sum_20[36]));
  AL_FADD comp20_37 (
    .a(i20[37]),
    .b(sum_19[37]),
    .c(cout_20[36]),
    .cout(cout_20[37]),
    .sum(sum_20[37]));
  AL_FADD comp20_38 (
    .a(i20[38]),
    .b(sum_19[38]),
    .c(cout_20[37]),
    .cout(cout_20[38]),
    .sum(sum_20[38]));
  AL_FADD comp20_39 (
    .a(i20[39]),
    .b(sum_19[39]),
    .c(cout_20[38]),
    .cout(cout_20[39]),
    .sum(sum_20[39]));
  AL_FADD comp20_4 (
    .a(i20[4]),
    .b(sum_19[4]),
    .c(cout_20[3]),
    .cout(cout_20[4]),
    .sum(sum_20[4]));
  AL_FADD comp20_40 (
    .a(i20[40]),
    .b(sum_19[40]),
    .c(cout_20[39]),
    .cout(cout_20[40]),
    .sum(sum_20[40]));
  AL_FADD comp20_41 (
    .a(i20[41]),
    .b(sum_19[41]),
    .c(cout_20[40]),
    .cout(cout_20[41]),
    .sum(sum_20[41]));
  AL_FADD comp20_42 (
    .a(i20[42]),
    .b(sum_19[42]),
    .c(cout_20[41]),
    .cout(cout_20[42]),
    .sum(sum_20[42]));
  AL_FADD comp20_43 (
    .a(1'b0),
    .b(sum_19[43]),
    .c(cout_20[42]),
    .cout(cout_20[43]),
    .sum(sum_20[43]));
  AL_FADD comp20_44 (
    .a(1'b0),
    .b(sum_19[44]),
    .c(cout_20[43]),
    .cout(cout_20[44]),
    .sum(sum_20[44]));
  AL_FADD comp20_45 (
    .a(1'b0),
    .b(sum_19[45]),
    .c(cout_20[44]),
    .cout(cout_20[45]),
    .sum(sum_20[45]));
  AL_FADD comp20_46 (
    .a(1'b0),
    .b(sum_19[46]),
    .c(cout_20[45]),
    .cout(cout_20[46]),
    .sum(sum_20[46]));
  AL_FADD comp20_47 (
    .a(1'b0),
    .b(sum_19[47]),
    .c(cout_20[46]),
    .cout(cout_20[47]),
    .sum(sum_20[47]));
  AL_FADD comp20_48 (
    .a(1'b0),
    .b(sum_19[48]),
    .c(cout_20[47]),
    .cout(cout_20[48]),
    .sum(sum_20[48]));
  AL_FADD comp20_49 (
    .a(1'b0),
    .b(sum_19[49]),
    .c(cout_20[48]),
    .cout(cout_20[49]),
    .sum(sum_20[49]));
  AL_FADD comp20_5 (
    .a(i20[5]),
    .b(sum_19[5]),
    .c(cout_20[4]),
    .cout(cout_20[5]),
    .sum(sum_20[5]));
  AL_FADD comp20_50 (
    .a(1'b0),
    .b(sum_19[50]),
    .c(cout_20[49]),
    .cout(cout_20[50]),
    .sum(sum_20[50]));
  AL_FADD comp20_51 (
    .a(1'b0),
    .b(sum_19[51]),
    .c(cout_20[50]),
    .cout(cout_20[51]),
    .sum(sum_20[51]));
  AL_FADD comp20_52 (
    .a(1'b0),
    .b(sum_19[52]),
    .c(cout_20[51]),
    .cout(cout_20[52]),
    .sum(sum_20[52]));
  AL_FADD comp20_53 (
    .a(1'b0),
    .b(sum_19[53]),
    .c(cout_20[52]),
    .cout(cout_20[53]),
    .sum(sum_20[53]));
  AL_FADD comp20_54 (
    .a(1'b0),
    .b(sum_19[54]),
    .c(cout_20[53]),
    .cout(cout_20[54]),
    .sum(sum_20[54]));
  AL_FADD comp20_55 (
    .a(1'b0),
    .b(sum_19[55]),
    .c(cout_20[54]),
    .cout(cout_20[55]),
    .sum(sum_20[55]));
  AL_FADD comp20_56 (
    .a(1'b0),
    .b(sum_19[56]),
    .c(cout_20[55]),
    .cout(cout_20[56]),
    .sum(sum_20[56]));
  AL_FADD comp20_57 (
    .a(1'b0),
    .b(sum_19[57]),
    .c(cout_20[56]),
    .cout(cout_20[57]),
    .sum(sum_20[57]));
  AL_FADD comp20_58 (
    .a(1'b0),
    .b(sum_19[58]),
    .c(cout_20[57]),
    .cout(cout_20[58]),
    .sum(sum_20[58]));
  AL_FADD comp20_59 (
    .a(1'b0),
    .b(sum_19[59]),
    .c(cout_20[58]),
    .cout(cout_20[59]),
    .sum(sum_20[59]));
  AL_FADD comp20_6 (
    .a(i20[6]),
    .b(sum_19[6]),
    .c(cout_20[5]),
    .cout(cout_20[6]),
    .sum(sum_20[6]));
  AL_FADD comp20_60 (
    .a(1'b0),
    .b(sum_19[60]),
    .c(cout_20[59]),
    .cout(cout_20[60]),
    .sum(sum_20[60]));
  AL_FADD comp20_61 (
    .a(1'b0),
    .b(sum_19[61]),
    .c(cout_20[60]),
    .cout(cout_20[61]),
    .sum(sum_20[61]));
  AL_FADD comp20_62 (
    .a(1'b0),
    .b(sum_19[62]),
    .c(cout_20[61]),
    .cout(cout_20[62]),
    .sum(sum_20[62]));
  AL_FADD comp20_63 (
    .a(1'b0),
    .b(sum_19[63]),
    .c(cout_20[62]),
    .cout(cout_20[63]),
    .sum(sum_20[63]));
  AL_FADD comp20_7 (
    .a(i20[7]),
    .b(sum_19[7]),
    .c(cout_20[6]),
    .cout(cout_20[7]),
    .sum(sum_20[7]));
  AL_FADD comp20_8 (
    .a(i20[8]),
    .b(sum_19[8]),
    .c(cout_20[7]),
    .cout(cout_20[8]),
    .sum(sum_20[8]));
  AL_FADD comp20_9 (
    .a(i20[9]),
    .b(sum_19[9]),
    .c(cout_20[8]),
    .cout(cout_20[9]),
    .sum(sum_20[9]));
  AL_FADD comp21_0 (
    .a(i21[0]),
    .b(sum_20[0]),
    .c(1'b0),
    .cout(cout_21[0]),
    .sum(sum_21[0]));
  AL_FADD comp21_1 (
    .a(i21[1]),
    .b(sum_20[1]),
    .c(cout_21[0]),
    .cout(cout_21[1]),
    .sum(sum_21[1]));
  AL_FADD comp21_10 (
    .a(i21[10]),
    .b(sum_20[10]),
    .c(cout_21[9]),
    .cout(cout_21[10]),
    .sum(sum_21[10]));
  AL_FADD comp21_11 (
    .a(i21[11]),
    .b(sum_20[11]),
    .c(cout_21[10]),
    .cout(cout_21[11]),
    .sum(sum_21[11]));
  AL_FADD comp21_12 (
    .a(i21[12]),
    .b(sum_20[12]),
    .c(cout_21[11]),
    .cout(cout_21[12]),
    .sum(sum_21[12]));
  AL_FADD comp21_13 (
    .a(i21[13]),
    .b(sum_20[13]),
    .c(cout_21[12]),
    .cout(cout_21[13]),
    .sum(sum_21[13]));
  AL_FADD comp21_14 (
    .a(i21[14]),
    .b(sum_20[14]),
    .c(cout_21[13]),
    .cout(cout_21[14]),
    .sum(sum_21[14]));
  AL_FADD comp21_15 (
    .a(i21[15]),
    .b(sum_20[15]),
    .c(cout_21[14]),
    .cout(cout_21[15]),
    .sum(sum_21[15]));
  AL_FADD comp21_16 (
    .a(i21[16]),
    .b(sum_20[16]),
    .c(cout_21[15]),
    .cout(cout_21[16]),
    .sum(sum_21[16]));
  AL_FADD comp21_17 (
    .a(i21[17]),
    .b(sum_20[17]),
    .c(cout_21[16]),
    .cout(cout_21[17]),
    .sum(sum_21[17]));
  AL_FADD comp21_18 (
    .a(i21[18]),
    .b(sum_20[18]),
    .c(cout_21[17]),
    .cout(cout_21[18]),
    .sum(sum_21[18]));
  AL_FADD comp21_19 (
    .a(i21[19]),
    .b(sum_20[19]),
    .c(cout_21[18]),
    .cout(cout_21[19]),
    .sum(sum_21[19]));
  AL_FADD comp21_2 (
    .a(i21[2]),
    .b(sum_20[2]),
    .c(cout_21[1]),
    .cout(cout_21[2]),
    .sum(sum_21[2]));
  AL_FADD comp21_20 (
    .a(i21[20]),
    .b(sum_20[20]),
    .c(cout_21[19]),
    .cout(cout_21[20]),
    .sum(sum_21[20]));
  AL_FADD comp21_21 (
    .a(i21[21]),
    .b(sum_20[21]),
    .c(cout_21[20]),
    .cout(cout_21[21]),
    .sum(sum_21[21]));
  AL_FADD comp21_22 (
    .a(i21[22]),
    .b(sum_20[22]),
    .c(cout_21[21]),
    .cout(cout_21[22]),
    .sum(sum_21[22]));
  AL_FADD comp21_23 (
    .a(i21[23]),
    .b(sum_20[23]),
    .c(cout_21[22]),
    .cout(cout_21[23]),
    .sum(sum_21[23]));
  AL_FADD comp21_24 (
    .a(i21[24]),
    .b(sum_20[24]),
    .c(cout_21[23]),
    .cout(cout_21[24]),
    .sum(sum_21[24]));
  AL_FADD comp21_25 (
    .a(i21[25]),
    .b(sum_20[25]),
    .c(cout_21[24]),
    .cout(cout_21[25]),
    .sum(sum_21[25]));
  AL_FADD comp21_26 (
    .a(i21[26]),
    .b(sum_20[26]),
    .c(cout_21[25]),
    .cout(cout_21[26]),
    .sum(sum_21[26]));
  AL_FADD comp21_27 (
    .a(i21[27]),
    .b(sum_20[27]),
    .c(cout_21[26]),
    .cout(cout_21[27]),
    .sum(sum_21[27]));
  AL_FADD comp21_28 (
    .a(i21[28]),
    .b(sum_20[28]),
    .c(cout_21[27]),
    .cout(cout_21[28]),
    .sum(sum_21[28]));
  AL_FADD comp21_29 (
    .a(i21[29]),
    .b(sum_20[29]),
    .c(cout_21[28]),
    .cout(cout_21[29]),
    .sum(sum_21[29]));
  AL_FADD comp21_3 (
    .a(i21[3]),
    .b(sum_20[3]),
    .c(cout_21[2]),
    .cout(cout_21[3]),
    .sum(sum_21[3]));
  AL_FADD comp21_30 (
    .a(i21[30]),
    .b(sum_20[30]),
    .c(cout_21[29]),
    .cout(cout_21[30]),
    .sum(sum_21[30]));
  AL_FADD comp21_31 (
    .a(i21[31]),
    .b(sum_20[31]),
    .c(cout_21[30]),
    .cout(cout_21[31]),
    .sum(sum_21[31]));
  AL_FADD comp21_32 (
    .a(i21[32]),
    .b(sum_20[32]),
    .c(cout_21[31]),
    .cout(cout_21[32]),
    .sum(sum_21[32]));
  AL_FADD comp21_33 (
    .a(i21[33]),
    .b(sum_20[33]),
    .c(cout_21[32]),
    .cout(cout_21[33]),
    .sum(sum_21[33]));
  AL_FADD comp21_34 (
    .a(i21[34]),
    .b(sum_20[34]),
    .c(cout_21[33]),
    .cout(cout_21[34]),
    .sum(sum_21[34]));
  AL_FADD comp21_35 (
    .a(i21[35]),
    .b(sum_20[35]),
    .c(cout_21[34]),
    .cout(cout_21[35]),
    .sum(sum_21[35]));
  AL_FADD comp21_36 (
    .a(i21[36]),
    .b(sum_20[36]),
    .c(cout_21[35]),
    .cout(cout_21[36]),
    .sum(sum_21[36]));
  AL_FADD comp21_37 (
    .a(i21[37]),
    .b(sum_20[37]),
    .c(cout_21[36]),
    .cout(cout_21[37]),
    .sum(sum_21[37]));
  AL_FADD comp21_38 (
    .a(i21[38]),
    .b(sum_20[38]),
    .c(cout_21[37]),
    .cout(cout_21[38]),
    .sum(sum_21[38]));
  AL_FADD comp21_39 (
    .a(i21[39]),
    .b(sum_20[39]),
    .c(cout_21[38]),
    .cout(cout_21[39]),
    .sum(sum_21[39]));
  AL_FADD comp21_4 (
    .a(i21[4]),
    .b(sum_20[4]),
    .c(cout_21[3]),
    .cout(cout_21[4]),
    .sum(sum_21[4]));
  AL_FADD comp21_40 (
    .a(i21[40]),
    .b(sum_20[40]),
    .c(cout_21[39]),
    .cout(cout_21[40]),
    .sum(sum_21[40]));
  AL_FADD comp21_41 (
    .a(i21[41]),
    .b(sum_20[41]),
    .c(cout_21[40]),
    .cout(cout_21[41]),
    .sum(sum_21[41]));
  AL_FADD comp21_42 (
    .a(1'b0),
    .b(sum_20[42]),
    .c(cout_21[41]),
    .cout(cout_21[42]),
    .sum(sum_21[42]));
  AL_FADD comp21_43 (
    .a(1'b0),
    .b(sum_20[43]),
    .c(cout_21[42]),
    .cout(cout_21[43]),
    .sum(sum_21[43]));
  AL_FADD comp21_44 (
    .a(1'b0),
    .b(sum_20[44]),
    .c(cout_21[43]),
    .cout(cout_21[44]),
    .sum(sum_21[44]));
  AL_FADD comp21_45 (
    .a(1'b0),
    .b(sum_20[45]),
    .c(cout_21[44]),
    .cout(cout_21[45]),
    .sum(sum_21[45]));
  AL_FADD comp21_46 (
    .a(1'b0),
    .b(sum_20[46]),
    .c(cout_21[45]),
    .cout(cout_21[46]),
    .sum(sum_21[46]));
  AL_FADD comp21_47 (
    .a(1'b0),
    .b(sum_20[47]),
    .c(cout_21[46]),
    .cout(cout_21[47]),
    .sum(sum_21[47]));
  AL_FADD comp21_48 (
    .a(1'b0),
    .b(sum_20[48]),
    .c(cout_21[47]),
    .cout(cout_21[48]),
    .sum(sum_21[48]));
  AL_FADD comp21_49 (
    .a(1'b0),
    .b(sum_20[49]),
    .c(cout_21[48]),
    .cout(cout_21[49]),
    .sum(sum_21[49]));
  AL_FADD comp21_5 (
    .a(i21[5]),
    .b(sum_20[5]),
    .c(cout_21[4]),
    .cout(cout_21[5]),
    .sum(sum_21[5]));
  AL_FADD comp21_50 (
    .a(1'b0),
    .b(sum_20[50]),
    .c(cout_21[49]),
    .cout(cout_21[50]),
    .sum(sum_21[50]));
  AL_FADD comp21_51 (
    .a(1'b0),
    .b(sum_20[51]),
    .c(cout_21[50]),
    .cout(cout_21[51]),
    .sum(sum_21[51]));
  AL_FADD comp21_52 (
    .a(1'b0),
    .b(sum_20[52]),
    .c(cout_21[51]),
    .cout(cout_21[52]),
    .sum(sum_21[52]));
  AL_FADD comp21_53 (
    .a(1'b0),
    .b(sum_20[53]),
    .c(cout_21[52]),
    .cout(cout_21[53]),
    .sum(sum_21[53]));
  AL_FADD comp21_54 (
    .a(1'b0),
    .b(sum_20[54]),
    .c(cout_21[53]),
    .cout(cout_21[54]),
    .sum(sum_21[54]));
  AL_FADD comp21_55 (
    .a(1'b0),
    .b(sum_20[55]),
    .c(cout_21[54]),
    .cout(cout_21[55]),
    .sum(sum_21[55]));
  AL_FADD comp21_56 (
    .a(1'b0),
    .b(sum_20[56]),
    .c(cout_21[55]),
    .cout(cout_21[56]),
    .sum(sum_21[56]));
  AL_FADD comp21_57 (
    .a(1'b0),
    .b(sum_20[57]),
    .c(cout_21[56]),
    .cout(cout_21[57]),
    .sum(sum_21[57]));
  AL_FADD comp21_58 (
    .a(1'b0),
    .b(sum_20[58]),
    .c(cout_21[57]),
    .cout(cout_21[58]),
    .sum(sum_21[58]));
  AL_FADD comp21_59 (
    .a(1'b0),
    .b(sum_20[59]),
    .c(cout_21[58]),
    .cout(cout_21[59]),
    .sum(sum_21[59]));
  AL_FADD comp21_6 (
    .a(i21[6]),
    .b(sum_20[6]),
    .c(cout_21[5]),
    .cout(cout_21[6]),
    .sum(sum_21[6]));
  AL_FADD comp21_60 (
    .a(1'b0),
    .b(sum_20[60]),
    .c(cout_21[59]),
    .cout(cout_21[60]),
    .sum(sum_21[60]));
  AL_FADD comp21_61 (
    .a(1'b0),
    .b(sum_20[61]),
    .c(cout_21[60]),
    .cout(cout_21[61]),
    .sum(sum_21[61]));
  AL_FADD comp21_62 (
    .a(1'b0),
    .b(sum_20[62]),
    .c(cout_21[61]),
    .cout(cout_21[62]),
    .sum(sum_21[62]));
  AL_FADD comp21_63 (
    .a(1'b0),
    .b(sum_20[63]),
    .c(cout_21[62]),
    .cout(cout_21[63]),
    .sum(sum_21[63]));
  AL_FADD comp21_7 (
    .a(i21[7]),
    .b(sum_20[7]),
    .c(cout_21[6]),
    .cout(cout_21[7]),
    .sum(sum_21[7]));
  AL_FADD comp21_8 (
    .a(i21[8]),
    .b(sum_20[8]),
    .c(cout_21[7]),
    .cout(cout_21[8]),
    .sum(sum_21[8]));
  AL_FADD comp21_9 (
    .a(i21[9]),
    .b(sum_20[9]),
    .c(cout_21[8]),
    .cout(cout_21[9]),
    .sum(sum_21[9]));
  AL_FADD comp22_0 (
    .a(i22[0]),
    .b(sum_21[0]),
    .c(1'b0),
    .cout(cout_22[0]),
    .sum(sum_22[0]));
  AL_FADD comp22_1 (
    .a(i22[1]),
    .b(sum_21[1]),
    .c(cout_22[0]),
    .cout(cout_22[1]),
    .sum(sum_22[1]));
  AL_FADD comp22_10 (
    .a(i22[10]),
    .b(sum_21[10]),
    .c(cout_22[9]),
    .cout(cout_22[10]),
    .sum(sum_22[10]));
  AL_FADD comp22_11 (
    .a(i22[11]),
    .b(sum_21[11]),
    .c(cout_22[10]),
    .cout(cout_22[11]),
    .sum(sum_22[11]));
  AL_FADD comp22_12 (
    .a(i22[12]),
    .b(sum_21[12]),
    .c(cout_22[11]),
    .cout(cout_22[12]),
    .sum(sum_22[12]));
  AL_FADD comp22_13 (
    .a(i22[13]),
    .b(sum_21[13]),
    .c(cout_22[12]),
    .cout(cout_22[13]),
    .sum(sum_22[13]));
  AL_FADD comp22_14 (
    .a(i22[14]),
    .b(sum_21[14]),
    .c(cout_22[13]),
    .cout(cout_22[14]),
    .sum(sum_22[14]));
  AL_FADD comp22_15 (
    .a(i22[15]),
    .b(sum_21[15]),
    .c(cout_22[14]),
    .cout(cout_22[15]),
    .sum(sum_22[15]));
  AL_FADD comp22_16 (
    .a(i22[16]),
    .b(sum_21[16]),
    .c(cout_22[15]),
    .cout(cout_22[16]),
    .sum(sum_22[16]));
  AL_FADD comp22_17 (
    .a(i22[17]),
    .b(sum_21[17]),
    .c(cout_22[16]),
    .cout(cout_22[17]),
    .sum(sum_22[17]));
  AL_FADD comp22_18 (
    .a(i22[18]),
    .b(sum_21[18]),
    .c(cout_22[17]),
    .cout(cout_22[18]),
    .sum(sum_22[18]));
  AL_FADD comp22_19 (
    .a(i22[19]),
    .b(sum_21[19]),
    .c(cout_22[18]),
    .cout(cout_22[19]),
    .sum(sum_22[19]));
  AL_FADD comp22_2 (
    .a(i22[2]),
    .b(sum_21[2]),
    .c(cout_22[1]),
    .cout(cout_22[2]),
    .sum(sum_22[2]));
  AL_FADD comp22_20 (
    .a(i22[20]),
    .b(sum_21[20]),
    .c(cout_22[19]),
    .cout(cout_22[20]),
    .sum(sum_22[20]));
  AL_FADD comp22_21 (
    .a(i22[21]),
    .b(sum_21[21]),
    .c(cout_22[20]),
    .cout(cout_22[21]),
    .sum(sum_22[21]));
  AL_FADD comp22_22 (
    .a(i22[22]),
    .b(sum_21[22]),
    .c(cout_22[21]),
    .cout(cout_22[22]),
    .sum(sum_22[22]));
  AL_FADD comp22_23 (
    .a(i22[23]),
    .b(sum_21[23]),
    .c(cout_22[22]),
    .cout(cout_22[23]),
    .sum(sum_22[23]));
  AL_FADD comp22_24 (
    .a(i22[24]),
    .b(sum_21[24]),
    .c(cout_22[23]),
    .cout(cout_22[24]),
    .sum(sum_22[24]));
  AL_FADD comp22_25 (
    .a(i22[25]),
    .b(sum_21[25]),
    .c(cout_22[24]),
    .cout(cout_22[25]),
    .sum(sum_22[25]));
  AL_FADD comp22_26 (
    .a(i22[26]),
    .b(sum_21[26]),
    .c(cout_22[25]),
    .cout(cout_22[26]),
    .sum(sum_22[26]));
  AL_FADD comp22_27 (
    .a(i22[27]),
    .b(sum_21[27]),
    .c(cout_22[26]),
    .cout(cout_22[27]),
    .sum(sum_22[27]));
  AL_FADD comp22_28 (
    .a(i22[28]),
    .b(sum_21[28]),
    .c(cout_22[27]),
    .cout(cout_22[28]),
    .sum(sum_22[28]));
  AL_FADD comp22_29 (
    .a(i22[29]),
    .b(sum_21[29]),
    .c(cout_22[28]),
    .cout(cout_22[29]),
    .sum(sum_22[29]));
  AL_FADD comp22_3 (
    .a(i22[3]),
    .b(sum_21[3]),
    .c(cout_22[2]),
    .cout(cout_22[3]),
    .sum(sum_22[3]));
  AL_FADD comp22_30 (
    .a(i22[30]),
    .b(sum_21[30]),
    .c(cout_22[29]),
    .cout(cout_22[30]),
    .sum(sum_22[30]));
  AL_FADD comp22_31 (
    .a(i22[31]),
    .b(sum_21[31]),
    .c(cout_22[30]),
    .cout(cout_22[31]),
    .sum(sum_22[31]));
  AL_FADD comp22_32 (
    .a(i22[32]),
    .b(sum_21[32]),
    .c(cout_22[31]),
    .cout(cout_22[32]),
    .sum(sum_22[32]));
  AL_FADD comp22_33 (
    .a(i22[33]),
    .b(sum_21[33]),
    .c(cout_22[32]),
    .cout(cout_22[33]),
    .sum(sum_22[33]));
  AL_FADD comp22_34 (
    .a(i22[34]),
    .b(sum_21[34]),
    .c(cout_22[33]),
    .cout(cout_22[34]),
    .sum(sum_22[34]));
  AL_FADD comp22_35 (
    .a(i22[35]),
    .b(sum_21[35]),
    .c(cout_22[34]),
    .cout(cout_22[35]),
    .sum(sum_22[35]));
  AL_FADD comp22_36 (
    .a(i22[36]),
    .b(sum_21[36]),
    .c(cout_22[35]),
    .cout(cout_22[36]),
    .sum(sum_22[36]));
  AL_FADD comp22_37 (
    .a(i22[37]),
    .b(sum_21[37]),
    .c(cout_22[36]),
    .cout(cout_22[37]),
    .sum(sum_22[37]));
  AL_FADD comp22_38 (
    .a(i22[38]),
    .b(sum_21[38]),
    .c(cout_22[37]),
    .cout(cout_22[38]),
    .sum(sum_22[38]));
  AL_FADD comp22_39 (
    .a(i22[39]),
    .b(sum_21[39]),
    .c(cout_22[38]),
    .cout(cout_22[39]),
    .sum(sum_22[39]));
  AL_FADD comp22_4 (
    .a(i22[4]),
    .b(sum_21[4]),
    .c(cout_22[3]),
    .cout(cout_22[4]),
    .sum(sum_22[4]));
  AL_FADD comp22_40 (
    .a(i22[40]),
    .b(sum_21[40]),
    .c(cout_22[39]),
    .cout(cout_22[40]),
    .sum(sum_22[40]));
  AL_FADD comp22_41 (
    .a(1'b0),
    .b(sum_21[41]),
    .c(cout_22[40]),
    .cout(cout_22[41]),
    .sum(sum_22[41]));
  AL_FADD comp22_42 (
    .a(1'b0),
    .b(sum_21[42]),
    .c(cout_22[41]),
    .cout(cout_22[42]),
    .sum(sum_22[42]));
  AL_FADD comp22_43 (
    .a(1'b0),
    .b(sum_21[43]),
    .c(cout_22[42]),
    .cout(cout_22[43]),
    .sum(sum_22[43]));
  AL_FADD comp22_44 (
    .a(1'b0),
    .b(sum_21[44]),
    .c(cout_22[43]),
    .cout(cout_22[44]),
    .sum(sum_22[44]));
  AL_FADD comp22_45 (
    .a(1'b0),
    .b(sum_21[45]),
    .c(cout_22[44]),
    .cout(cout_22[45]),
    .sum(sum_22[45]));
  AL_FADD comp22_46 (
    .a(1'b0),
    .b(sum_21[46]),
    .c(cout_22[45]),
    .cout(cout_22[46]),
    .sum(sum_22[46]));
  AL_FADD comp22_47 (
    .a(1'b0),
    .b(sum_21[47]),
    .c(cout_22[46]),
    .cout(cout_22[47]),
    .sum(sum_22[47]));
  AL_FADD comp22_48 (
    .a(1'b0),
    .b(sum_21[48]),
    .c(cout_22[47]),
    .cout(cout_22[48]),
    .sum(sum_22[48]));
  AL_FADD comp22_49 (
    .a(1'b0),
    .b(sum_21[49]),
    .c(cout_22[48]),
    .cout(cout_22[49]),
    .sum(sum_22[49]));
  AL_FADD comp22_5 (
    .a(i22[5]),
    .b(sum_21[5]),
    .c(cout_22[4]),
    .cout(cout_22[5]),
    .sum(sum_22[5]));
  AL_FADD comp22_50 (
    .a(1'b0),
    .b(sum_21[50]),
    .c(cout_22[49]),
    .cout(cout_22[50]),
    .sum(sum_22[50]));
  AL_FADD comp22_51 (
    .a(1'b0),
    .b(sum_21[51]),
    .c(cout_22[50]),
    .cout(cout_22[51]),
    .sum(sum_22[51]));
  AL_FADD comp22_52 (
    .a(1'b0),
    .b(sum_21[52]),
    .c(cout_22[51]),
    .cout(cout_22[52]),
    .sum(sum_22[52]));
  AL_FADD comp22_53 (
    .a(1'b0),
    .b(sum_21[53]),
    .c(cout_22[52]),
    .cout(cout_22[53]),
    .sum(sum_22[53]));
  AL_FADD comp22_54 (
    .a(1'b0),
    .b(sum_21[54]),
    .c(cout_22[53]),
    .cout(cout_22[54]),
    .sum(sum_22[54]));
  AL_FADD comp22_55 (
    .a(1'b0),
    .b(sum_21[55]),
    .c(cout_22[54]),
    .cout(cout_22[55]),
    .sum(sum_22[55]));
  AL_FADD comp22_56 (
    .a(1'b0),
    .b(sum_21[56]),
    .c(cout_22[55]),
    .cout(cout_22[56]),
    .sum(sum_22[56]));
  AL_FADD comp22_57 (
    .a(1'b0),
    .b(sum_21[57]),
    .c(cout_22[56]),
    .cout(cout_22[57]),
    .sum(sum_22[57]));
  AL_FADD comp22_58 (
    .a(1'b0),
    .b(sum_21[58]),
    .c(cout_22[57]),
    .cout(cout_22[58]),
    .sum(sum_22[58]));
  AL_FADD comp22_59 (
    .a(1'b0),
    .b(sum_21[59]),
    .c(cout_22[58]),
    .cout(cout_22[59]),
    .sum(sum_22[59]));
  AL_FADD comp22_6 (
    .a(i22[6]),
    .b(sum_21[6]),
    .c(cout_22[5]),
    .cout(cout_22[6]),
    .sum(sum_22[6]));
  AL_FADD comp22_60 (
    .a(1'b0),
    .b(sum_21[60]),
    .c(cout_22[59]),
    .cout(cout_22[60]),
    .sum(sum_22[60]));
  AL_FADD comp22_61 (
    .a(1'b0),
    .b(sum_21[61]),
    .c(cout_22[60]),
    .cout(cout_22[61]),
    .sum(sum_22[61]));
  AL_FADD comp22_62 (
    .a(1'b0),
    .b(sum_21[62]),
    .c(cout_22[61]),
    .cout(cout_22[62]),
    .sum(sum_22[62]));
  AL_FADD comp22_63 (
    .a(1'b0),
    .b(sum_21[63]),
    .c(cout_22[62]),
    .cout(cout_22[63]),
    .sum(sum_22[63]));
  AL_FADD comp22_7 (
    .a(i22[7]),
    .b(sum_21[7]),
    .c(cout_22[6]),
    .cout(cout_22[7]),
    .sum(sum_22[7]));
  AL_FADD comp22_8 (
    .a(i22[8]),
    .b(sum_21[8]),
    .c(cout_22[7]),
    .cout(cout_22[8]),
    .sum(sum_22[8]));
  AL_FADD comp22_9 (
    .a(i22[9]),
    .b(sum_21[9]),
    .c(cout_22[8]),
    .cout(cout_22[9]),
    .sum(sum_22[9]));
  AL_FADD comp23_0 (
    .a(i23[0]),
    .b(sum_22[0]),
    .c(1'b0),
    .cout(cout_23[0]),
    .sum(sum_23[0]));
  AL_FADD comp23_1 (
    .a(i23[1]),
    .b(sum_22[1]),
    .c(cout_23[0]),
    .cout(cout_23[1]),
    .sum(sum_23[1]));
  AL_FADD comp23_10 (
    .a(i23[10]),
    .b(sum_22[10]),
    .c(cout_23[9]),
    .cout(cout_23[10]),
    .sum(sum_23[10]));
  AL_FADD comp23_11 (
    .a(i23[11]),
    .b(sum_22[11]),
    .c(cout_23[10]),
    .cout(cout_23[11]),
    .sum(sum_23[11]));
  AL_FADD comp23_12 (
    .a(i23[12]),
    .b(sum_22[12]),
    .c(cout_23[11]),
    .cout(cout_23[12]),
    .sum(sum_23[12]));
  AL_FADD comp23_13 (
    .a(i23[13]),
    .b(sum_22[13]),
    .c(cout_23[12]),
    .cout(cout_23[13]),
    .sum(sum_23[13]));
  AL_FADD comp23_14 (
    .a(i23[14]),
    .b(sum_22[14]),
    .c(cout_23[13]),
    .cout(cout_23[14]),
    .sum(sum_23[14]));
  AL_FADD comp23_15 (
    .a(i23[15]),
    .b(sum_22[15]),
    .c(cout_23[14]),
    .cout(cout_23[15]),
    .sum(sum_23[15]));
  AL_FADD comp23_16 (
    .a(i23[16]),
    .b(sum_22[16]),
    .c(cout_23[15]),
    .cout(cout_23[16]),
    .sum(sum_23[16]));
  AL_FADD comp23_17 (
    .a(i23[17]),
    .b(sum_22[17]),
    .c(cout_23[16]),
    .cout(cout_23[17]),
    .sum(sum_23[17]));
  AL_FADD comp23_18 (
    .a(i23[18]),
    .b(sum_22[18]),
    .c(cout_23[17]),
    .cout(cout_23[18]),
    .sum(sum_23[18]));
  AL_FADD comp23_19 (
    .a(i23[19]),
    .b(sum_22[19]),
    .c(cout_23[18]),
    .cout(cout_23[19]),
    .sum(sum_23[19]));
  AL_FADD comp23_2 (
    .a(i23[2]),
    .b(sum_22[2]),
    .c(cout_23[1]),
    .cout(cout_23[2]),
    .sum(sum_23[2]));
  AL_FADD comp23_20 (
    .a(i23[20]),
    .b(sum_22[20]),
    .c(cout_23[19]),
    .cout(cout_23[20]),
    .sum(sum_23[20]));
  AL_FADD comp23_21 (
    .a(i23[21]),
    .b(sum_22[21]),
    .c(cout_23[20]),
    .cout(cout_23[21]),
    .sum(sum_23[21]));
  AL_FADD comp23_22 (
    .a(i23[22]),
    .b(sum_22[22]),
    .c(cout_23[21]),
    .cout(cout_23[22]),
    .sum(sum_23[22]));
  AL_FADD comp23_23 (
    .a(i23[23]),
    .b(sum_22[23]),
    .c(cout_23[22]),
    .cout(cout_23[23]),
    .sum(sum_23[23]));
  AL_FADD comp23_24 (
    .a(i23[24]),
    .b(sum_22[24]),
    .c(cout_23[23]),
    .cout(cout_23[24]),
    .sum(sum_23[24]));
  AL_FADD comp23_25 (
    .a(i23[25]),
    .b(sum_22[25]),
    .c(cout_23[24]),
    .cout(cout_23[25]),
    .sum(sum_23[25]));
  AL_FADD comp23_26 (
    .a(i23[26]),
    .b(sum_22[26]),
    .c(cout_23[25]),
    .cout(cout_23[26]),
    .sum(sum_23[26]));
  AL_FADD comp23_27 (
    .a(i23[27]),
    .b(sum_22[27]),
    .c(cout_23[26]),
    .cout(cout_23[27]),
    .sum(sum_23[27]));
  AL_FADD comp23_28 (
    .a(i23[28]),
    .b(sum_22[28]),
    .c(cout_23[27]),
    .cout(cout_23[28]),
    .sum(sum_23[28]));
  AL_FADD comp23_29 (
    .a(i23[29]),
    .b(sum_22[29]),
    .c(cout_23[28]),
    .cout(cout_23[29]),
    .sum(sum_23[29]));
  AL_FADD comp23_3 (
    .a(i23[3]),
    .b(sum_22[3]),
    .c(cout_23[2]),
    .cout(cout_23[3]),
    .sum(sum_23[3]));
  AL_FADD comp23_30 (
    .a(i23[30]),
    .b(sum_22[30]),
    .c(cout_23[29]),
    .cout(cout_23[30]),
    .sum(sum_23[30]));
  AL_FADD comp23_31 (
    .a(i23[31]),
    .b(sum_22[31]),
    .c(cout_23[30]),
    .cout(cout_23[31]),
    .sum(sum_23[31]));
  AL_FADD comp23_32 (
    .a(i23[32]),
    .b(sum_22[32]),
    .c(cout_23[31]),
    .cout(cout_23[32]),
    .sum(sum_23[32]));
  AL_FADD comp23_33 (
    .a(i23[33]),
    .b(sum_22[33]),
    .c(cout_23[32]),
    .cout(cout_23[33]),
    .sum(sum_23[33]));
  AL_FADD comp23_34 (
    .a(i23[34]),
    .b(sum_22[34]),
    .c(cout_23[33]),
    .cout(cout_23[34]),
    .sum(sum_23[34]));
  AL_FADD comp23_35 (
    .a(i23[35]),
    .b(sum_22[35]),
    .c(cout_23[34]),
    .cout(cout_23[35]),
    .sum(sum_23[35]));
  AL_FADD comp23_36 (
    .a(i23[36]),
    .b(sum_22[36]),
    .c(cout_23[35]),
    .cout(cout_23[36]),
    .sum(sum_23[36]));
  AL_FADD comp23_37 (
    .a(i23[37]),
    .b(sum_22[37]),
    .c(cout_23[36]),
    .cout(cout_23[37]),
    .sum(sum_23[37]));
  AL_FADD comp23_38 (
    .a(i23[38]),
    .b(sum_22[38]),
    .c(cout_23[37]),
    .cout(cout_23[38]),
    .sum(sum_23[38]));
  AL_FADD comp23_39 (
    .a(i23[39]),
    .b(sum_22[39]),
    .c(cout_23[38]),
    .cout(cout_23[39]),
    .sum(sum_23[39]));
  AL_FADD comp23_4 (
    .a(i23[4]),
    .b(sum_22[4]),
    .c(cout_23[3]),
    .cout(cout_23[4]),
    .sum(sum_23[4]));
  AL_FADD comp23_40 (
    .a(1'b0),
    .b(sum_22[40]),
    .c(cout_23[39]),
    .cout(cout_23[40]),
    .sum(sum_23[40]));
  AL_FADD comp23_41 (
    .a(1'b0),
    .b(sum_22[41]),
    .c(cout_23[40]),
    .cout(cout_23[41]),
    .sum(sum_23[41]));
  AL_FADD comp23_42 (
    .a(1'b0),
    .b(sum_22[42]),
    .c(cout_23[41]),
    .cout(cout_23[42]),
    .sum(sum_23[42]));
  AL_FADD comp23_43 (
    .a(1'b0),
    .b(sum_22[43]),
    .c(cout_23[42]),
    .cout(cout_23[43]),
    .sum(sum_23[43]));
  AL_FADD comp23_44 (
    .a(1'b0),
    .b(sum_22[44]),
    .c(cout_23[43]),
    .cout(cout_23[44]),
    .sum(sum_23[44]));
  AL_FADD comp23_45 (
    .a(1'b0),
    .b(sum_22[45]),
    .c(cout_23[44]),
    .cout(cout_23[45]),
    .sum(sum_23[45]));
  AL_FADD comp23_46 (
    .a(1'b0),
    .b(sum_22[46]),
    .c(cout_23[45]),
    .cout(cout_23[46]),
    .sum(sum_23[46]));
  AL_FADD comp23_47 (
    .a(1'b0),
    .b(sum_22[47]),
    .c(cout_23[46]),
    .cout(cout_23[47]),
    .sum(sum_23[47]));
  AL_FADD comp23_48 (
    .a(1'b0),
    .b(sum_22[48]),
    .c(cout_23[47]),
    .cout(cout_23[48]),
    .sum(sum_23[48]));
  AL_FADD comp23_49 (
    .a(1'b0),
    .b(sum_22[49]),
    .c(cout_23[48]),
    .cout(cout_23[49]),
    .sum(sum_23[49]));
  AL_FADD comp23_5 (
    .a(i23[5]),
    .b(sum_22[5]),
    .c(cout_23[4]),
    .cout(cout_23[5]),
    .sum(sum_23[5]));
  AL_FADD comp23_50 (
    .a(1'b0),
    .b(sum_22[50]),
    .c(cout_23[49]),
    .cout(cout_23[50]),
    .sum(sum_23[50]));
  AL_FADD comp23_51 (
    .a(1'b0),
    .b(sum_22[51]),
    .c(cout_23[50]),
    .cout(cout_23[51]),
    .sum(sum_23[51]));
  AL_FADD comp23_52 (
    .a(1'b0),
    .b(sum_22[52]),
    .c(cout_23[51]),
    .cout(cout_23[52]),
    .sum(sum_23[52]));
  AL_FADD comp23_53 (
    .a(1'b0),
    .b(sum_22[53]),
    .c(cout_23[52]),
    .cout(cout_23[53]),
    .sum(sum_23[53]));
  AL_FADD comp23_54 (
    .a(1'b0),
    .b(sum_22[54]),
    .c(cout_23[53]),
    .cout(cout_23[54]),
    .sum(sum_23[54]));
  AL_FADD comp23_55 (
    .a(1'b0),
    .b(sum_22[55]),
    .c(cout_23[54]),
    .cout(cout_23[55]),
    .sum(sum_23[55]));
  AL_FADD comp23_56 (
    .a(1'b0),
    .b(sum_22[56]),
    .c(cout_23[55]),
    .cout(cout_23[56]),
    .sum(sum_23[56]));
  AL_FADD comp23_57 (
    .a(1'b0),
    .b(sum_22[57]),
    .c(cout_23[56]),
    .cout(cout_23[57]),
    .sum(sum_23[57]));
  AL_FADD comp23_58 (
    .a(1'b0),
    .b(sum_22[58]),
    .c(cout_23[57]),
    .cout(cout_23[58]),
    .sum(sum_23[58]));
  AL_FADD comp23_59 (
    .a(1'b0),
    .b(sum_22[59]),
    .c(cout_23[58]),
    .cout(cout_23[59]),
    .sum(sum_23[59]));
  AL_FADD comp23_6 (
    .a(i23[6]),
    .b(sum_22[6]),
    .c(cout_23[5]),
    .cout(cout_23[6]),
    .sum(sum_23[6]));
  AL_FADD comp23_60 (
    .a(1'b0),
    .b(sum_22[60]),
    .c(cout_23[59]),
    .cout(cout_23[60]),
    .sum(sum_23[60]));
  AL_FADD comp23_61 (
    .a(1'b0),
    .b(sum_22[61]),
    .c(cout_23[60]),
    .cout(cout_23[61]),
    .sum(sum_23[61]));
  AL_FADD comp23_62 (
    .a(1'b0),
    .b(sum_22[62]),
    .c(cout_23[61]),
    .cout(cout_23[62]),
    .sum(sum_23[62]));
  AL_FADD comp23_63 (
    .a(1'b0),
    .b(sum_22[63]),
    .c(cout_23[62]),
    .cout(cout_23[63]),
    .sum(sum_23[63]));
  AL_FADD comp23_7 (
    .a(i23[7]),
    .b(sum_22[7]),
    .c(cout_23[6]),
    .cout(cout_23[7]),
    .sum(sum_23[7]));
  AL_FADD comp23_8 (
    .a(i23[8]),
    .b(sum_22[8]),
    .c(cout_23[7]),
    .cout(cout_23[8]),
    .sum(sum_23[8]));
  AL_FADD comp23_9 (
    .a(i23[9]),
    .b(sum_22[9]),
    .c(cout_23[8]),
    .cout(cout_23[9]),
    .sum(sum_23[9]));
  AL_FADD comp24_0 (
    .a(i24[0]),
    .b(sum_23[0]),
    .c(1'b0),
    .cout(cout_24[0]),
    .sum(sum_24[0]));
  AL_FADD comp24_1 (
    .a(i24[1]),
    .b(sum_23[1]),
    .c(cout_24[0]),
    .cout(cout_24[1]),
    .sum(sum_24[1]));
  AL_FADD comp24_10 (
    .a(i24[10]),
    .b(sum_23[10]),
    .c(cout_24[9]),
    .cout(cout_24[10]),
    .sum(sum_24[10]));
  AL_FADD comp24_11 (
    .a(i24[11]),
    .b(sum_23[11]),
    .c(cout_24[10]),
    .cout(cout_24[11]),
    .sum(sum_24[11]));
  AL_FADD comp24_12 (
    .a(i24[12]),
    .b(sum_23[12]),
    .c(cout_24[11]),
    .cout(cout_24[12]),
    .sum(sum_24[12]));
  AL_FADD comp24_13 (
    .a(i24[13]),
    .b(sum_23[13]),
    .c(cout_24[12]),
    .cout(cout_24[13]),
    .sum(sum_24[13]));
  AL_FADD comp24_14 (
    .a(i24[14]),
    .b(sum_23[14]),
    .c(cout_24[13]),
    .cout(cout_24[14]),
    .sum(sum_24[14]));
  AL_FADD comp24_15 (
    .a(i24[15]),
    .b(sum_23[15]),
    .c(cout_24[14]),
    .cout(cout_24[15]),
    .sum(sum_24[15]));
  AL_FADD comp24_16 (
    .a(i24[16]),
    .b(sum_23[16]),
    .c(cout_24[15]),
    .cout(cout_24[16]),
    .sum(sum_24[16]));
  AL_FADD comp24_17 (
    .a(i24[17]),
    .b(sum_23[17]),
    .c(cout_24[16]),
    .cout(cout_24[17]),
    .sum(sum_24[17]));
  AL_FADD comp24_18 (
    .a(i24[18]),
    .b(sum_23[18]),
    .c(cout_24[17]),
    .cout(cout_24[18]),
    .sum(sum_24[18]));
  AL_FADD comp24_19 (
    .a(i24[19]),
    .b(sum_23[19]),
    .c(cout_24[18]),
    .cout(cout_24[19]),
    .sum(sum_24[19]));
  AL_FADD comp24_2 (
    .a(i24[2]),
    .b(sum_23[2]),
    .c(cout_24[1]),
    .cout(cout_24[2]),
    .sum(sum_24[2]));
  AL_FADD comp24_20 (
    .a(i24[20]),
    .b(sum_23[20]),
    .c(cout_24[19]),
    .cout(cout_24[20]),
    .sum(sum_24[20]));
  AL_FADD comp24_21 (
    .a(i24[21]),
    .b(sum_23[21]),
    .c(cout_24[20]),
    .cout(cout_24[21]),
    .sum(sum_24[21]));
  AL_FADD comp24_22 (
    .a(i24[22]),
    .b(sum_23[22]),
    .c(cout_24[21]),
    .cout(cout_24[22]),
    .sum(sum_24[22]));
  AL_FADD comp24_23 (
    .a(i24[23]),
    .b(sum_23[23]),
    .c(cout_24[22]),
    .cout(cout_24[23]),
    .sum(sum_24[23]));
  AL_FADD comp24_24 (
    .a(i24[24]),
    .b(sum_23[24]),
    .c(cout_24[23]),
    .cout(cout_24[24]),
    .sum(sum_24[24]));
  AL_FADD comp24_25 (
    .a(i24[25]),
    .b(sum_23[25]),
    .c(cout_24[24]),
    .cout(cout_24[25]),
    .sum(sum_24[25]));
  AL_FADD comp24_26 (
    .a(i24[26]),
    .b(sum_23[26]),
    .c(cout_24[25]),
    .cout(cout_24[26]),
    .sum(sum_24[26]));
  AL_FADD comp24_27 (
    .a(i24[27]),
    .b(sum_23[27]),
    .c(cout_24[26]),
    .cout(cout_24[27]),
    .sum(sum_24[27]));
  AL_FADD comp24_28 (
    .a(i24[28]),
    .b(sum_23[28]),
    .c(cout_24[27]),
    .cout(cout_24[28]),
    .sum(sum_24[28]));
  AL_FADD comp24_29 (
    .a(i24[29]),
    .b(sum_23[29]),
    .c(cout_24[28]),
    .cout(cout_24[29]),
    .sum(sum_24[29]));
  AL_FADD comp24_3 (
    .a(i24[3]),
    .b(sum_23[3]),
    .c(cout_24[2]),
    .cout(cout_24[3]),
    .sum(sum_24[3]));
  AL_FADD comp24_30 (
    .a(i24[30]),
    .b(sum_23[30]),
    .c(cout_24[29]),
    .cout(cout_24[30]),
    .sum(sum_24[30]));
  AL_FADD comp24_31 (
    .a(i24[31]),
    .b(sum_23[31]),
    .c(cout_24[30]),
    .cout(cout_24[31]),
    .sum(sum_24[31]));
  AL_FADD comp24_32 (
    .a(i24[32]),
    .b(sum_23[32]),
    .c(cout_24[31]),
    .cout(cout_24[32]),
    .sum(sum_24[32]));
  AL_FADD comp24_33 (
    .a(i24[33]),
    .b(sum_23[33]),
    .c(cout_24[32]),
    .cout(cout_24[33]),
    .sum(sum_24[33]));
  AL_FADD comp24_34 (
    .a(i24[34]),
    .b(sum_23[34]),
    .c(cout_24[33]),
    .cout(cout_24[34]),
    .sum(sum_24[34]));
  AL_FADD comp24_35 (
    .a(i24[35]),
    .b(sum_23[35]),
    .c(cout_24[34]),
    .cout(cout_24[35]),
    .sum(sum_24[35]));
  AL_FADD comp24_36 (
    .a(i24[36]),
    .b(sum_23[36]),
    .c(cout_24[35]),
    .cout(cout_24[36]),
    .sum(sum_24[36]));
  AL_FADD comp24_37 (
    .a(i24[37]),
    .b(sum_23[37]),
    .c(cout_24[36]),
    .cout(cout_24[37]),
    .sum(sum_24[37]));
  AL_FADD comp24_38 (
    .a(i24[38]),
    .b(sum_23[38]),
    .c(cout_24[37]),
    .cout(cout_24[38]),
    .sum(sum_24[38]));
  AL_FADD comp24_39 (
    .a(1'b0),
    .b(sum_23[39]),
    .c(cout_24[38]),
    .cout(cout_24[39]),
    .sum(sum_24[39]));
  AL_FADD comp24_4 (
    .a(i24[4]),
    .b(sum_23[4]),
    .c(cout_24[3]),
    .cout(cout_24[4]),
    .sum(sum_24[4]));
  AL_FADD comp24_40 (
    .a(1'b0),
    .b(sum_23[40]),
    .c(cout_24[39]),
    .cout(cout_24[40]),
    .sum(sum_24[40]));
  AL_FADD comp24_41 (
    .a(1'b0),
    .b(sum_23[41]),
    .c(cout_24[40]),
    .cout(cout_24[41]),
    .sum(sum_24[41]));
  AL_FADD comp24_42 (
    .a(1'b0),
    .b(sum_23[42]),
    .c(cout_24[41]),
    .cout(cout_24[42]),
    .sum(sum_24[42]));
  AL_FADD comp24_43 (
    .a(1'b0),
    .b(sum_23[43]),
    .c(cout_24[42]),
    .cout(cout_24[43]),
    .sum(sum_24[43]));
  AL_FADD comp24_44 (
    .a(1'b0),
    .b(sum_23[44]),
    .c(cout_24[43]),
    .cout(cout_24[44]),
    .sum(sum_24[44]));
  AL_FADD comp24_45 (
    .a(1'b0),
    .b(sum_23[45]),
    .c(cout_24[44]),
    .cout(cout_24[45]),
    .sum(sum_24[45]));
  AL_FADD comp24_46 (
    .a(1'b0),
    .b(sum_23[46]),
    .c(cout_24[45]),
    .cout(cout_24[46]),
    .sum(sum_24[46]));
  AL_FADD comp24_47 (
    .a(1'b0),
    .b(sum_23[47]),
    .c(cout_24[46]),
    .cout(cout_24[47]),
    .sum(sum_24[47]));
  AL_FADD comp24_48 (
    .a(1'b0),
    .b(sum_23[48]),
    .c(cout_24[47]),
    .cout(cout_24[48]),
    .sum(sum_24[48]));
  AL_FADD comp24_49 (
    .a(1'b0),
    .b(sum_23[49]),
    .c(cout_24[48]),
    .cout(cout_24[49]),
    .sum(sum_24[49]));
  AL_FADD comp24_5 (
    .a(i24[5]),
    .b(sum_23[5]),
    .c(cout_24[4]),
    .cout(cout_24[5]),
    .sum(sum_24[5]));
  AL_FADD comp24_50 (
    .a(1'b0),
    .b(sum_23[50]),
    .c(cout_24[49]),
    .cout(cout_24[50]),
    .sum(sum_24[50]));
  AL_FADD comp24_51 (
    .a(1'b0),
    .b(sum_23[51]),
    .c(cout_24[50]),
    .cout(cout_24[51]),
    .sum(sum_24[51]));
  AL_FADD comp24_52 (
    .a(1'b0),
    .b(sum_23[52]),
    .c(cout_24[51]),
    .cout(cout_24[52]),
    .sum(sum_24[52]));
  AL_FADD comp24_53 (
    .a(1'b0),
    .b(sum_23[53]),
    .c(cout_24[52]),
    .cout(cout_24[53]),
    .sum(sum_24[53]));
  AL_FADD comp24_54 (
    .a(1'b0),
    .b(sum_23[54]),
    .c(cout_24[53]),
    .cout(cout_24[54]),
    .sum(sum_24[54]));
  AL_FADD comp24_55 (
    .a(1'b0),
    .b(sum_23[55]),
    .c(cout_24[54]),
    .cout(cout_24[55]),
    .sum(sum_24[55]));
  AL_FADD comp24_56 (
    .a(1'b0),
    .b(sum_23[56]),
    .c(cout_24[55]),
    .cout(cout_24[56]),
    .sum(sum_24[56]));
  AL_FADD comp24_57 (
    .a(1'b0),
    .b(sum_23[57]),
    .c(cout_24[56]),
    .cout(cout_24[57]),
    .sum(sum_24[57]));
  AL_FADD comp24_58 (
    .a(1'b0),
    .b(sum_23[58]),
    .c(cout_24[57]),
    .cout(cout_24[58]),
    .sum(sum_24[58]));
  AL_FADD comp24_59 (
    .a(1'b0),
    .b(sum_23[59]),
    .c(cout_24[58]),
    .cout(cout_24[59]),
    .sum(sum_24[59]));
  AL_FADD comp24_6 (
    .a(i24[6]),
    .b(sum_23[6]),
    .c(cout_24[5]),
    .cout(cout_24[6]),
    .sum(sum_24[6]));
  AL_FADD comp24_60 (
    .a(1'b0),
    .b(sum_23[60]),
    .c(cout_24[59]),
    .cout(cout_24[60]),
    .sum(sum_24[60]));
  AL_FADD comp24_61 (
    .a(1'b0),
    .b(sum_23[61]),
    .c(cout_24[60]),
    .cout(cout_24[61]),
    .sum(sum_24[61]));
  AL_FADD comp24_62 (
    .a(1'b0),
    .b(sum_23[62]),
    .c(cout_24[61]),
    .cout(cout_24[62]),
    .sum(sum_24[62]));
  AL_FADD comp24_63 (
    .a(1'b0),
    .b(sum_23[63]),
    .c(cout_24[62]),
    .cout(cout_24[63]),
    .sum(sum_24[63]));
  AL_FADD comp24_7 (
    .a(i24[7]),
    .b(sum_23[7]),
    .c(cout_24[6]),
    .cout(cout_24[7]),
    .sum(sum_24[7]));
  AL_FADD comp24_8 (
    .a(i24[8]),
    .b(sum_23[8]),
    .c(cout_24[7]),
    .cout(cout_24[8]),
    .sum(sum_24[8]));
  AL_FADD comp24_9 (
    .a(i24[9]),
    .b(sum_23[9]),
    .c(cout_24[8]),
    .cout(cout_24[9]),
    .sum(sum_24[9]));
  AL_FADD comp25_0 (
    .a(i25[0]),
    .b(sum_24[0]),
    .c(1'b0),
    .cout(cout_25[0]),
    .sum(sum_25[0]));
  AL_FADD comp25_1 (
    .a(i25[1]),
    .b(sum_24[1]),
    .c(cout_25[0]),
    .cout(cout_25[1]),
    .sum(sum_25[1]));
  AL_FADD comp25_10 (
    .a(i25[10]),
    .b(sum_24[10]),
    .c(cout_25[9]),
    .cout(cout_25[10]),
    .sum(sum_25[10]));
  AL_FADD comp25_11 (
    .a(i25[11]),
    .b(sum_24[11]),
    .c(cout_25[10]),
    .cout(cout_25[11]),
    .sum(sum_25[11]));
  AL_FADD comp25_12 (
    .a(i25[12]),
    .b(sum_24[12]),
    .c(cout_25[11]),
    .cout(cout_25[12]),
    .sum(sum_25[12]));
  AL_FADD comp25_13 (
    .a(i25[13]),
    .b(sum_24[13]),
    .c(cout_25[12]),
    .cout(cout_25[13]),
    .sum(sum_25[13]));
  AL_FADD comp25_14 (
    .a(i25[14]),
    .b(sum_24[14]),
    .c(cout_25[13]),
    .cout(cout_25[14]),
    .sum(sum_25[14]));
  AL_FADD comp25_15 (
    .a(i25[15]),
    .b(sum_24[15]),
    .c(cout_25[14]),
    .cout(cout_25[15]),
    .sum(sum_25[15]));
  AL_FADD comp25_16 (
    .a(i25[16]),
    .b(sum_24[16]),
    .c(cout_25[15]),
    .cout(cout_25[16]),
    .sum(sum_25[16]));
  AL_FADD comp25_17 (
    .a(i25[17]),
    .b(sum_24[17]),
    .c(cout_25[16]),
    .cout(cout_25[17]),
    .sum(sum_25[17]));
  AL_FADD comp25_18 (
    .a(i25[18]),
    .b(sum_24[18]),
    .c(cout_25[17]),
    .cout(cout_25[18]),
    .sum(sum_25[18]));
  AL_FADD comp25_19 (
    .a(i25[19]),
    .b(sum_24[19]),
    .c(cout_25[18]),
    .cout(cout_25[19]),
    .sum(sum_25[19]));
  AL_FADD comp25_2 (
    .a(i25[2]),
    .b(sum_24[2]),
    .c(cout_25[1]),
    .cout(cout_25[2]),
    .sum(sum_25[2]));
  AL_FADD comp25_20 (
    .a(i25[20]),
    .b(sum_24[20]),
    .c(cout_25[19]),
    .cout(cout_25[20]),
    .sum(sum_25[20]));
  AL_FADD comp25_21 (
    .a(i25[21]),
    .b(sum_24[21]),
    .c(cout_25[20]),
    .cout(cout_25[21]),
    .sum(sum_25[21]));
  AL_FADD comp25_22 (
    .a(i25[22]),
    .b(sum_24[22]),
    .c(cout_25[21]),
    .cout(cout_25[22]),
    .sum(sum_25[22]));
  AL_FADD comp25_23 (
    .a(i25[23]),
    .b(sum_24[23]),
    .c(cout_25[22]),
    .cout(cout_25[23]),
    .sum(sum_25[23]));
  AL_FADD comp25_24 (
    .a(i25[24]),
    .b(sum_24[24]),
    .c(cout_25[23]),
    .cout(cout_25[24]),
    .sum(sum_25[24]));
  AL_FADD comp25_25 (
    .a(i25[25]),
    .b(sum_24[25]),
    .c(cout_25[24]),
    .cout(cout_25[25]),
    .sum(sum_25[25]));
  AL_FADD comp25_26 (
    .a(i25[26]),
    .b(sum_24[26]),
    .c(cout_25[25]),
    .cout(cout_25[26]),
    .sum(sum_25[26]));
  AL_FADD comp25_27 (
    .a(i25[27]),
    .b(sum_24[27]),
    .c(cout_25[26]),
    .cout(cout_25[27]),
    .sum(sum_25[27]));
  AL_FADD comp25_28 (
    .a(i25[28]),
    .b(sum_24[28]),
    .c(cout_25[27]),
    .cout(cout_25[28]),
    .sum(sum_25[28]));
  AL_FADD comp25_29 (
    .a(i25[29]),
    .b(sum_24[29]),
    .c(cout_25[28]),
    .cout(cout_25[29]),
    .sum(sum_25[29]));
  AL_FADD comp25_3 (
    .a(i25[3]),
    .b(sum_24[3]),
    .c(cout_25[2]),
    .cout(cout_25[3]),
    .sum(sum_25[3]));
  AL_FADD comp25_30 (
    .a(i25[30]),
    .b(sum_24[30]),
    .c(cout_25[29]),
    .cout(cout_25[30]),
    .sum(sum_25[30]));
  AL_FADD comp25_31 (
    .a(i25[31]),
    .b(sum_24[31]),
    .c(cout_25[30]),
    .cout(cout_25[31]),
    .sum(sum_25[31]));
  AL_FADD comp25_32 (
    .a(i25[32]),
    .b(sum_24[32]),
    .c(cout_25[31]),
    .cout(cout_25[32]),
    .sum(sum_25[32]));
  AL_FADD comp25_33 (
    .a(i25[33]),
    .b(sum_24[33]),
    .c(cout_25[32]),
    .cout(cout_25[33]),
    .sum(sum_25[33]));
  AL_FADD comp25_34 (
    .a(i25[34]),
    .b(sum_24[34]),
    .c(cout_25[33]),
    .cout(cout_25[34]),
    .sum(sum_25[34]));
  AL_FADD comp25_35 (
    .a(i25[35]),
    .b(sum_24[35]),
    .c(cout_25[34]),
    .cout(cout_25[35]),
    .sum(sum_25[35]));
  AL_FADD comp25_36 (
    .a(i25[36]),
    .b(sum_24[36]),
    .c(cout_25[35]),
    .cout(cout_25[36]),
    .sum(sum_25[36]));
  AL_FADD comp25_37 (
    .a(i25[37]),
    .b(sum_24[37]),
    .c(cout_25[36]),
    .cout(cout_25[37]),
    .sum(sum_25[37]));
  AL_FADD comp25_38 (
    .a(1'b0),
    .b(sum_24[38]),
    .c(cout_25[37]),
    .cout(cout_25[38]),
    .sum(sum_25[38]));
  AL_FADD comp25_39 (
    .a(1'b0),
    .b(sum_24[39]),
    .c(cout_25[38]),
    .cout(cout_25[39]),
    .sum(sum_25[39]));
  AL_FADD comp25_4 (
    .a(i25[4]),
    .b(sum_24[4]),
    .c(cout_25[3]),
    .cout(cout_25[4]),
    .sum(sum_25[4]));
  AL_FADD comp25_40 (
    .a(1'b0),
    .b(sum_24[40]),
    .c(cout_25[39]),
    .cout(cout_25[40]),
    .sum(sum_25[40]));
  AL_FADD comp25_41 (
    .a(1'b0),
    .b(sum_24[41]),
    .c(cout_25[40]),
    .cout(cout_25[41]),
    .sum(sum_25[41]));
  AL_FADD comp25_42 (
    .a(1'b0),
    .b(sum_24[42]),
    .c(cout_25[41]),
    .cout(cout_25[42]),
    .sum(sum_25[42]));
  AL_FADD comp25_43 (
    .a(1'b0),
    .b(sum_24[43]),
    .c(cout_25[42]),
    .cout(cout_25[43]),
    .sum(sum_25[43]));
  AL_FADD comp25_44 (
    .a(1'b0),
    .b(sum_24[44]),
    .c(cout_25[43]),
    .cout(cout_25[44]),
    .sum(sum_25[44]));
  AL_FADD comp25_45 (
    .a(1'b0),
    .b(sum_24[45]),
    .c(cout_25[44]),
    .cout(cout_25[45]),
    .sum(sum_25[45]));
  AL_FADD comp25_46 (
    .a(1'b0),
    .b(sum_24[46]),
    .c(cout_25[45]),
    .cout(cout_25[46]),
    .sum(sum_25[46]));
  AL_FADD comp25_47 (
    .a(1'b0),
    .b(sum_24[47]),
    .c(cout_25[46]),
    .cout(cout_25[47]),
    .sum(sum_25[47]));
  AL_FADD comp25_48 (
    .a(1'b0),
    .b(sum_24[48]),
    .c(cout_25[47]),
    .cout(cout_25[48]),
    .sum(sum_25[48]));
  AL_FADD comp25_49 (
    .a(1'b0),
    .b(sum_24[49]),
    .c(cout_25[48]),
    .cout(cout_25[49]),
    .sum(sum_25[49]));
  AL_FADD comp25_5 (
    .a(i25[5]),
    .b(sum_24[5]),
    .c(cout_25[4]),
    .cout(cout_25[5]),
    .sum(sum_25[5]));
  AL_FADD comp25_50 (
    .a(1'b0),
    .b(sum_24[50]),
    .c(cout_25[49]),
    .cout(cout_25[50]),
    .sum(sum_25[50]));
  AL_FADD comp25_51 (
    .a(1'b0),
    .b(sum_24[51]),
    .c(cout_25[50]),
    .cout(cout_25[51]),
    .sum(sum_25[51]));
  AL_FADD comp25_52 (
    .a(1'b0),
    .b(sum_24[52]),
    .c(cout_25[51]),
    .cout(cout_25[52]),
    .sum(sum_25[52]));
  AL_FADD comp25_53 (
    .a(1'b0),
    .b(sum_24[53]),
    .c(cout_25[52]),
    .cout(cout_25[53]),
    .sum(sum_25[53]));
  AL_FADD comp25_54 (
    .a(1'b0),
    .b(sum_24[54]),
    .c(cout_25[53]),
    .cout(cout_25[54]),
    .sum(sum_25[54]));
  AL_FADD comp25_55 (
    .a(1'b0),
    .b(sum_24[55]),
    .c(cout_25[54]),
    .cout(cout_25[55]),
    .sum(sum_25[55]));
  AL_FADD comp25_56 (
    .a(1'b0),
    .b(sum_24[56]),
    .c(cout_25[55]),
    .cout(cout_25[56]),
    .sum(sum_25[56]));
  AL_FADD comp25_57 (
    .a(1'b0),
    .b(sum_24[57]),
    .c(cout_25[56]),
    .cout(cout_25[57]),
    .sum(sum_25[57]));
  AL_FADD comp25_58 (
    .a(1'b0),
    .b(sum_24[58]),
    .c(cout_25[57]),
    .cout(cout_25[58]),
    .sum(sum_25[58]));
  AL_FADD comp25_59 (
    .a(1'b0),
    .b(sum_24[59]),
    .c(cout_25[58]),
    .cout(cout_25[59]),
    .sum(sum_25[59]));
  AL_FADD comp25_6 (
    .a(i25[6]),
    .b(sum_24[6]),
    .c(cout_25[5]),
    .cout(cout_25[6]),
    .sum(sum_25[6]));
  AL_FADD comp25_60 (
    .a(1'b0),
    .b(sum_24[60]),
    .c(cout_25[59]),
    .cout(cout_25[60]),
    .sum(sum_25[60]));
  AL_FADD comp25_61 (
    .a(1'b0),
    .b(sum_24[61]),
    .c(cout_25[60]),
    .cout(cout_25[61]),
    .sum(sum_25[61]));
  AL_FADD comp25_62 (
    .a(1'b0),
    .b(sum_24[62]),
    .c(cout_25[61]),
    .cout(cout_25[62]),
    .sum(sum_25[62]));
  AL_FADD comp25_63 (
    .a(1'b0),
    .b(sum_24[63]),
    .c(cout_25[62]),
    .cout(cout_25[63]),
    .sum(sum_25[63]));
  AL_FADD comp25_7 (
    .a(i25[7]),
    .b(sum_24[7]),
    .c(cout_25[6]),
    .cout(cout_25[7]),
    .sum(sum_25[7]));
  AL_FADD comp25_8 (
    .a(i25[8]),
    .b(sum_24[8]),
    .c(cout_25[7]),
    .cout(cout_25[8]),
    .sum(sum_25[8]));
  AL_FADD comp25_9 (
    .a(i25[9]),
    .b(sum_24[9]),
    .c(cout_25[8]),
    .cout(cout_25[9]),
    .sum(sum_25[9]));
  AL_FADD comp26_0 (
    .a(i26[0]),
    .b(sum_25[0]),
    .c(1'b0),
    .cout(cout_26[0]),
    .sum(sum_26[0]));
  AL_FADD comp26_1 (
    .a(i26[1]),
    .b(sum_25[1]),
    .c(cout_26[0]),
    .cout(cout_26[1]),
    .sum(sum_26[1]));
  AL_FADD comp26_10 (
    .a(i26[10]),
    .b(sum_25[10]),
    .c(cout_26[9]),
    .cout(cout_26[10]),
    .sum(sum_26[10]));
  AL_FADD comp26_11 (
    .a(i26[11]),
    .b(sum_25[11]),
    .c(cout_26[10]),
    .cout(cout_26[11]),
    .sum(sum_26[11]));
  AL_FADD comp26_12 (
    .a(i26[12]),
    .b(sum_25[12]),
    .c(cout_26[11]),
    .cout(cout_26[12]),
    .sum(sum_26[12]));
  AL_FADD comp26_13 (
    .a(i26[13]),
    .b(sum_25[13]),
    .c(cout_26[12]),
    .cout(cout_26[13]),
    .sum(sum_26[13]));
  AL_FADD comp26_14 (
    .a(i26[14]),
    .b(sum_25[14]),
    .c(cout_26[13]),
    .cout(cout_26[14]),
    .sum(sum_26[14]));
  AL_FADD comp26_15 (
    .a(i26[15]),
    .b(sum_25[15]),
    .c(cout_26[14]),
    .cout(cout_26[15]),
    .sum(sum_26[15]));
  AL_FADD comp26_16 (
    .a(i26[16]),
    .b(sum_25[16]),
    .c(cout_26[15]),
    .cout(cout_26[16]),
    .sum(sum_26[16]));
  AL_FADD comp26_17 (
    .a(i26[17]),
    .b(sum_25[17]),
    .c(cout_26[16]),
    .cout(cout_26[17]),
    .sum(sum_26[17]));
  AL_FADD comp26_18 (
    .a(i26[18]),
    .b(sum_25[18]),
    .c(cout_26[17]),
    .cout(cout_26[18]),
    .sum(sum_26[18]));
  AL_FADD comp26_19 (
    .a(i26[19]),
    .b(sum_25[19]),
    .c(cout_26[18]),
    .cout(cout_26[19]),
    .sum(sum_26[19]));
  AL_FADD comp26_2 (
    .a(i26[2]),
    .b(sum_25[2]),
    .c(cout_26[1]),
    .cout(cout_26[2]),
    .sum(sum_26[2]));
  AL_FADD comp26_20 (
    .a(i26[20]),
    .b(sum_25[20]),
    .c(cout_26[19]),
    .cout(cout_26[20]),
    .sum(sum_26[20]));
  AL_FADD comp26_21 (
    .a(i26[21]),
    .b(sum_25[21]),
    .c(cout_26[20]),
    .cout(cout_26[21]),
    .sum(sum_26[21]));
  AL_FADD comp26_22 (
    .a(i26[22]),
    .b(sum_25[22]),
    .c(cout_26[21]),
    .cout(cout_26[22]),
    .sum(sum_26[22]));
  AL_FADD comp26_23 (
    .a(i26[23]),
    .b(sum_25[23]),
    .c(cout_26[22]),
    .cout(cout_26[23]),
    .sum(sum_26[23]));
  AL_FADD comp26_24 (
    .a(i26[24]),
    .b(sum_25[24]),
    .c(cout_26[23]),
    .cout(cout_26[24]),
    .sum(sum_26[24]));
  AL_FADD comp26_25 (
    .a(i26[25]),
    .b(sum_25[25]),
    .c(cout_26[24]),
    .cout(cout_26[25]),
    .sum(sum_26[25]));
  AL_FADD comp26_26 (
    .a(i26[26]),
    .b(sum_25[26]),
    .c(cout_26[25]),
    .cout(cout_26[26]),
    .sum(sum_26[26]));
  AL_FADD comp26_27 (
    .a(i26[27]),
    .b(sum_25[27]),
    .c(cout_26[26]),
    .cout(cout_26[27]),
    .sum(sum_26[27]));
  AL_FADD comp26_28 (
    .a(i26[28]),
    .b(sum_25[28]),
    .c(cout_26[27]),
    .cout(cout_26[28]),
    .sum(sum_26[28]));
  AL_FADD comp26_29 (
    .a(i26[29]),
    .b(sum_25[29]),
    .c(cout_26[28]),
    .cout(cout_26[29]),
    .sum(sum_26[29]));
  AL_FADD comp26_3 (
    .a(i26[3]),
    .b(sum_25[3]),
    .c(cout_26[2]),
    .cout(cout_26[3]),
    .sum(sum_26[3]));
  AL_FADD comp26_30 (
    .a(i26[30]),
    .b(sum_25[30]),
    .c(cout_26[29]),
    .cout(cout_26[30]),
    .sum(sum_26[30]));
  AL_FADD comp26_31 (
    .a(i26[31]),
    .b(sum_25[31]),
    .c(cout_26[30]),
    .cout(cout_26[31]),
    .sum(sum_26[31]));
  AL_FADD comp26_32 (
    .a(i26[32]),
    .b(sum_25[32]),
    .c(cout_26[31]),
    .cout(cout_26[32]),
    .sum(sum_26[32]));
  AL_FADD comp26_33 (
    .a(i26[33]),
    .b(sum_25[33]),
    .c(cout_26[32]),
    .cout(cout_26[33]),
    .sum(sum_26[33]));
  AL_FADD comp26_34 (
    .a(i26[34]),
    .b(sum_25[34]),
    .c(cout_26[33]),
    .cout(cout_26[34]),
    .sum(sum_26[34]));
  AL_FADD comp26_35 (
    .a(i26[35]),
    .b(sum_25[35]),
    .c(cout_26[34]),
    .cout(cout_26[35]),
    .sum(sum_26[35]));
  AL_FADD comp26_36 (
    .a(i26[36]),
    .b(sum_25[36]),
    .c(cout_26[35]),
    .cout(cout_26[36]),
    .sum(sum_26[36]));
  AL_FADD comp26_37 (
    .a(1'b0),
    .b(sum_25[37]),
    .c(cout_26[36]),
    .cout(cout_26[37]),
    .sum(sum_26[37]));
  AL_FADD comp26_38 (
    .a(1'b0),
    .b(sum_25[38]),
    .c(cout_26[37]),
    .cout(cout_26[38]),
    .sum(sum_26[38]));
  AL_FADD comp26_39 (
    .a(1'b0),
    .b(sum_25[39]),
    .c(cout_26[38]),
    .cout(cout_26[39]),
    .sum(sum_26[39]));
  AL_FADD comp26_4 (
    .a(i26[4]),
    .b(sum_25[4]),
    .c(cout_26[3]),
    .cout(cout_26[4]),
    .sum(sum_26[4]));
  AL_FADD comp26_40 (
    .a(1'b0),
    .b(sum_25[40]),
    .c(cout_26[39]),
    .cout(cout_26[40]),
    .sum(sum_26[40]));
  AL_FADD comp26_41 (
    .a(1'b0),
    .b(sum_25[41]),
    .c(cout_26[40]),
    .cout(cout_26[41]),
    .sum(sum_26[41]));
  AL_FADD comp26_42 (
    .a(1'b0),
    .b(sum_25[42]),
    .c(cout_26[41]),
    .cout(cout_26[42]),
    .sum(sum_26[42]));
  AL_FADD comp26_43 (
    .a(1'b0),
    .b(sum_25[43]),
    .c(cout_26[42]),
    .cout(cout_26[43]),
    .sum(sum_26[43]));
  AL_FADD comp26_44 (
    .a(1'b0),
    .b(sum_25[44]),
    .c(cout_26[43]),
    .cout(cout_26[44]),
    .sum(sum_26[44]));
  AL_FADD comp26_45 (
    .a(1'b0),
    .b(sum_25[45]),
    .c(cout_26[44]),
    .cout(cout_26[45]),
    .sum(sum_26[45]));
  AL_FADD comp26_46 (
    .a(1'b0),
    .b(sum_25[46]),
    .c(cout_26[45]),
    .cout(cout_26[46]),
    .sum(sum_26[46]));
  AL_FADD comp26_47 (
    .a(1'b0),
    .b(sum_25[47]),
    .c(cout_26[46]),
    .cout(cout_26[47]),
    .sum(sum_26[47]));
  AL_FADD comp26_48 (
    .a(1'b0),
    .b(sum_25[48]),
    .c(cout_26[47]),
    .cout(cout_26[48]),
    .sum(sum_26[48]));
  AL_FADD comp26_49 (
    .a(1'b0),
    .b(sum_25[49]),
    .c(cout_26[48]),
    .cout(cout_26[49]),
    .sum(sum_26[49]));
  AL_FADD comp26_5 (
    .a(i26[5]),
    .b(sum_25[5]),
    .c(cout_26[4]),
    .cout(cout_26[5]),
    .sum(sum_26[5]));
  AL_FADD comp26_50 (
    .a(1'b0),
    .b(sum_25[50]),
    .c(cout_26[49]),
    .cout(cout_26[50]),
    .sum(sum_26[50]));
  AL_FADD comp26_51 (
    .a(1'b0),
    .b(sum_25[51]),
    .c(cout_26[50]),
    .cout(cout_26[51]),
    .sum(sum_26[51]));
  AL_FADD comp26_52 (
    .a(1'b0),
    .b(sum_25[52]),
    .c(cout_26[51]),
    .cout(cout_26[52]),
    .sum(sum_26[52]));
  AL_FADD comp26_53 (
    .a(1'b0),
    .b(sum_25[53]),
    .c(cout_26[52]),
    .cout(cout_26[53]),
    .sum(sum_26[53]));
  AL_FADD comp26_54 (
    .a(1'b0),
    .b(sum_25[54]),
    .c(cout_26[53]),
    .cout(cout_26[54]),
    .sum(sum_26[54]));
  AL_FADD comp26_55 (
    .a(1'b0),
    .b(sum_25[55]),
    .c(cout_26[54]),
    .cout(cout_26[55]),
    .sum(sum_26[55]));
  AL_FADD comp26_56 (
    .a(1'b0),
    .b(sum_25[56]),
    .c(cout_26[55]),
    .cout(cout_26[56]),
    .sum(sum_26[56]));
  AL_FADD comp26_57 (
    .a(1'b0),
    .b(sum_25[57]),
    .c(cout_26[56]),
    .cout(cout_26[57]),
    .sum(sum_26[57]));
  AL_FADD comp26_58 (
    .a(1'b0),
    .b(sum_25[58]),
    .c(cout_26[57]),
    .cout(cout_26[58]),
    .sum(sum_26[58]));
  AL_FADD comp26_59 (
    .a(1'b0),
    .b(sum_25[59]),
    .c(cout_26[58]),
    .cout(cout_26[59]),
    .sum(sum_26[59]));
  AL_FADD comp26_6 (
    .a(i26[6]),
    .b(sum_25[6]),
    .c(cout_26[5]),
    .cout(cout_26[6]),
    .sum(sum_26[6]));
  AL_FADD comp26_60 (
    .a(1'b0),
    .b(sum_25[60]),
    .c(cout_26[59]),
    .cout(cout_26[60]),
    .sum(sum_26[60]));
  AL_FADD comp26_61 (
    .a(1'b0),
    .b(sum_25[61]),
    .c(cout_26[60]),
    .cout(cout_26[61]),
    .sum(sum_26[61]));
  AL_FADD comp26_62 (
    .a(1'b0),
    .b(sum_25[62]),
    .c(cout_26[61]),
    .cout(cout_26[62]),
    .sum(sum_26[62]));
  AL_FADD comp26_63 (
    .a(1'b0),
    .b(sum_25[63]),
    .c(cout_26[62]),
    .cout(cout_26[63]),
    .sum(sum_26[63]));
  AL_FADD comp26_7 (
    .a(i26[7]),
    .b(sum_25[7]),
    .c(cout_26[6]),
    .cout(cout_26[7]),
    .sum(sum_26[7]));
  AL_FADD comp26_8 (
    .a(i26[8]),
    .b(sum_25[8]),
    .c(cout_26[7]),
    .cout(cout_26[8]),
    .sum(sum_26[8]));
  AL_FADD comp26_9 (
    .a(i26[9]),
    .b(sum_25[9]),
    .c(cout_26[8]),
    .cout(cout_26[9]),
    .sum(sum_26[9]));
  AL_FADD comp27_0 (
    .a(i27[0]),
    .b(sum_26[0]),
    .c(1'b0),
    .cout(cout_27[0]),
    .sum(sum_27[0]));
  AL_FADD comp27_1 (
    .a(i27[1]),
    .b(sum_26[1]),
    .c(cout_27[0]),
    .cout(cout_27[1]),
    .sum(sum_27[1]));
  AL_FADD comp27_10 (
    .a(i27[10]),
    .b(sum_26[10]),
    .c(cout_27[9]),
    .cout(cout_27[10]),
    .sum(sum_27[10]));
  AL_FADD comp27_11 (
    .a(i27[11]),
    .b(sum_26[11]),
    .c(cout_27[10]),
    .cout(cout_27[11]),
    .sum(sum_27[11]));
  AL_FADD comp27_12 (
    .a(i27[12]),
    .b(sum_26[12]),
    .c(cout_27[11]),
    .cout(cout_27[12]),
    .sum(sum_27[12]));
  AL_FADD comp27_13 (
    .a(i27[13]),
    .b(sum_26[13]),
    .c(cout_27[12]),
    .cout(cout_27[13]),
    .sum(sum_27[13]));
  AL_FADD comp27_14 (
    .a(i27[14]),
    .b(sum_26[14]),
    .c(cout_27[13]),
    .cout(cout_27[14]),
    .sum(sum_27[14]));
  AL_FADD comp27_15 (
    .a(i27[15]),
    .b(sum_26[15]),
    .c(cout_27[14]),
    .cout(cout_27[15]),
    .sum(sum_27[15]));
  AL_FADD comp27_16 (
    .a(i27[16]),
    .b(sum_26[16]),
    .c(cout_27[15]),
    .cout(cout_27[16]),
    .sum(sum_27[16]));
  AL_FADD comp27_17 (
    .a(i27[17]),
    .b(sum_26[17]),
    .c(cout_27[16]),
    .cout(cout_27[17]),
    .sum(sum_27[17]));
  AL_FADD comp27_18 (
    .a(i27[18]),
    .b(sum_26[18]),
    .c(cout_27[17]),
    .cout(cout_27[18]),
    .sum(sum_27[18]));
  AL_FADD comp27_19 (
    .a(i27[19]),
    .b(sum_26[19]),
    .c(cout_27[18]),
    .cout(cout_27[19]),
    .sum(sum_27[19]));
  AL_FADD comp27_2 (
    .a(i27[2]),
    .b(sum_26[2]),
    .c(cout_27[1]),
    .cout(cout_27[2]),
    .sum(sum_27[2]));
  AL_FADD comp27_20 (
    .a(i27[20]),
    .b(sum_26[20]),
    .c(cout_27[19]),
    .cout(cout_27[20]),
    .sum(sum_27[20]));
  AL_FADD comp27_21 (
    .a(i27[21]),
    .b(sum_26[21]),
    .c(cout_27[20]),
    .cout(cout_27[21]),
    .sum(sum_27[21]));
  AL_FADD comp27_22 (
    .a(i27[22]),
    .b(sum_26[22]),
    .c(cout_27[21]),
    .cout(cout_27[22]),
    .sum(sum_27[22]));
  AL_FADD comp27_23 (
    .a(i27[23]),
    .b(sum_26[23]),
    .c(cout_27[22]),
    .cout(cout_27[23]),
    .sum(sum_27[23]));
  AL_FADD comp27_24 (
    .a(i27[24]),
    .b(sum_26[24]),
    .c(cout_27[23]),
    .cout(cout_27[24]),
    .sum(sum_27[24]));
  AL_FADD comp27_25 (
    .a(i27[25]),
    .b(sum_26[25]),
    .c(cout_27[24]),
    .cout(cout_27[25]),
    .sum(sum_27[25]));
  AL_FADD comp27_26 (
    .a(i27[26]),
    .b(sum_26[26]),
    .c(cout_27[25]),
    .cout(cout_27[26]),
    .sum(sum_27[26]));
  AL_FADD comp27_27 (
    .a(i27[27]),
    .b(sum_26[27]),
    .c(cout_27[26]),
    .cout(cout_27[27]),
    .sum(sum_27[27]));
  AL_FADD comp27_28 (
    .a(i27[28]),
    .b(sum_26[28]),
    .c(cout_27[27]),
    .cout(cout_27[28]),
    .sum(sum_27[28]));
  AL_FADD comp27_29 (
    .a(i27[29]),
    .b(sum_26[29]),
    .c(cout_27[28]),
    .cout(cout_27[29]),
    .sum(sum_27[29]));
  AL_FADD comp27_3 (
    .a(i27[3]),
    .b(sum_26[3]),
    .c(cout_27[2]),
    .cout(cout_27[3]),
    .sum(sum_27[3]));
  AL_FADD comp27_30 (
    .a(i27[30]),
    .b(sum_26[30]),
    .c(cout_27[29]),
    .cout(cout_27[30]),
    .sum(sum_27[30]));
  AL_FADD comp27_31 (
    .a(i27[31]),
    .b(sum_26[31]),
    .c(cout_27[30]),
    .cout(cout_27[31]),
    .sum(sum_27[31]));
  AL_FADD comp27_32 (
    .a(i27[32]),
    .b(sum_26[32]),
    .c(cout_27[31]),
    .cout(cout_27[32]),
    .sum(sum_27[32]));
  AL_FADD comp27_33 (
    .a(i27[33]),
    .b(sum_26[33]),
    .c(cout_27[32]),
    .cout(cout_27[33]),
    .sum(sum_27[33]));
  AL_FADD comp27_34 (
    .a(i27[34]),
    .b(sum_26[34]),
    .c(cout_27[33]),
    .cout(cout_27[34]),
    .sum(sum_27[34]));
  AL_FADD comp27_35 (
    .a(i27[35]),
    .b(sum_26[35]),
    .c(cout_27[34]),
    .cout(cout_27[35]),
    .sum(sum_27[35]));
  AL_FADD comp27_36 (
    .a(1'b0),
    .b(sum_26[36]),
    .c(cout_27[35]),
    .cout(cout_27[36]),
    .sum(sum_27[36]));
  AL_FADD comp27_37 (
    .a(1'b0),
    .b(sum_26[37]),
    .c(cout_27[36]),
    .cout(cout_27[37]),
    .sum(sum_27[37]));
  AL_FADD comp27_38 (
    .a(1'b0),
    .b(sum_26[38]),
    .c(cout_27[37]),
    .cout(cout_27[38]),
    .sum(sum_27[38]));
  AL_FADD comp27_39 (
    .a(1'b0),
    .b(sum_26[39]),
    .c(cout_27[38]),
    .cout(cout_27[39]),
    .sum(sum_27[39]));
  AL_FADD comp27_4 (
    .a(i27[4]),
    .b(sum_26[4]),
    .c(cout_27[3]),
    .cout(cout_27[4]),
    .sum(sum_27[4]));
  AL_FADD comp27_40 (
    .a(1'b0),
    .b(sum_26[40]),
    .c(cout_27[39]),
    .cout(cout_27[40]),
    .sum(sum_27[40]));
  AL_FADD comp27_41 (
    .a(1'b0),
    .b(sum_26[41]),
    .c(cout_27[40]),
    .cout(cout_27[41]),
    .sum(sum_27[41]));
  AL_FADD comp27_42 (
    .a(1'b0),
    .b(sum_26[42]),
    .c(cout_27[41]),
    .cout(cout_27[42]),
    .sum(sum_27[42]));
  AL_FADD comp27_43 (
    .a(1'b0),
    .b(sum_26[43]),
    .c(cout_27[42]),
    .cout(cout_27[43]),
    .sum(sum_27[43]));
  AL_FADD comp27_44 (
    .a(1'b0),
    .b(sum_26[44]),
    .c(cout_27[43]),
    .cout(cout_27[44]),
    .sum(sum_27[44]));
  AL_FADD comp27_45 (
    .a(1'b0),
    .b(sum_26[45]),
    .c(cout_27[44]),
    .cout(cout_27[45]),
    .sum(sum_27[45]));
  AL_FADD comp27_46 (
    .a(1'b0),
    .b(sum_26[46]),
    .c(cout_27[45]),
    .cout(cout_27[46]),
    .sum(sum_27[46]));
  AL_FADD comp27_47 (
    .a(1'b0),
    .b(sum_26[47]),
    .c(cout_27[46]),
    .cout(cout_27[47]),
    .sum(sum_27[47]));
  AL_FADD comp27_48 (
    .a(1'b0),
    .b(sum_26[48]),
    .c(cout_27[47]),
    .cout(cout_27[48]),
    .sum(sum_27[48]));
  AL_FADD comp27_49 (
    .a(1'b0),
    .b(sum_26[49]),
    .c(cout_27[48]),
    .cout(cout_27[49]),
    .sum(sum_27[49]));
  AL_FADD comp27_5 (
    .a(i27[5]),
    .b(sum_26[5]),
    .c(cout_27[4]),
    .cout(cout_27[5]),
    .sum(sum_27[5]));
  AL_FADD comp27_50 (
    .a(1'b0),
    .b(sum_26[50]),
    .c(cout_27[49]),
    .cout(cout_27[50]),
    .sum(sum_27[50]));
  AL_FADD comp27_51 (
    .a(1'b0),
    .b(sum_26[51]),
    .c(cout_27[50]),
    .cout(cout_27[51]),
    .sum(sum_27[51]));
  AL_FADD comp27_52 (
    .a(1'b0),
    .b(sum_26[52]),
    .c(cout_27[51]),
    .cout(cout_27[52]),
    .sum(sum_27[52]));
  AL_FADD comp27_53 (
    .a(1'b0),
    .b(sum_26[53]),
    .c(cout_27[52]),
    .cout(cout_27[53]),
    .sum(sum_27[53]));
  AL_FADD comp27_54 (
    .a(1'b0),
    .b(sum_26[54]),
    .c(cout_27[53]),
    .cout(cout_27[54]),
    .sum(sum_27[54]));
  AL_FADD comp27_55 (
    .a(1'b0),
    .b(sum_26[55]),
    .c(cout_27[54]),
    .cout(cout_27[55]),
    .sum(sum_27[55]));
  AL_FADD comp27_56 (
    .a(1'b0),
    .b(sum_26[56]),
    .c(cout_27[55]),
    .cout(cout_27[56]),
    .sum(sum_27[56]));
  AL_FADD comp27_57 (
    .a(1'b0),
    .b(sum_26[57]),
    .c(cout_27[56]),
    .cout(cout_27[57]),
    .sum(sum_27[57]));
  AL_FADD comp27_58 (
    .a(1'b0),
    .b(sum_26[58]),
    .c(cout_27[57]),
    .cout(cout_27[58]),
    .sum(sum_27[58]));
  AL_FADD comp27_59 (
    .a(1'b0),
    .b(sum_26[59]),
    .c(cout_27[58]),
    .cout(cout_27[59]),
    .sum(sum_27[59]));
  AL_FADD comp27_6 (
    .a(i27[6]),
    .b(sum_26[6]),
    .c(cout_27[5]),
    .cout(cout_27[6]),
    .sum(sum_27[6]));
  AL_FADD comp27_60 (
    .a(1'b0),
    .b(sum_26[60]),
    .c(cout_27[59]),
    .cout(cout_27[60]),
    .sum(sum_27[60]));
  AL_FADD comp27_61 (
    .a(1'b0),
    .b(sum_26[61]),
    .c(cout_27[60]),
    .cout(cout_27[61]),
    .sum(sum_27[61]));
  AL_FADD comp27_62 (
    .a(1'b0),
    .b(sum_26[62]),
    .c(cout_27[61]),
    .cout(cout_27[62]),
    .sum(sum_27[62]));
  AL_FADD comp27_63 (
    .a(1'b0),
    .b(sum_26[63]),
    .c(cout_27[62]),
    .cout(cout_27[63]),
    .sum(sum_27[63]));
  AL_FADD comp27_7 (
    .a(i27[7]),
    .b(sum_26[7]),
    .c(cout_27[6]),
    .cout(cout_27[7]),
    .sum(sum_27[7]));
  AL_FADD comp27_8 (
    .a(i27[8]),
    .b(sum_26[8]),
    .c(cout_27[7]),
    .cout(cout_27[8]),
    .sum(sum_27[8]));
  AL_FADD comp27_9 (
    .a(i27[9]),
    .b(sum_26[9]),
    .c(cout_27[8]),
    .cout(cout_27[9]),
    .sum(sum_27[9]));
  AL_FADD comp28_0 (
    .a(i28[0]),
    .b(sum_27[0]),
    .c(1'b0),
    .cout(cout_28[0]),
    .sum(sum_28[0]));
  AL_FADD comp28_1 (
    .a(i28[1]),
    .b(sum_27[1]),
    .c(cout_28[0]),
    .cout(cout_28[1]),
    .sum(sum_28[1]));
  AL_FADD comp28_10 (
    .a(i28[10]),
    .b(sum_27[10]),
    .c(cout_28[9]),
    .cout(cout_28[10]),
    .sum(sum_28[10]));
  AL_FADD comp28_11 (
    .a(i28[11]),
    .b(sum_27[11]),
    .c(cout_28[10]),
    .cout(cout_28[11]),
    .sum(sum_28[11]));
  AL_FADD comp28_12 (
    .a(i28[12]),
    .b(sum_27[12]),
    .c(cout_28[11]),
    .cout(cout_28[12]),
    .sum(sum_28[12]));
  AL_FADD comp28_13 (
    .a(i28[13]),
    .b(sum_27[13]),
    .c(cout_28[12]),
    .cout(cout_28[13]),
    .sum(sum_28[13]));
  AL_FADD comp28_14 (
    .a(i28[14]),
    .b(sum_27[14]),
    .c(cout_28[13]),
    .cout(cout_28[14]),
    .sum(sum_28[14]));
  AL_FADD comp28_15 (
    .a(i28[15]),
    .b(sum_27[15]),
    .c(cout_28[14]),
    .cout(cout_28[15]),
    .sum(sum_28[15]));
  AL_FADD comp28_16 (
    .a(i28[16]),
    .b(sum_27[16]),
    .c(cout_28[15]),
    .cout(cout_28[16]),
    .sum(sum_28[16]));
  AL_FADD comp28_17 (
    .a(i28[17]),
    .b(sum_27[17]),
    .c(cout_28[16]),
    .cout(cout_28[17]),
    .sum(sum_28[17]));
  AL_FADD comp28_18 (
    .a(i28[18]),
    .b(sum_27[18]),
    .c(cout_28[17]),
    .cout(cout_28[18]),
    .sum(sum_28[18]));
  AL_FADD comp28_19 (
    .a(i28[19]),
    .b(sum_27[19]),
    .c(cout_28[18]),
    .cout(cout_28[19]),
    .sum(sum_28[19]));
  AL_FADD comp28_2 (
    .a(i28[2]),
    .b(sum_27[2]),
    .c(cout_28[1]),
    .cout(cout_28[2]),
    .sum(sum_28[2]));
  AL_FADD comp28_20 (
    .a(i28[20]),
    .b(sum_27[20]),
    .c(cout_28[19]),
    .cout(cout_28[20]),
    .sum(sum_28[20]));
  AL_FADD comp28_21 (
    .a(i28[21]),
    .b(sum_27[21]),
    .c(cout_28[20]),
    .cout(cout_28[21]),
    .sum(sum_28[21]));
  AL_FADD comp28_22 (
    .a(i28[22]),
    .b(sum_27[22]),
    .c(cout_28[21]),
    .cout(cout_28[22]),
    .sum(sum_28[22]));
  AL_FADD comp28_23 (
    .a(i28[23]),
    .b(sum_27[23]),
    .c(cout_28[22]),
    .cout(cout_28[23]),
    .sum(sum_28[23]));
  AL_FADD comp28_24 (
    .a(i28[24]),
    .b(sum_27[24]),
    .c(cout_28[23]),
    .cout(cout_28[24]),
    .sum(sum_28[24]));
  AL_FADD comp28_25 (
    .a(i28[25]),
    .b(sum_27[25]),
    .c(cout_28[24]),
    .cout(cout_28[25]),
    .sum(sum_28[25]));
  AL_FADD comp28_26 (
    .a(i28[26]),
    .b(sum_27[26]),
    .c(cout_28[25]),
    .cout(cout_28[26]),
    .sum(sum_28[26]));
  AL_FADD comp28_27 (
    .a(i28[27]),
    .b(sum_27[27]),
    .c(cout_28[26]),
    .cout(cout_28[27]),
    .sum(sum_28[27]));
  AL_FADD comp28_28 (
    .a(i28[28]),
    .b(sum_27[28]),
    .c(cout_28[27]),
    .cout(cout_28[28]),
    .sum(sum_28[28]));
  AL_FADD comp28_29 (
    .a(i28[29]),
    .b(sum_27[29]),
    .c(cout_28[28]),
    .cout(cout_28[29]),
    .sum(sum_28[29]));
  AL_FADD comp28_3 (
    .a(i28[3]),
    .b(sum_27[3]),
    .c(cout_28[2]),
    .cout(cout_28[3]),
    .sum(sum_28[3]));
  AL_FADD comp28_30 (
    .a(i28[30]),
    .b(sum_27[30]),
    .c(cout_28[29]),
    .cout(cout_28[30]),
    .sum(sum_28[30]));
  AL_FADD comp28_31 (
    .a(i28[31]),
    .b(sum_27[31]),
    .c(cout_28[30]),
    .cout(cout_28[31]),
    .sum(sum_28[31]));
  AL_FADD comp28_32 (
    .a(i28[32]),
    .b(sum_27[32]),
    .c(cout_28[31]),
    .cout(cout_28[32]),
    .sum(sum_28[32]));
  AL_FADD comp28_33 (
    .a(i28[33]),
    .b(sum_27[33]),
    .c(cout_28[32]),
    .cout(cout_28[33]),
    .sum(sum_28[33]));
  AL_FADD comp28_34 (
    .a(i28[34]),
    .b(sum_27[34]),
    .c(cout_28[33]),
    .cout(cout_28[34]),
    .sum(sum_28[34]));
  AL_FADD comp28_35 (
    .a(1'b0),
    .b(sum_27[35]),
    .c(cout_28[34]),
    .cout(cout_28[35]),
    .sum(sum_28[35]));
  AL_FADD comp28_36 (
    .a(1'b0),
    .b(sum_27[36]),
    .c(cout_28[35]),
    .cout(cout_28[36]),
    .sum(sum_28[36]));
  AL_FADD comp28_37 (
    .a(1'b0),
    .b(sum_27[37]),
    .c(cout_28[36]),
    .cout(cout_28[37]),
    .sum(sum_28[37]));
  AL_FADD comp28_38 (
    .a(1'b0),
    .b(sum_27[38]),
    .c(cout_28[37]),
    .cout(cout_28[38]),
    .sum(sum_28[38]));
  AL_FADD comp28_39 (
    .a(1'b0),
    .b(sum_27[39]),
    .c(cout_28[38]),
    .cout(cout_28[39]),
    .sum(sum_28[39]));
  AL_FADD comp28_4 (
    .a(i28[4]),
    .b(sum_27[4]),
    .c(cout_28[3]),
    .cout(cout_28[4]),
    .sum(sum_28[4]));
  AL_FADD comp28_40 (
    .a(1'b0),
    .b(sum_27[40]),
    .c(cout_28[39]),
    .cout(cout_28[40]),
    .sum(sum_28[40]));
  AL_FADD comp28_41 (
    .a(1'b0),
    .b(sum_27[41]),
    .c(cout_28[40]),
    .cout(cout_28[41]),
    .sum(sum_28[41]));
  AL_FADD comp28_42 (
    .a(1'b0),
    .b(sum_27[42]),
    .c(cout_28[41]),
    .cout(cout_28[42]),
    .sum(sum_28[42]));
  AL_FADD comp28_43 (
    .a(1'b0),
    .b(sum_27[43]),
    .c(cout_28[42]),
    .cout(cout_28[43]),
    .sum(sum_28[43]));
  AL_FADD comp28_44 (
    .a(1'b0),
    .b(sum_27[44]),
    .c(cout_28[43]),
    .cout(cout_28[44]),
    .sum(sum_28[44]));
  AL_FADD comp28_45 (
    .a(1'b0),
    .b(sum_27[45]),
    .c(cout_28[44]),
    .cout(cout_28[45]),
    .sum(sum_28[45]));
  AL_FADD comp28_46 (
    .a(1'b0),
    .b(sum_27[46]),
    .c(cout_28[45]),
    .cout(cout_28[46]),
    .sum(sum_28[46]));
  AL_FADD comp28_47 (
    .a(1'b0),
    .b(sum_27[47]),
    .c(cout_28[46]),
    .cout(cout_28[47]),
    .sum(sum_28[47]));
  AL_FADD comp28_48 (
    .a(1'b0),
    .b(sum_27[48]),
    .c(cout_28[47]),
    .cout(cout_28[48]),
    .sum(sum_28[48]));
  AL_FADD comp28_49 (
    .a(1'b0),
    .b(sum_27[49]),
    .c(cout_28[48]),
    .cout(cout_28[49]),
    .sum(sum_28[49]));
  AL_FADD comp28_5 (
    .a(i28[5]),
    .b(sum_27[5]),
    .c(cout_28[4]),
    .cout(cout_28[5]),
    .sum(sum_28[5]));
  AL_FADD comp28_50 (
    .a(1'b0),
    .b(sum_27[50]),
    .c(cout_28[49]),
    .cout(cout_28[50]),
    .sum(sum_28[50]));
  AL_FADD comp28_51 (
    .a(1'b0),
    .b(sum_27[51]),
    .c(cout_28[50]),
    .cout(cout_28[51]),
    .sum(sum_28[51]));
  AL_FADD comp28_52 (
    .a(1'b0),
    .b(sum_27[52]),
    .c(cout_28[51]),
    .cout(cout_28[52]),
    .sum(sum_28[52]));
  AL_FADD comp28_53 (
    .a(1'b0),
    .b(sum_27[53]),
    .c(cout_28[52]),
    .cout(cout_28[53]),
    .sum(sum_28[53]));
  AL_FADD comp28_54 (
    .a(1'b0),
    .b(sum_27[54]),
    .c(cout_28[53]),
    .cout(cout_28[54]),
    .sum(sum_28[54]));
  AL_FADD comp28_55 (
    .a(1'b0),
    .b(sum_27[55]),
    .c(cout_28[54]),
    .cout(cout_28[55]),
    .sum(sum_28[55]));
  AL_FADD comp28_56 (
    .a(1'b0),
    .b(sum_27[56]),
    .c(cout_28[55]),
    .cout(cout_28[56]),
    .sum(sum_28[56]));
  AL_FADD comp28_57 (
    .a(1'b0),
    .b(sum_27[57]),
    .c(cout_28[56]),
    .cout(cout_28[57]),
    .sum(sum_28[57]));
  AL_FADD comp28_58 (
    .a(1'b0),
    .b(sum_27[58]),
    .c(cout_28[57]),
    .cout(cout_28[58]),
    .sum(sum_28[58]));
  AL_FADD comp28_59 (
    .a(1'b0),
    .b(sum_27[59]),
    .c(cout_28[58]),
    .cout(cout_28[59]),
    .sum(sum_28[59]));
  AL_FADD comp28_6 (
    .a(i28[6]),
    .b(sum_27[6]),
    .c(cout_28[5]),
    .cout(cout_28[6]),
    .sum(sum_28[6]));
  AL_FADD comp28_60 (
    .a(1'b0),
    .b(sum_27[60]),
    .c(cout_28[59]),
    .cout(cout_28[60]),
    .sum(sum_28[60]));
  AL_FADD comp28_61 (
    .a(1'b0),
    .b(sum_27[61]),
    .c(cout_28[60]),
    .cout(cout_28[61]),
    .sum(sum_28[61]));
  AL_FADD comp28_62 (
    .a(1'b0),
    .b(sum_27[62]),
    .c(cout_28[61]),
    .cout(cout_28[62]),
    .sum(sum_28[62]));
  AL_FADD comp28_63 (
    .a(1'b0),
    .b(sum_27[63]),
    .c(cout_28[62]),
    .cout(cout_28[63]),
    .sum(sum_28[63]));
  AL_FADD comp28_7 (
    .a(i28[7]),
    .b(sum_27[7]),
    .c(cout_28[6]),
    .cout(cout_28[7]),
    .sum(sum_28[7]));
  AL_FADD comp28_8 (
    .a(i28[8]),
    .b(sum_27[8]),
    .c(cout_28[7]),
    .cout(cout_28[8]),
    .sum(sum_28[8]));
  AL_FADD comp28_9 (
    .a(i28[9]),
    .b(sum_27[9]),
    .c(cout_28[8]),
    .cout(cout_28[9]),
    .sum(sum_28[9]));
  AL_FADD comp29_0 (
    .a(i29[0]),
    .b(sum_28[0]),
    .c(1'b0),
    .cout(cout_29[0]),
    .sum(sum_29[0]));
  AL_FADD comp29_1 (
    .a(i29[1]),
    .b(sum_28[1]),
    .c(cout_29[0]),
    .cout(cout_29[1]),
    .sum(sum_29[1]));
  AL_FADD comp29_10 (
    .a(i29[10]),
    .b(sum_28[10]),
    .c(cout_29[9]),
    .cout(cout_29[10]),
    .sum(sum_29[10]));
  AL_FADD comp29_11 (
    .a(i29[11]),
    .b(sum_28[11]),
    .c(cout_29[10]),
    .cout(cout_29[11]),
    .sum(sum_29[11]));
  AL_FADD comp29_12 (
    .a(i29[12]),
    .b(sum_28[12]),
    .c(cout_29[11]),
    .cout(cout_29[12]),
    .sum(sum_29[12]));
  AL_FADD comp29_13 (
    .a(i29[13]),
    .b(sum_28[13]),
    .c(cout_29[12]),
    .cout(cout_29[13]),
    .sum(sum_29[13]));
  AL_FADD comp29_14 (
    .a(i29[14]),
    .b(sum_28[14]),
    .c(cout_29[13]),
    .cout(cout_29[14]),
    .sum(sum_29[14]));
  AL_FADD comp29_15 (
    .a(i29[15]),
    .b(sum_28[15]),
    .c(cout_29[14]),
    .cout(cout_29[15]),
    .sum(sum_29[15]));
  AL_FADD comp29_16 (
    .a(i29[16]),
    .b(sum_28[16]),
    .c(cout_29[15]),
    .cout(cout_29[16]),
    .sum(sum_29[16]));
  AL_FADD comp29_17 (
    .a(i29[17]),
    .b(sum_28[17]),
    .c(cout_29[16]),
    .cout(cout_29[17]),
    .sum(sum_29[17]));
  AL_FADD comp29_18 (
    .a(i29[18]),
    .b(sum_28[18]),
    .c(cout_29[17]),
    .cout(cout_29[18]),
    .sum(sum_29[18]));
  AL_FADD comp29_19 (
    .a(i29[19]),
    .b(sum_28[19]),
    .c(cout_29[18]),
    .cout(cout_29[19]),
    .sum(sum_29[19]));
  AL_FADD comp29_2 (
    .a(i29[2]),
    .b(sum_28[2]),
    .c(cout_29[1]),
    .cout(cout_29[2]),
    .sum(sum_29[2]));
  AL_FADD comp29_20 (
    .a(i29[20]),
    .b(sum_28[20]),
    .c(cout_29[19]),
    .cout(cout_29[20]),
    .sum(sum_29[20]));
  AL_FADD comp29_21 (
    .a(i29[21]),
    .b(sum_28[21]),
    .c(cout_29[20]),
    .cout(cout_29[21]),
    .sum(sum_29[21]));
  AL_FADD comp29_22 (
    .a(i29[22]),
    .b(sum_28[22]),
    .c(cout_29[21]),
    .cout(cout_29[22]),
    .sum(sum_29[22]));
  AL_FADD comp29_23 (
    .a(i29[23]),
    .b(sum_28[23]),
    .c(cout_29[22]),
    .cout(cout_29[23]),
    .sum(sum_29[23]));
  AL_FADD comp29_24 (
    .a(i29[24]),
    .b(sum_28[24]),
    .c(cout_29[23]),
    .cout(cout_29[24]),
    .sum(sum_29[24]));
  AL_FADD comp29_25 (
    .a(i29[25]),
    .b(sum_28[25]),
    .c(cout_29[24]),
    .cout(cout_29[25]),
    .sum(sum_29[25]));
  AL_FADD comp29_26 (
    .a(i29[26]),
    .b(sum_28[26]),
    .c(cout_29[25]),
    .cout(cout_29[26]),
    .sum(sum_29[26]));
  AL_FADD comp29_27 (
    .a(i29[27]),
    .b(sum_28[27]),
    .c(cout_29[26]),
    .cout(cout_29[27]),
    .sum(sum_29[27]));
  AL_FADD comp29_28 (
    .a(i29[28]),
    .b(sum_28[28]),
    .c(cout_29[27]),
    .cout(cout_29[28]),
    .sum(sum_29[28]));
  AL_FADD comp29_29 (
    .a(i29[29]),
    .b(sum_28[29]),
    .c(cout_29[28]),
    .cout(cout_29[29]),
    .sum(sum_29[29]));
  AL_FADD comp29_3 (
    .a(i29[3]),
    .b(sum_28[3]),
    .c(cout_29[2]),
    .cout(cout_29[3]),
    .sum(sum_29[3]));
  AL_FADD comp29_30 (
    .a(i29[30]),
    .b(sum_28[30]),
    .c(cout_29[29]),
    .cout(cout_29[30]),
    .sum(sum_29[30]));
  AL_FADD comp29_31 (
    .a(i29[31]),
    .b(sum_28[31]),
    .c(cout_29[30]),
    .cout(cout_29[31]),
    .sum(sum_29[31]));
  AL_FADD comp29_32 (
    .a(i29[32]),
    .b(sum_28[32]),
    .c(cout_29[31]),
    .cout(cout_29[32]),
    .sum(sum_29[32]));
  AL_FADD comp29_33 (
    .a(i29[33]),
    .b(sum_28[33]),
    .c(cout_29[32]),
    .cout(cout_29[33]),
    .sum(sum_29[33]));
  AL_FADD comp29_34 (
    .a(1'b0),
    .b(sum_28[34]),
    .c(cout_29[33]),
    .cout(cout_29[34]),
    .sum(sum_29[34]));
  AL_FADD comp29_35 (
    .a(1'b0),
    .b(sum_28[35]),
    .c(cout_29[34]),
    .cout(cout_29[35]),
    .sum(sum_29[35]));
  AL_FADD comp29_36 (
    .a(1'b0),
    .b(sum_28[36]),
    .c(cout_29[35]),
    .cout(cout_29[36]),
    .sum(sum_29[36]));
  AL_FADD comp29_37 (
    .a(1'b0),
    .b(sum_28[37]),
    .c(cout_29[36]),
    .cout(cout_29[37]),
    .sum(sum_29[37]));
  AL_FADD comp29_38 (
    .a(1'b0),
    .b(sum_28[38]),
    .c(cout_29[37]),
    .cout(cout_29[38]),
    .sum(sum_29[38]));
  AL_FADD comp29_39 (
    .a(1'b0),
    .b(sum_28[39]),
    .c(cout_29[38]),
    .cout(cout_29[39]),
    .sum(sum_29[39]));
  AL_FADD comp29_4 (
    .a(i29[4]),
    .b(sum_28[4]),
    .c(cout_29[3]),
    .cout(cout_29[4]),
    .sum(sum_29[4]));
  AL_FADD comp29_40 (
    .a(1'b0),
    .b(sum_28[40]),
    .c(cout_29[39]),
    .cout(cout_29[40]),
    .sum(sum_29[40]));
  AL_FADD comp29_41 (
    .a(1'b0),
    .b(sum_28[41]),
    .c(cout_29[40]),
    .cout(cout_29[41]),
    .sum(sum_29[41]));
  AL_FADD comp29_42 (
    .a(1'b0),
    .b(sum_28[42]),
    .c(cout_29[41]),
    .cout(cout_29[42]),
    .sum(sum_29[42]));
  AL_FADD comp29_43 (
    .a(1'b0),
    .b(sum_28[43]),
    .c(cout_29[42]),
    .cout(cout_29[43]),
    .sum(sum_29[43]));
  AL_FADD comp29_44 (
    .a(1'b0),
    .b(sum_28[44]),
    .c(cout_29[43]),
    .cout(cout_29[44]),
    .sum(sum_29[44]));
  AL_FADD comp29_45 (
    .a(1'b0),
    .b(sum_28[45]),
    .c(cout_29[44]),
    .cout(cout_29[45]),
    .sum(sum_29[45]));
  AL_FADD comp29_46 (
    .a(1'b0),
    .b(sum_28[46]),
    .c(cout_29[45]),
    .cout(cout_29[46]),
    .sum(sum_29[46]));
  AL_FADD comp29_47 (
    .a(1'b0),
    .b(sum_28[47]),
    .c(cout_29[46]),
    .cout(cout_29[47]),
    .sum(sum_29[47]));
  AL_FADD comp29_48 (
    .a(1'b0),
    .b(sum_28[48]),
    .c(cout_29[47]),
    .cout(cout_29[48]),
    .sum(sum_29[48]));
  AL_FADD comp29_49 (
    .a(1'b0),
    .b(sum_28[49]),
    .c(cout_29[48]),
    .cout(cout_29[49]),
    .sum(sum_29[49]));
  AL_FADD comp29_5 (
    .a(i29[5]),
    .b(sum_28[5]),
    .c(cout_29[4]),
    .cout(cout_29[5]),
    .sum(sum_29[5]));
  AL_FADD comp29_50 (
    .a(1'b0),
    .b(sum_28[50]),
    .c(cout_29[49]),
    .cout(cout_29[50]),
    .sum(sum_29[50]));
  AL_FADD comp29_51 (
    .a(1'b0),
    .b(sum_28[51]),
    .c(cout_29[50]),
    .cout(cout_29[51]),
    .sum(sum_29[51]));
  AL_FADD comp29_52 (
    .a(1'b0),
    .b(sum_28[52]),
    .c(cout_29[51]),
    .cout(cout_29[52]),
    .sum(sum_29[52]));
  AL_FADD comp29_53 (
    .a(1'b0),
    .b(sum_28[53]),
    .c(cout_29[52]),
    .cout(cout_29[53]),
    .sum(sum_29[53]));
  AL_FADD comp29_54 (
    .a(1'b0),
    .b(sum_28[54]),
    .c(cout_29[53]),
    .cout(cout_29[54]),
    .sum(sum_29[54]));
  AL_FADD comp29_55 (
    .a(1'b0),
    .b(sum_28[55]),
    .c(cout_29[54]),
    .cout(cout_29[55]),
    .sum(sum_29[55]));
  AL_FADD comp29_56 (
    .a(1'b0),
    .b(sum_28[56]),
    .c(cout_29[55]),
    .cout(cout_29[56]),
    .sum(sum_29[56]));
  AL_FADD comp29_57 (
    .a(1'b0),
    .b(sum_28[57]),
    .c(cout_29[56]),
    .cout(cout_29[57]),
    .sum(sum_29[57]));
  AL_FADD comp29_58 (
    .a(1'b0),
    .b(sum_28[58]),
    .c(cout_29[57]),
    .cout(cout_29[58]),
    .sum(sum_29[58]));
  AL_FADD comp29_59 (
    .a(1'b0),
    .b(sum_28[59]),
    .c(cout_29[58]),
    .cout(cout_29[59]),
    .sum(sum_29[59]));
  AL_FADD comp29_6 (
    .a(i29[6]),
    .b(sum_28[6]),
    .c(cout_29[5]),
    .cout(cout_29[6]),
    .sum(sum_29[6]));
  AL_FADD comp29_60 (
    .a(1'b0),
    .b(sum_28[60]),
    .c(cout_29[59]),
    .cout(cout_29[60]),
    .sum(sum_29[60]));
  AL_FADD comp29_61 (
    .a(1'b0),
    .b(sum_28[61]),
    .c(cout_29[60]),
    .cout(cout_29[61]),
    .sum(sum_29[61]));
  AL_FADD comp29_62 (
    .a(1'b0),
    .b(sum_28[62]),
    .c(cout_29[61]),
    .cout(cout_29[62]),
    .sum(sum_29[62]));
  AL_FADD comp29_63 (
    .a(1'b0),
    .b(sum_28[63]),
    .c(cout_29[62]),
    .cout(cout_29[63]),
    .sum(sum_29[63]));
  AL_FADD comp29_7 (
    .a(i29[7]),
    .b(sum_28[7]),
    .c(cout_29[6]),
    .cout(cout_29[7]),
    .sum(sum_29[7]));
  AL_FADD comp29_8 (
    .a(i29[8]),
    .b(sum_28[8]),
    .c(cout_29[7]),
    .cout(cout_29[8]),
    .sum(sum_29[8]));
  AL_FADD comp29_9 (
    .a(i29[9]),
    .b(sum_28[9]),
    .c(cout_29[8]),
    .cout(cout_29[9]),
    .sum(sum_29[9]));
  AL_FADD comp2_0 (
    .a(i2[0]),
    .b(sum_1[0]),
    .c(1'b0),
    .cout(cout_2[0]),
    .sum(sum_2[0]));
  AL_FADD comp2_1 (
    .a(i2[1]),
    .b(sum_1[1]),
    .c(cout_2[0]),
    .cout(cout_2[1]),
    .sum(sum_2[1]));
  AL_FADD comp2_10 (
    .a(i2[10]),
    .b(sum_1[10]),
    .c(cout_2[9]),
    .cout(cout_2[10]),
    .sum(sum_2[10]));
  AL_FADD comp2_11 (
    .a(i2[11]),
    .b(sum_1[11]),
    .c(cout_2[10]),
    .cout(cout_2[11]),
    .sum(sum_2[11]));
  AL_FADD comp2_12 (
    .a(i2[12]),
    .b(sum_1[12]),
    .c(cout_2[11]),
    .cout(cout_2[12]),
    .sum(sum_2[12]));
  AL_FADD comp2_13 (
    .a(i2[13]),
    .b(sum_1[13]),
    .c(cout_2[12]),
    .cout(cout_2[13]),
    .sum(sum_2[13]));
  AL_FADD comp2_14 (
    .a(i2[14]),
    .b(sum_1[14]),
    .c(cout_2[13]),
    .cout(cout_2[14]),
    .sum(sum_2[14]));
  AL_FADD comp2_15 (
    .a(i2[15]),
    .b(sum_1[15]),
    .c(cout_2[14]),
    .cout(cout_2[15]),
    .sum(sum_2[15]));
  AL_FADD comp2_16 (
    .a(i2[16]),
    .b(sum_1[16]),
    .c(cout_2[15]),
    .cout(cout_2[16]),
    .sum(sum_2[16]));
  AL_FADD comp2_17 (
    .a(i2[17]),
    .b(sum_1[17]),
    .c(cout_2[16]),
    .cout(cout_2[17]),
    .sum(sum_2[17]));
  AL_FADD comp2_18 (
    .a(i2[18]),
    .b(sum_1[18]),
    .c(cout_2[17]),
    .cout(cout_2[18]),
    .sum(sum_2[18]));
  AL_FADD comp2_19 (
    .a(i2[19]),
    .b(sum_1[19]),
    .c(cout_2[18]),
    .cout(cout_2[19]),
    .sum(sum_2[19]));
  AL_FADD comp2_2 (
    .a(i2[2]),
    .b(sum_1[2]),
    .c(cout_2[1]),
    .cout(cout_2[2]),
    .sum(sum_2[2]));
  AL_FADD comp2_20 (
    .a(i2[20]),
    .b(sum_1[20]),
    .c(cout_2[19]),
    .cout(cout_2[20]),
    .sum(sum_2[20]));
  AL_FADD comp2_21 (
    .a(i2[21]),
    .b(sum_1[21]),
    .c(cout_2[20]),
    .cout(cout_2[21]),
    .sum(sum_2[21]));
  AL_FADD comp2_22 (
    .a(i2[22]),
    .b(sum_1[22]),
    .c(cout_2[21]),
    .cout(cout_2[22]),
    .sum(sum_2[22]));
  AL_FADD comp2_23 (
    .a(i2[23]),
    .b(sum_1[23]),
    .c(cout_2[22]),
    .cout(cout_2[23]),
    .sum(sum_2[23]));
  AL_FADD comp2_24 (
    .a(i2[24]),
    .b(sum_1[24]),
    .c(cout_2[23]),
    .cout(cout_2[24]),
    .sum(sum_2[24]));
  AL_FADD comp2_25 (
    .a(i2[25]),
    .b(sum_1[25]),
    .c(cout_2[24]),
    .cout(cout_2[25]),
    .sum(sum_2[25]));
  AL_FADD comp2_26 (
    .a(i2[26]),
    .b(sum_1[26]),
    .c(cout_2[25]),
    .cout(cout_2[26]),
    .sum(sum_2[26]));
  AL_FADD comp2_27 (
    .a(i2[27]),
    .b(sum_1[27]),
    .c(cout_2[26]),
    .cout(cout_2[27]),
    .sum(sum_2[27]));
  AL_FADD comp2_28 (
    .a(i2[28]),
    .b(sum_1[28]),
    .c(cout_2[27]),
    .cout(cout_2[28]),
    .sum(sum_2[28]));
  AL_FADD comp2_29 (
    .a(i2[29]),
    .b(sum_1[29]),
    .c(cout_2[28]),
    .cout(cout_2[29]),
    .sum(sum_2[29]));
  AL_FADD comp2_3 (
    .a(i2[3]),
    .b(sum_1[3]),
    .c(cout_2[2]),
    .cout(cout_2[3]),
    .sum(sum_2[3]));
  AL_FADD comp2_30 (
    .a(i2[30]),
    .b(sum_1[30]),
    .c(cout_2[29]),
    .cout(cout_2[30]),
    .sum(sum_2[30]));
  AL_FADD comp2_31 (
    .a(i2[31]),
    .b(sum_1[31]),
    .c(cout_2[30]),
    .cout(cout_2[31]),
    .sum(sum_2[31]));
  AL_FADD comp2_32 (
    .a(i2[32]),
    .b(sum_1[32]),
    .c(cout_2[31]),
    .cout(cout_2[32]),
    .sum(sum_2[32]));
  AL_FADD comp2_33 (
    .a(i2[33]),
    .b(sum_1[33]),
    .c(cout_2[32]),
    .cout(cout_2[33]),
    .sum(sum_2[33]));
  AL_FADD comp2_34 (
    .a(i2[34]),
    .b(sum_1[34]),
    .c(cout_2[33]),
    .cout(cout_2[34]),
    .sum(sum_2[34]));
  AL_FADD comp2_35 (
    .a(i2[35]),
    .b(sum_1[35]),
    .c(cout_2[34]),
    .cout(cout_2[35]),
    .sum(sum_2[35]));
  AL_FADD comp2_36 (
    .a(i2[36]),
    .b(sum_1[36]),
    .c(cout_2[35]),
    .cout(cout_2[36]),
    .sum(sum_2[36]));
  AL_FADD comp2_37 (
    .a(i2[37]),
    .b(sum_1[37]),
    .c(cout_2[36]),
    .cout(cout_2[37]),
    .sum(sum_2[37]));
  AL_FADD comp2_38 (
    .a(i2[38]),
    .b(sum_1[38]),
    .c(cout_2[37]),
    .cout(cout_2[38]),
    .sum(sum_2[38]));
  AL_FADD comp2_39 (
    .a(i2[39]),
    .b(sum_1[39]),
    .c(cout_2[38]),
    .cout(cout_2[39]),
    .sum(sum_2[39]));
  AL_FADD comp2_4 (
    .a(i2[4]),
    .b(sum_1[4]),
    .c(cout_2[3]),
    .cout(cout_2[4]),
    .sum(sum_2[4]));
  AL_FADD comp2_40 (
    .a(i2[40]),
    .b(sum_1[40]),
    .c(cout_2[39]),
    .cout(cout_2[40]),
    .sum(sum_2[40]));
  AL_FADD comp2_41 (
    .a(i2[41]),
    .b(sum_1[41]),
    .c(cout_2[40]),
    .cout(cout_2[41]),
    .sum(sum_2[41]));
  AL_FADD comp2_42 (
    .a(i2[42]),
    .b(sum_1[42]),
    .c(cout_2[41]),
    .cout(cout_2[42]),
    .sum(sum_2[42]));
  AL_FADD comp2_43 (
    .a(i2[43]),
    .b(sum_1[43]),
    .c(cout_2[42]),
    .cout(cout_2[43]),
    .sum(sum_2[43]));
  AL_FADD comp2_44 (
    .a(i2[44]),
    .b(sum_1[44]),
    .c(cout_2[43]),
    .cout(cout_2[44]),
    .sum(sum_2[44]));
  AL_FADD comp2_45 (
    .a(i2[45]),
    .b(sum_1[45]),
    .c(cout_2[44]),
    .cout(cout_2[45]),
    .sum(sum_2[45]));
  AL_FADD comp2_46 (
    .a(i2[46]),
    .b(sum_1[46]),
    .c(cout_2[45]),
    .cout(cout_2[46]),
    .sum(sum_2[46]));
  AL_FADD comp2_47 (
    .a(i2[47]),
    .b(sum_1[47]),
    .c(cout_2[46]),
    .cout(cout_2[47]),
    .sum(sum_2[47]));
  AL_FADD comp2_48 (
    .a(i2[48]),
    .b(sum_1[48]),
    .c(cout_2[47]),
    .cout(cout_2[48]),
    .sum(sum_2[48]));
  AL_FADD comp2_49 (
    .a(i2[49]),
    .b(sum_1[49]),
    .c(cout_2[48]),
    .cout(cout_2[49]),
    .sum(sum_2[49]));
  AL_FADD comp2_5 (
    .a(i2[5]),
    .b(sum_1[5]),
    .c(cout_2[4]),
    .cout(cout_2[5]),
    .sum(sum_2[5]));
  AL_FADD comp2_50 (
    .a(i2[50]),
    .b(sum_1[50]),
    .c(cout_2[49]),
    .cout(cout_2[50]),
    .sum(sum_2[50]));
  AL_FADD comp2_51 (
    .a(i2[51]),
    .b(sum_1[51]),
    .c(cout_2[50]),
    .cout(cout_2[51]),
    .sum(sum_2[51]));
  AL_FADD comp2_52 (
    .a(i2[52]),
    .b(sum_1[52]),
    .c(cout_2[51]),
    .cout(cout_2[52]),
    .sum(sum_2[52]));
  AL_FADD comp2_53 (
    .a(i2[53]),
    .b(sum_1[53]),
    .c(cout_2[52]),
    .cout(cout_2[53]),
    .sum(sum_2[53]));
  AL_FADD comp2_54 (
    .a(i2[54]),
    .b(sum_1[54]),
    .c(cout_2[53]),
    .cout(cout_2[54]),
    .sum(sum_2[54]));
  AL_FADD comp2_55 (
    .a(i2[55]),
    .b(sum_1[55]),
    .c(cout_2[54]),
    .cout(cout_2[55]),
    .sum(sum_2[55]));
  AL_FADD comp2_56 (
    .a(i2[56]),
    .b(sum_1[56]),
    .c(cout_2[55]),
    .cout(cout_2[56]),
    .sum(sum_2[56]));
  AL_FADD comp2_57 (
    .a(i2[57]),
    .b(sum_1[57]),
    .c(cout_2[56]),
    .cout(cout_2[57]),
    .sum(sum_2[57]));
  AL_FADD comp2_58 (
    .a(i2[58]),
    .b(sum_1[58]),
    .c(cout_2[57]),
    .cout(cout_2[58]),
    .sum(sum_2[58]));
  AL_FADD comp2_59 (
    .a(i2[59]),
    .b(sum_1[59]),
    .c(cout_2[58]),
    .cout(cout_2[59]),
    .sum(sum_2[59]));
  AL_FADD comp2_6 (
    .a(i2[6]),
    .b(sum_1[6]),
    .c(cout_2[5]),
    .cout(cout_2[6]),
    .sum(sum_2[6]));
  AL_FADD comp2_60 (
    .a(i2[60]),
    .b(sum_1[60]),
    .c(cout_2[59]),
    .cout(cout_2[60]),
    .sum(sum_2[60]));
  AL_FADD comp2_61 (
    .a(1'b0),
    .b(sum_1[61]),
    .c(cout_2[60]),
    .cout(cout_2[61]),
    .sum(sum_2[61]));
  AL_FADD comp2_62 (
    .a(1'b0),
    .b(sum_1[62]),
    .c(cout_2[61]),
    .cout(cout_2[62]),
    .sum(sum_2[62]));
  AL_FADD comp2_63 (
    .a(1'b0),
    .b(cout_1[62]),
    .c(cout_2[62]),
    .cout(cout_2[63]),
    .sum(sum_2[63]));
  AL_FADD comp2_7 (
    .a(i2[7]),
    .b(sum_1[7]),
    .c(cout_2[6]),
    .cout(cout_2[7]),
    .sum(sum_2[7]));
  AL_FADD comp2_8 (
    .a(i2[8]),
    .b(sum_1[8]),
    .c(cout_2[7]),
    .cout(cout_2[8]),
    .sum(sum_2[8]));
  AL_FADD comp2_9 (
    .a(i2[9]),
    .b(sum_1[9]),
    .c(cout_2[8]),
    .cout(cout_2[9]),
    .sum(sum_2[9]));
  AL_FADD comp30_0 (
    .a(i30[0]),
    .b(sum_29[0]),
    .c(1'b0),
    .cout(cout_30[0]),
    .sum(sum_30[0]));
  AL_FADD comp30_1 (
    .a(i30[1]),
    .b(sum_29[1]),
    .c(cout_30[0]),
    .cout(cout_30[1]),
    .sum(sum_30[1]));
  AL_FADD comp30_10 (
    .a(i30[10]),
    .b(sum_29[10]),
    .c(cout_30[9]),
    .cout(cout_30[10]),
    .sum(sum_30[10]));
  AL_FADD comp30_11 (
    .a(i30[11]),
    .b(sum_29[11]),
    .c(cout_30[10]),
    .cout(cout_30[11]),
    .sum(sum_30[11]));
  AL_FADD comp30_12 (
    .a(i30[12]),
    .b(sum_29[12]),
    .c(cout_30[11]),
    .cout(cout_30[12]),
    .sum(sum_30[12]));
  AL_FADD comp30_13 (
    .a(i30[13]),
    .b(sum_29[13]),
    .c(cout_30[12]),
    .cout(cout_30[13]),
    .sum(sum_30[13]));
  AL_FADD comp30_14 (
    .a(i30[14]),
    .b(sum_29[14]),
    .c(cout_30[13]),
    .cout(cout_30[14]),
    .sum(sum_30[14]));
  AL_FADD comp30_15 (
    .a(i30[15]),
    .b(sum_29[15]),
    .c(cout_30[14]),
    .cout(cout_30[15]),
    .sum(sum_30[15]));
  AL_FADD comp30_16 (
    .a(i30[16]),
    .b(sum_29[16]),
    .c(cout_30[15]),
    .cout(cout_30[16]),
    .sum(sum_30[16]));
  AL_FADD comp30_17 (
    .a(i30[17]),
    .b(sum_29[17]),
    .c(cout_30[16]),
    .cout(cout_30[17]),
    .sum(sum_30[17]));
  AL_FADD comp30_18 (
    .a(i30[18]),
    .b(sum_29[18]),
    .c(cout_30[17]),
    .cout(cout_30[18]),
    .sum(sum_30[18]));
  AL_FADD comp30_19 (
    .a(i30[19]),
    .b(sum_29[19]),
    .c(cout_30[18]),
    .cout(cout_30[19]),
    .sum(sum_30[19]));
  AL_FADD comp30_2 (
    .a(i30[2]),
    .b(sum_29[2]),
    .c(cout_30[1]),
    .cout(cout_30[2]),
    .sum(sum_30[2]));
  AL_FADD comp30_20 (
    .a(i30[20]),
    .b(sum_29[20]),
    .c(cout_30[19]),
    .cout(cout_30[20]),
    .sum(sum_30[20]));
  AL_FADD comp30_21 (
    .a(i30[21]),
    .b(sum_29[21]),
    .c(cout_30[20]),
    .cout(cout_30[21]),
    .sum(sum_30[21]));
  AL_FADD comp30_22 (
    .a(i30[22]),
    .b(sum_29[22]),
    .c(cout_30[21]),
    .cout(cout_30[22]),
    .sum(sum_30[22]));
  AL_FADD comp30_23 (
    .a(i30[23]),
    .b(sum_29[23]),
    .c(cout_30[22]),
    .cout(cout_30[23]),
    .sum(sum_30[23]));
  AL_FADD comp30_24 (
    .a(i30[24]),
    .b(sum_29[24]),
    .c(cout_30[23]),
    .cout(cout_30[24]),
    .sum(sum_30[24]));
  AL_FADD comp30_25 (
    .a(i30[25]),
    .b(sum_29[25]),
    .c(cout_30[24]),
    .cout(cout_30[25]),
    .sum(sum_30[25]));
  AL_FADD comp30_26 (
    .a(i30[26]),
    .b(sum_29[26]),
    .c(cout_30[25]),
    .cout(cout_30[26]),
    .sum(sum_30[26]));
  AL_FADD comp30_27 (
    .a(i30[27]),
    .b(sum_29[27]),
    .c(cout_30[26]),
    .cout(cout_30[27]),
    .sum(sum_30[27]));
  AL_FADD comp30_28 (
    .a(i30[28]),
    .b(sum_29[28]),
    .c(cout_30[27]),
    .cout(cout_30[28]),
    .sum(sum_30[28]));
  AL_FADD comp30_29 (
    .a(i30[29]),
    .b(sum_29[29]),
    .c(cout_30[28]),
    .cout(cout_30[29]),
    .sum(sum_30[29]));
  AL_FADD comp30_3 (
    .a(i30[3]),
    .b(sum_29[3]),
    .c(cout_30[2]),
    .cout(cout_30[3]),
    .sum(sum_30[3]));
  AL_FADD comp30_30 (
    .a(i30[30]),
    .b(sum_29[30]),
    .c(cout_30[29]),
    .cout(cout_30[30]),
    .sum(sum_30[30]));
  AL_FADD comp30_31 (
    .a(i30[31]),
    .b(sum_29[31]),
    .c(cout_30[30]),
    .cout(cout_30[31]),
    .sum(sum_30[31]));
  AL_FADD comp30_32 (
    .a(i30[32]),
    .b(sum_29[32]),
    .c(cout_30[31]),
    .cout(cout_30[32]),
    .sum(sum_30[32]));
  AL_FADD comp30_33 (
    .a(1'b0),
    .b(sum_29[33]),
    .c(cout_30[32]),
    .cout(cout_30[33]),
    .sum(sum_30[33]));
  AL_FADD comp30_34 (
    .a(1'b0),
    .b(sum_29[34]),
    .c(cout_30[33]),
    .cout(cout_30[34]),
    .sum(sum_30[34]));
  AL_FADD comp30_35 (
    .a(1'b0),
    .b(sum_29[35]),
    .c(cout_30[34]),
    .cout(cout_30[35]),
    .sum(sum_30[35]));
  AL_FADD comp30_36 (
    .a(1'b0),
    .b(sum_29[36]),
    .c(cout_30[35]),
    .cout(cout_30[36]),
    .sum(sum_30[36]));
  AL_FADD comp30_37 (
    .a(1'b0),
    .b(sum_29[37]),
    .c(cout_30[36]),
    .cout(cout_30[37]),
    .sum(sum_30[37]));
  AL_FADD comp30_38 (
    .a(1'b0),
    .b(sum_29[38]),
    .c(cout_30[37]),
    .cout(cout_30[38]),
    .sum(sum_30[38]));
  AL_FADD comp30_39 (
    .a(1'b0),
    .b(sum_29[39]),
    .c(cout_30[38]),
    .cout(cout_30[39]),
    .sum(sum_30[39]));
  AL_FADD comp30_4 (
    .a(i30[4]),
    .b(sum_29[4]),
    .c(cout_30[3]),
    .cout(cout_30[4]),
    .sum(sum_30[4]));
  AL_FADD comp30_40 (
    .a(1'b0),
    .b(sum_29[40]),
    .c(cout_30[39]),
    .cout(cout_30[40]),
    .sum(sum_30[40]));
  AL_FADD comp30_41 (
    .a(1'b0),
    .b(sum_29[41]),
    .c(cout_30[40]),
    .cout(cout_30[41]),
    .sum(sum_30[41]));
  AL_FADD comp30_42 (
    .a(1'b0),
    .b(sum_29[42]),
    .c(cout_30[41]),
    .cout(cout_30[42]),
    .sum(sum_30[42]));
  AL_FADD comp30_43 (
    .a(1'b0),
    .b(sum_29[43]),
    .c(cout_30[42]),
    .cout(cout_30[43]),
    .sum(sum_30[43]));
  AL_FADD comp30_44 (
    .a(1'b0),
    .b(sum_29[44]),
    .c(cout_30[43]),
    .cout(cout_30[44]),
    .sum(sum_30[44]));
  AL_FADD comp30_45 (
    .a(1'b0),
    .b(sum_29[45]),
    .c(cout_30[44]),
    .cout(cout_30[45]),
    .sum(sum_30[45]));
  AL_FADD comp30_46 (
    .a(1'b0),
    .b(sum_29[46]),
    .c(cout_30[45]),
    .cout(cout_30[46]),
    .sum(sum_30[46]));
  AL_FADD comp30_47 (
    .a(1'b0),
    .b(sum_29[47]),
    .c(cout_30[46]),
    .cout(cout_30[47]),
    .sum(sum_30[47]));
  AL_FADD comp30_48 (
    .a(1'b0),
    .b(sum_29[48]),
    .c(cout_30[47]),
    .cout(cout_30[48]),
    .sum(sum_30[48]));
  AL_FADD comp30_49 (
    .a(1'b0),
    .b(sum_29[49]),
    .c(cout_30[48]),
    .cout(cout_30[49]),
    .sum(sum_30[49]));
  AL_FADD comp30_5 (
    .a(i30[5]),
    .b(sum_29[5]),
    .c(cout_30[4]),
    .cout(cout_30[5]),
    .sum(sum_30[5]));
  AL_FADD comp30_50 (
    .a(1'b0),
    .b(sum_29[50]),
    .c(cout_30[49]),
    .cout(cout_30[50]),
    .sum(sum_30[50]));
  AL_FADD comp30_51 (
    .a(1'b0),
    .b(sum_29[51]),
    .c(cout_30[50]),
    .cout(cout_30[51]),
    .sum(sum_30[51]));
  AL_FADD comp30_52 (
    .a(1'b0),
    .b(sum_29[52]),
    .c(cout_30[51]),
    .cout(cout_30[52]),
    .sum(sum_30[52]));
  AL_FADD comp30_53 (
    .a(1'b0),
    .b(sum_29[53]),
    .c(cout_30[52]),
    .cout(cout_30[53]),
    .sum(sum_30[53]));
  AL_FADD comp30_54 (
    .a(1'b0),
    .b(sum_29[54]),
    .c(cout_30[53]),
    .cout(cout_30[54]),
    .sum(sum_30[54]));
  AL_FADD comp30_55 (
    .a(1'b0),
    .b(sum_29[55]),
    .c(cout_30[54]),
    .cout(cout_30[55]),
    .sum(sum_30[55]));
  AL_FADD comp30_56 (
    .a(1'b0),
    .b(sum_29[56]),
    .c(cout_30[55]),
    .cout(cout_30[56]),
    .sum(sum_30[56]));
  AL_FADD comp30_57 (
    .a(1'b0),
    .b(sum_29[57]),
    .c(cout_30[56]),
    .cout(cout_30[57]),
    .sum(sum_30[57]));
  AL_FADD comp30_58 (
    .a(1'b0),
    .b(sum_29[58]),
    .c(cout_30[57]),
    .cout(cout_30[58]),
    .sum(sum_30[58]));
  AL_FADD comp30_59 (
    .a(1'b0),
    .b(sum_29[59]),
    .c(cout_30[58]),
    .cout(cout_30[59]),
    .sum(sum_30[59]));
  AL_FADD comp30_6 (
    .a(i30[6]),
    .b(sum_29[6]),
    .c(cout_30[5]),
    .cout(cout_30[6]),
    .sum(sum_30[6]));
  AL_FADD comp30_60 (
    .a(1'b0),
    .b(sum_29[60]),
    .c(cout_30[59]),
    .cout(cout_30[60]),
    .sum(sum_30[60]));
  AL_FADD comp30_61 (
    .a(1'b0),
    .b(sum_29[61]),
    .c(cout_30[60]),
    .cout(cout_30[61]),
    .sum(sum_30[61]));
  AL_FADD comp30_62 (
    .a(1'b0),
    .b(sum_29[62]),
    .c(cout_30[61]),
    .cout(cout_30[62]),
    .sum(sum_30[62]));
  AL_FADD comp30_63 (
    .a(1'b0),
    .b(sum_29[63]),
    .c(cout_30[62]),
    .cout(cout_30[63]),
    .sum(sum_30[63]));
  AL_FADD comp30_7 (
    .a(i30[7]),
    .b(sum_29[7]),
    .c(cout_30[6]),
    .cout(cout_30[7]),
    .sum(sum_30[7]));
  AL_FADD comp30_8 (
    .a(i30[8]),
    .b(sum_29[8]),
    .c(cout_30[7]),
    .cout(cout_30[8]),
    .sum(sum_30[8]));
  AL_FADD comp30_9 (
    .a(i30[9]),
    .b(sum_29[9]),
    .c(cout_30[8]),
    .cout(cout_30[9]),
    .sum(sum_30[9]));
  AL_FADD comp31_0 (
    .a(i31[0]),
    .b(sum_30[0]),
    .c(1'b0),
    .cout(cout_31[0]),
    .sum(sum_31[0]));
  AL_FADD comp31_1 (
    .a(i31[1]),
    .b(sum_30[1]),
    .c(cout_31[0]),
    .cout(cout_31[1]),
    .sum(sum_31[1]));
  AL_FADD comp31_10 (
    .a(i31[10]),
    .b(sum_30[10]),
    .c(cout_31[9]),
    .cout(cout_31[10]),
    .sum(sum_31[10]));
  AL_FADD comp31_11 (
    .a(i31[11]),
    .b(sum_30[11]),
    .c(cout_31[10]),
    .cout(cout_31[11]),
    .sum(sum_31[11]));
  AL_FADD comp31_12 (
    .a(i31[12]),
    .b(sum_30[12]),
    .c(cout_31[11]),
    .cout(cout_31[12]),
    .sum(sum_31[12]));
  AL_FADD comp31_13 (
    .a(i31[13]),
    .b(sum_30[13]),
    .c(cout_31[12]),
    .cout(cout_31[13]),
    .sum(sum_31[13]));
  AL_FADD comp31_14 (
    .a(i31[14]),
    .b(sum_30[14]),
    .c(cout_31[13]),
    .cout(cout_31[14]),
    .sum(sum_31[14]));
  AL_FADD comp31_15 (
    .a(i31[15]),
    .b(sum_30[15]),
    .c(cout_31[14]),
    .cout(cout_31[15]),
    .sum(sum_31[15]));
  AL_FADD comp31_16 (
    .a(i31[16]),
    .b(sum_30[16]),
    .c(cout_31[15]),
    .cout(cout_31[16]),
    .sum(sum_31[16]));
  AL_FADD comp31_17 (
    .a(i31[17]),
    .b(sum_30[17]),
    .c(cout_31[16]),
    .cout(cout_31[17]),
    .sum(sum_31[17]));
  AL_FADD comp31_18 (
    .a(i31[18]),
    .b(sum_30[18]),
    .c(cout_31[17]),
    .cout(cout_31[18]),
    .sum(sum_31[18]));
  AL_FADD comp31_19 (
    .a(i31[19]),
    .b(sum_30[19]),
    .c(cout_31[18]),
    .cout(cout_31[19]),
    .sum(sum_31[19]));
  AL_FADD comp31_2 (
    .a(i31[2]),
    .b(sum_30[2]),
    .c(cout_31[1]),
    .cout(cout_31[2]),
    .sum(sum_31[2]));
  AL_FADD comp31_20 (
    .a(i31[20]),
    .b(sum_30[20]),
    .c(cout_31[19]),
    .cout(cout_31[20]),
    .sum(sum_31[20]));
  AL_FADD comp31_21 (
    .a(i31[21]),
    .b(sum_30[21]),
    .c(cout_31[20]),
    .cout(cout_31[21]),
    .sum(sum_31[21]));
  AL_FADD comp31_22 (
    .a(i31[22]),
    .b(sum_30[22]),
    .c(cout_31[21]),
    .cout(cout_31[22]),
    .sum(sum_31[22]));
  AL_FADD comp31_23 (
    .a(i31[23]),
    .b(sum_30[23]),
    .c(cout_31[22]),
    .cout(cout_31[23]),
    .sum(sum_31[23]));
  AL_FADD comp31_24 (
    .a(i31[24]),
    .b(sum_30[24]),
    .c(cout_31[23]),
    .cout(cout_31[24]),
    .sum(sum_31[24]));
  AL_FADD comp31_25 (
    .a(i31[25]),
    .b(sum_30[25]),
    .c(cout_31[24]),
    .cout(cout_31[25]),
    .sum(sum_31[25]));
  AL_FADD comp31_26 (
    .a(i31[26]),
    .b(sum_30[26]),
    .c(cout_31[25]),
    .cout(cout_31[26]),
    .sum(sum_31[26]));
  AL_FADD comp31_27 (
    .a(i31[27]),
    .b(sum_30[27]),
    .c(cout_31[26]),
    .cout(cout_31[27]),
    .sum(sum_31[27]));
  AL_FADD comp31_28 (
    .a(i31[28]),
    .b(sum_30[28]),
    .c(cout_31[27]),
    .cout(cout_31[28]),
    .sum(sum_31[28]));
  AL_FADD comp31_29 (
    .a(i31[29]),
    .b(sum_30[29]),
    .c(cout_31[28]),
    .cout(cout_31[29]),
    .sum(sum_31[29]));
  AL_FADD comp31_3 (
    .a(i31[3]),
    .b(sum_30[3]),
    .c(cout_31[2]),
    .cout(cout_31[3]),
    .sum(sum_31[3]));
  AL_FADD comp31_30 (
    .a(i31[30]),
    .b(sum_30[30]),
    .c(cout_31[29]),
    .cout(cout_31[30]),
    .sum(sum_31[30]));
  AL_FADD comp31_31 (
    .a(i31[31]),
    .b(sum_30[31]),
    .c(cout_31[30]),
    .cout(cout_31[31]),
    .sum(sum_31[31]));
  AL_FADD comp31_32 (
    .a(1'b0),
    .b(sum_30[32]),
    .c(cout_31[31]),
    .cout(cout_31[32]),
    .sum(sum_31[32]));
  AL_FADD comp31_33 (
    .a(1'b0),
    .b(sum_30[33]),
    .c(cout_31[32]),
    .cout(cout_31[33]),
    .sum(sum_31[33]));
  AL_FADD comp31_34 (
    .a(1'b0),
    .b(sum_30[34]),
    .c(cout_31[33]),
    .cout(cout_31[34]),
    .sum(sum_31[34]));
  AL_FADD comp31_35 (
    .a(1'b0),
    .b(sum_30[35]),
    .c(cout_31[34]),
    .cout(cout_31[35]),
    .sum(sum_31[35]));
  AL_FADD comp31_36 (
    .a(1'b0),
    .b(sum_30[36]),
    .c(cout_31[35]),
    .cout(cout_31[36]),
    .sum(sum_31[36]));
  AL_FADD comp31_37 (
    .a(1'b0),
    .b(sum_30[37]),
    .c(cout_31[36]),
    .cout(cout_31[37]),
    .sum(sum_31[37]));
  AL_FADD comp31_38 (
    .a(1'b0),
    .b(sum_30[38]),
    .c(cout_31[37]),
    .cout(cout_31[38]),
    .sum(sum_31[38]));
  AL_FADD comp31_39 (
    .a(1'b0),
    .b(sum_30[39]),
    .c(cout_31[38]),
    .cout(cout_31[39]),
    .sum(sum_31[39]));
  AL_FADD comp31_4 (
    .a(i31[4]),
    .b(sum_30[4]),
    .c(cout_31[3]),
    .cout(cout_31[4]),
    .sum(sum_31[4]));
  AL_FADD comp31_40 (
    .a(1'b0),
    .b(sum_30[40]),
    .c(cout_31[39]),
    .cout(cout_31[40]),
    .sum(sum_31[40]));
  AL_FADD comp31_41 (
    .a(1'b0),
    .b(sum_30[41]),
    .c(cout_31[40]),
    .cout(cout_31[41]),
    .sum(sum_31[41]));
  AL_FADD comp31_42 (
    .a(1'b0),
    .b(sum_30[42]),
    .c(cout_31[41]),
    .cout(cout_31[42]),
    .sum(sum_31[42]));
  AL_FADD comp31_43 (
    .a(1'b0),
    .b(sum_30[43]),
    .c(cout_31[42]),
    .cout(cout_31[43]),
    .sum(sum_31[43]));
  AL_FADD comp31_44 (
    .a(1'b0),
    .b(sum_30[44]),
    .c(cout_31[43]),
    .cout(cout_31[44]),
    .sum(sum_31[44]));
  AL_FADD comp31_45 (
    .a(1'b0),
    .b(sum_30[45]),
    .c(cout_31[44]),
    .cout(cout_31[45]),
    .sum(sum_31[45]));
  AL_FADD comp31_46 (
    .a(1'b0),
    .b(sum_30[46]),
    .c(cout_31[45]),
    .cout(cout_31[46]),
    .sum(sum_31[46]));
  AL_FADD comp31_47 (
    .a(1'b0),
    .b(sum_30[47]),
    .c(cout_31[46]),
    .cout(cout_31[47]),
    .sum(sum_31[47]));
  AL_FADD comp31_48 (
    .a(1'b0),
    .b(sum_30[48]),
    .c(cout_31[47]),
    .cout(cout_31[48]),
    .sum(sum_31[48]));
  AL_FADD comp31_49 (
    .a(1'b0),
    .b(sum_30[49]),
    .c(cout_31[48]),
    .cout(cout_31[49]),
    .sum(sum_31[49]));
  AL_FADD comp31_5 (
    .a(i31[5]),
    .b(sum_30[5]),
    .c(cout_31[4]),
    .cout(cout_31[5]),
    .sum(sum_31[5]));
  AL_FADD comp31_50 (
    .a(1'b0),
    .b(sum_30[50]),
    .c(cout_31[49]),
    .cout(cout_31[50]),
    .sum(sum_31[50]));
  AL_FADD comp31_51 (
    .a(1'b0),
    .b(sum_30[51]),
    .c(cout_31[50]),
    .cout(cout_31[51]),
    .sum(sum_31[51]));
  AL_FADD comp31_52 (
    .a(1'b0),
    .b(sum_30[52]),
    .c(cout_31[51]),
    .cout(cout_31[52]),
    .sum(sum_31[52]));
  AL_FADD comp31_53 (
    .a(1'b0),
    .b(sum_30[53]),
    .c(cout_31[52]),
    .cout(cout_31[53]),
    .sum(sum_31[53]));
  AL_FADD comp31_54 (
    .a(1'b0),
    .b(sum_30[54]),
    .c(cout_31[53]),
    .cout(cout_31[54]),
    .sum(sum_31[54]));
  AL_FADD comp31_55 (
    .a(1'b0),
    .b(sum_30[55]),
    .c(cout_31[54]),
    .cout(cout_31[55]),
    .sum(sum_31[55]));
  AL_FADD comp31_56 (
    .a(1'b0),
    .b(sum_30[56]),
    .c(cout_31[55]),
    .cout(cout_31[56]),
    .sum(sum_31[56]));
  AL_FADD comp31_57 (
    .a(1'b0),
    .b(sum_30[57]),
    .c(cout_31[56]),
    .cout(cout_31[57]),
    .sum(sum_31[57]));
  AL_FADD comp31_58 (
    .a(1'b0),
    .b(sum_30[58]),
    .c(cout_31[57]),
    .cout(cout_31[58]),
    .sum(sum_31[58]));
  AL_FADD comp31_59 (
    .a(1'b0),
    .b(sum_30[59]),
    .c(cout_31[58]),
    .cout(cout_31[59]),
    .sum(sum_31[59]));
  AL_FADD comp31_6 (
    .a(i31[6]),
    .b(sum_30[6]),
    .c(cout_31[5]),
    .cout(cout_31[6]),
    .sum(sum_31[6]));
  AL_FADD comp31_60 (
    .a(1'b0),
    .b(sum_30[60]),
    .c(cout_31[59]),
    .cout(cout_31[60]),
    .sum(sum_31[60]));
  AL_FADD comp31_61 (
    .a(1'b0),
    .b(sum_30[61]),
    .c(cout_31[60]),
    .cout(cout_31[61]),
    .sum(sum_31[61]));
  AL_FADD comp31_62 (
    .a(1'b0),
    .b(sum_30[62]),
    .c(cout_31[61]),
    .cout(cout_31[62]),
    .sum(sum_31[62]));
  AL_FADD comp31_63 (
    .a(1'b0),
    .b(sum_30[63]),
    .c(cout_31[62]),
    .cout(cout_31[63]),
    .sum(sum_31[63]));
  AL_FADD comp31_7 (
    .a(i31[7]),
    .b(sum_30[7]),
    .c(cout_31[6]),
    .cout(cout_31[7]),
    .sum(sum_31[7]));
  AL_FADD comp31_8 (
    .a(i31[8]),
    .b(sum_30[8]),
    .c(cout_31[7]),
    .cout(cout_31[8]),
    .sum(sum_31[8]));
  AL_FADD comp31_9 (
    .a(i31[9]),
    .b(sum_30[9]),
    .c(cout_31[8]),
    .cout(cout_31[9]),
    .sum(sum_31[9]));
  AL_FADD comp3_0 (
    .a(i3[0]),
    .b(sum_2[0]),
    .c(1'b0),
    .cout(cout_3[0]),
    .sum(sum_3[0]));
  AL_FADD comp3_1 (
    .a(i3[1]),
    .b(sum_2[1]),
    .c(cout_3[0]),
    .cout(cout_3[1]),
    .sum(sum_3[1]));
  AL_FADD comp3_10 (
    .a(i3[10]),
    .b(sum_2[10]),
    .c(cout_3[9]),
    .cout(cout_3[10]),
    .sum(sum_3[10]));
  AL_FADD comp3_11 (
    .a(i3[11]),
    .b(sum_2[11]),
    .c(cout_3[10]),
    .cout(cout_3[11]),
    .sum(sum_3[11]));
  AL_FADD comp3_12 (
    .a(i3[12]),
    .b(sum_2[12]),
    .c(cout_3[11]),
    .cout(cout_3[12]),
    .sum(sum_3[12]));
  AL_FADD comp3_13 (
    .a(i3[13]),
    .b(sum_2[13]),
    .c(cout_3[12]),
    .cout(cout_3[13]),
    .sum(sum_3[13]));
  AL_FADD comp3_14 (
    .a(i3[14]),
    .b(sum_2[14]),
    .c(cout_3[13]),
    .cout(cout_3[14]),
    .sum(sum_3[14]));
  AL_FADD comp3_15 (
    .a(i3[15]),
    .b(sum_2[15]),
    .c(cout_3[14]),
    .cout(cout_3[15]),
    .sum(sum_3[15]));
  AL_FADD comp3_16 (
    .a(i3[16]),
    .b(sum_2[16]),
    .c(cout_3[15]),
    .cout(cout_3[16]),
    .sum(sum_3[16]));
  AL_FADD comp3_17 (
    .a(i3[17]),
    .b(sum_2[17]),
    .c(cout_3[16]),
    .cout(cout_3[17]),
    .sum(sum_3[17]));
  AL_FADD comp3_18 (
    .a(i3[18]),
    .b(sum_2[18]),
    .c(cout_3[17]),
    .cout(cout_3[18]),
    .sum(sum_3[18]));
  AL_FADD comp3_19 (
    .a(i3[19]),
    .b(sum_2[19]),
    .c(cout_3[18]),
    .cout(cout_3[19]),
    .sum(sum_3[19]));
  AL_FADD comp3_2 (
    .a(i3[2]),
    .b(sum_2[2]),
    .c(cout_3[1]),
    .cout(cout_3[2]),
    .sum(sum_3[2]));
  AL_FADD comp3_20 (
    .a(i3[20]),
    .b(sum_2[20]),
    .c(cout_3[19]),
    .cout(cout_3[20]),
    .sum(sum_3[20]));
  AL_FADD comp3_21 (
    .a(i3[21]),
    .b(sum_2[21]),
    .c(cout_3[20]),
    .cout(cout_3[21]),
    .sum(sum_3[21]));
  AL_FADD comp3_22 (
    .a(i3[22]),
    .b(sum_2[22]),
    .c(cout_3[21]),
    .cout(cout_3[22]),
    .sum(sum_3[22]));
  AL_FADD comp3_23 (
    .a(i3[23]),
    .b(sum_2[23]),
    .c(cout_3[22]),
    .cout(cout_3[23]),
    .sum(sum_3[23]));
  AL_FADD comp3_24 (
    .a(i3[24]),
    .b(sum_2[24]),
    .c(cout_3[23]),
    .cout(cout_3[24]),
    .sum(sum_3[24]));
  AL_FADD comp3_25 (
    .a(i3[25]),
    .b(sum_2[25]),
    .c(cout_3[24]),
    .cout(cout_3[25]),
    .sum(sum_3[25]));
  AL_FADD comp3_26 (
    .a(i3[26]),
    .b(sum_2[26]),
    .c(cout_3[25]),
    .cout(cout_3[26]),
    .sum(sum_3[26]));
  AL_FADD comp3_27 (
    .a(i3[27]),
    .b(sum_2[27]),
    .c(cout_3[26]),
    .cout(cout_3[27]),
    .sum(sum_3[27]));
  AL_FADD comp3_28 (
    .a(i3[28]),
    .b(sum_2[28]),
    .c(cout_3[27]),
    .cout(cout_3[28]),
    .sum(sum_3[28]));
  AL_FADD comp3_29 (
    .a(i3[29]),
    .b(sum_2[29]),
    .c(cout_3[28]),
    .cout(cout_3[29]),
    .sum(sum_3[29]));
  AL_FADD comp3_3 (
    .a(i3[3]),
    .b(sum_2[3]),
    .c(cout_3[2]),
    .cout(cout_3[3]),
    .sum(sum_3[3]));
  AL_FADD comp3_30 (
    .a(i3[30]),
    .b(sum_2[30]),
    .c(cout_3[29]),
    .cout(cout_3[30]),
    .sum(sum_3[30]));
  AL_FADD comp3_31 (
    .a(i3[31]),
    .b(sum_2[31]),
    .c(cout_3[30]),
    .cout(cout_3[31]),
    .sum(sum_3[31]));
  AL_FADD comp3_32 (
    .a(i3[32]),
    .b(sum_2[32]),
    .c(cout_3[31]),
    .cout(cout_3[32]),
    .sum(sum_3[32]));
  AL_FADD comp3_33 (
    .a(i3[33]),
    .b(sum_2[33]),
    .c(cout_3[32]),
    .cout(cout_3[33]),
    .sum(sum_3[33]));
  AL_FADD comp3_34 (
    .a(i3[34]),
    .b(sum_2[34]),
    .c(cout_3[33]),
    .cout(cout_3[34]),
    .sum(sum_3[34]));
  AL_FADD comp3_35 (
    .a(i3[35]),
    .b(sum_2[35]),
    .c(cout_3[34]),
    .cout(cout_3[35]),
    .sum(sum_3[35]));
  AL_FADD comp3_36 (
    .a(i3[36]),
    .b(sum_2[36]),
    .c(cout_3[35]),
    .cout(cout_3[36]),
    .sum(sum_3[36]));
  AL_FADD comp3_37 (
    .a(i3[37]),
    .b(sum_2[37]),
    .c(cout_3[36]),
    .cout(cout_3[37]),
    .sum(sum_3[37]));
  AL_FADD comp3_38 (
    .a(i3[38]),
    .b(sum_2[38]),
    .c(cout_3[37]),
    .cout(cout_3[38]),
    .sum(sum_3[38]));
  AL_FADD comp3_39 (
    .a(i3[39]),
    .b(sum_2[39]),
    .c(cout_3[38]),
    .cout(cout_3[39]),
    .sum(sum_3[39]));
  AL_FADD comp3_4 (
    .a(i3[4]),
    .b(sum_2[4]),
    .c(cout_3[3]),
    .cout(cout_3[4]),
    .sum(sum_3[4]));
  AL_FADD comp3_40 (
    .a(i3[40]),
    .b(sum_2[40]),
    .c(cout_3[39]),
    .cout(cout_3[40]),
    .sum(sum_3[40]));
  AL_FADD comp3_41 (
    .a(i3[41]),
    .b(sum_2[41]),
    .c(cout_3[40]),
    .cout(cout_3[41]),
    .sum(sum_3[41]));
  AL_FADD comp3_42 (
    .a(i3[42]),
    .b(sum_2[42]),
    .c(cout_3[41]),
    .cout(cout_3[42]),
    .sum(sum_3[42]));
  AL_FADD comp3_43 (
    .a(i3[43]),
    .b(sum_2[43]),
    .c(cout_3[42]),
    .cout(cout_3[43]),
    .sum(sum_3[43]));
  AL_FADD comp3_44 (
    .a(i3[44]),
    .b(sum_2[44]),
    .c(cout_3[43]),
    .cout(cout_3[44]),
    .sum(sum_3[44]));
  AL_FADD comp3_45 (
    .a(i3[45]),
    .b(sum_2[45]),
    .c(cout_3[44]),
    .cout(cout_3[45]),
    .sum(sum_3[45]));
  AL_FADD comp3_46 (
    .a(i3[46]),
    .b(sum_2[46]),
    .c(cout_3[45]),
    .cout(cout_3[46]),
    .sum(sum_3[46]));
  AL_FADD comp3_47 (
    .a(i3[47]),
    .b(sum_2[47]),
    .c(cout_3[46]),
    .cout(cout_3[47]),
    .sum(sum_3[47]));
  AL_FADD comp3_48 (
    .a(i3[48]),
    .b(sum_2[48]),
    .c(cout_3[47]),
    .cout(cout_3[48]),
    .sum(sum_3[48]));
  AL_FADD comp3_49 (
    .a(i3[49]),
    .b(sum_2[49]),
    .c(cout_3[48]),
    .cout(cout_3[49]),
    .sum(sum_3[49]));
  AL_FADD comp3_5 (
    .a(i3[5]),
    .b(sum_2[5]),
    .c(cout_3[4]),
    .cout(cout_3[5]),
    .sum(sum_3[5]));
  AL_FADD comp3_50 (
    .a(i3[50]),
    .b(sum_2[50]),
    .c(cout_3[49]),
    .cout(cout_3[50]),
    .sum(sum_3[50]));
  AL_FADD comp3_51 (
    .a(i3[51]),
    .b(sum_2[51]),
    .c(cout_3[50]),
    .cout(cout_3[51]),
    .sum(sum_3[51]));
  AL_FADD comp3_52 (
    .a(i3[52]),
    .b(sum_2[52]),
    .c(cout_3[51]),
    .cout(cout_3[52]),
    .sum(sum_3[52]));
  AL_FADD comp3_53 (
    .a(i3[53]),
    .b(sum_2[53]),
    .c(cout_3[52]),
    .cout(cout_3[53]),
    .sum(sum_3[53]));
  AL_FADD comp3_54 (
    .a(i3[54]),
    .b(sum_2[54]),
    .c(cout_3[53]),
    .cout(cout_3[54]),
    .sum(sum_3[54]));
  AL_FADD comp3_55 (
    .a(i3[55]),
    .b(sum_2[55]),
    .c(cout_3[54]),
    .cout(cout_3[55]),
    .sum(sum_3[55]));
  AL_FADD comp3_56 (
    .a(i3[56]),
    .b(sum_2[56]),
    .c(cout_3[55]),
    .cout(cout_3[56]),
    .sum(sum_3[56]));
  AL_FADD comp3_57 (
    .a(i3[57]),
    .b(sum_2[57]),
    .c(cout_3[56]),
    .cout(cout_3[57]),
    .sum(sum_3[57]));
  AL_FADD comp3_58 (
    .a(i3[58]),
    .b(sum_2[58]),
    .c(cout_3[57]),
    .cout(cout_3[58]),
    .sum(sum_3[58]));
  AL_FADD comp3_59 (
    .a(i3[59]),
    .b(sum_2[59]),
    .c(cout_3[58]),
    .cout(cout_3[59]),
    .sum(sum_3[59]));
  AL_FADD comp3_6 (
    .a(i3[6]),
    .b(sum_2[6]),
    .c(cout_3[5]),
    .cout(cout_3[6]),
    .sum(sum_3[6]));
  AL_FADD comp3_60 (
    .a(1'b0),
    .b(sum_2[60]),
    .c(cout_3[59]),
    .cout(cout_3[60]),
    .sum(sum_3[60]));
  AL_FADD comp3_61 (
    .a(1'b0),
    .b(sum_2[61]),
    .c(cout_3[60]),
    .cout(cout_3[61]),
    .sum(sum_3[61]));
  AL_FADD comp3_62 (
    .a(1'b0),
    .b(sum_2[62]),
    .c(cout_3[61]),
    .cout(cout_3[62]),
    .sum(sum_3[62]));
  AL_FADD comp3_63 (
    .a(1'b0),
    .b(sum_2[63]),
    .c(cout_3[62]),
    .cout(cout_3[63]),
    .sum(sum_3[63]));
  AL_FADD comp3_7 (
    .a(i3[7]),
    .b(sum_2[7]),
    .c(cout_3[6]),
    .cout(cout_3[7]),
    .sum(sum_3[7]));
  AL_FADD comp3_8 (
    .a(i3[8]),
    .b(sum_2[8]),
    .c(cout_3[7]),
    .cout(cout_3[8]),
    .sum(sum_3[8]));
  AL_FADD comp3_9 (
    .a(i3[9]),
    .b(sum_2[9]),
    .c(cout_3[8]),
    .cout(cout_3[9]),
    .sum(sum_3[9]));
  AL_FADD comp4_0 (
    .a(i4[0]),
    .b(sum_3[0]),
    .c(1'b0),
    .cout(cout_4[0]),
    .sum(sum_4[0]));
  AL_FADD comp4_1 (
    .a(i4[1]),
    .b(sum_3[1]),
    .c(cout_4[0]),
    .cout(cout_4[1]),
    .sum(sum_4[1]));
  AL_FADD comp4_10 (
    .a(i4[10]),
    .b(sum_3[10]),
    .c(cout_4[9]),
    .cout(cout_4[10]),
    .sum(sum_4[10]));
  AL_FADD comp4_11 (
    .a(i4[11]),
    .b(sum_3[11]),
    .c(cout_4[10]),
    .cout(cout_4[11]),
    .sum(sum_4[11]));
  AL_FADD comp4_12 (
    .a(i4[12]),
    .b(sum_3[12]),
    .c(cout_4[11]),
    .cout(cout_4[12]),
    .sum(sum_4[12]));
  AL_FADD comp4_13 (
    .a(i4[13]),
    .b(sum_3[13]),
    .c(cout_4[12]),
    .cout(cout_4[13]),
    .sum(sum_4[13]));
  AL_FADD comp4_14 (
    .a(i4[14]),
    .b(sum_3[14]),
    .c(cout_4[13]),
    .cout(cout_4[14]),
    .sum(sum_4[14]));
  AL_FADD comp4_15 (
    .a(i4[15]),
    .b(sum_3[15]),
    .c(cout_4[14]),
    .cout(cout_4[15]),
    .sum(sum_4[15]));
  AL_FADD comp4_16 (
    .a(i4[16]),
    .b(sum_3[16]),
    .c(cout_4[15]),
    .cout(cout_4[16]),
    .sum(sum_4[16]));
  AL_FADD comp4_17 (
    .a(i4[17]),
    .b(sum_3[17]),
    .c(cout_4[16]),
    .cout(cout_4[17]),
    .sum(sum_4[17]));
  AL_FADD comp4_18 (
    .a(i4[18]),
    .b(sum_3[18]),
    .c(cout_4[17]),
    .cout(cout_4[18]),
    .sum(sum_4[18]));
  AL_FADD comp4_19 (
    .a(i4[19]),
    .b(sum_3[19]),
    .c(cout_4[18]),
    .cout(cout_4[19]),
    .sum(sum_4[19]));
  AL_FADD comp4_2 (
    .a(i4[2]),
    .b(sum_3[2]),
    .c(cout_4[1]),
    .cout(cout_4[2]),
    .sum(sum_4[2]));
  AL_FADD comp4_20 (
    .a(i4[20]),
    .b(sum_3[20]),
    .c(cout_4[19]),
    .cout(cout_4[20]),
    .sum(sum_4[20]));
  AL_FADD comp4_21 (
    .a(i4[21]),
    .b(sum_3[21]),
    .c(cout_4[20]),
    .cout(cout_4[21]),
    .sum(sum_4[21]));
  AL_FADD comp4_22 (
    .a(i4[22]),
    .b(sum_3[22]),
    .c(cout_4[21]),
    .cout(cout_4[22]),
    .sum(sum_4[22]));
  AL_FADD comp4_23 (
    .a(i4[23]),
    .b(sum_3[23]),
    .c(cout_4[22]),
    .cout(cout_4[23]),
    .sum(sum_4[23]));
  AL_FADD comp4_24 (
    .a(i4[24]),
    .b(sum_3[24]),
    .c(cout_4[23]),
    .cout(cout_4[24]),
    .sum(sum_4[24]));
  AL_FADD comp4_25 (
    .a(i4[25]),
    .b(sum_3[25]),
    .c(cout_4[24]),
    .cout(cout_4[25]),
    .sum(sum_4[25]));
  AL_FADD comp4_26 (
    .a(i4[26]),
    .b(sum_3[26]),
    .c(cout_4[25]),
    .cout(cout_4[26]),
    .sum(sum_4[26]));
  AL_FADD comp4_27 (
    .a(i4[27]),
    .b(sum_3[27]),
    .c(cout_4[26]),
    .cout(cout_4[27]),
    .sum(sum_4[27]));
  AL_FADD comp4_28 (
    .a(i4[28]),
    .b(sum_3[28]),
    .c(cout_4[27]),
    .cout(cout_4[28]),
    .sum(sum_4[28]));
  AL_FADD comp4_29 (
    .a(i4[29]),
    .b(sum_3[29]),
    .c(cout_4[28]),
    .cout(cout_4[29]),
    .sum(sum_4[29]));
  AL_FADD comp4_3 (
    .a(i4[3]),
    .b(sum_3[3]),
    .c(cout_4[2]),
    .cout(cout_4[3]),
    .sum(sum_4[3]));
  AL_FADD comp4_30 (
    .a(i4[30]),
    .b(sum_3[30]),
    .c(cout_4[29]),
    .cout(cout_4[30]),
    .sum(sum_4[30]));
  AL_FADD comp4_31 (
    .a(i4[31]),
    .b(sum_3[31]),
    .c(cout_4[30]),
    .cout(cout_4[31]),
    .sum(sum_4[31]));
  AL_FADD comp4_32 (
    .a(i4[32]),
    .b(sum_3[32]),
    .c(cout_4[31]),
    .cout(cout_4[32]),
    .sum(sum_4[32]));
  AL_FADD comp4_33 (
    .a(i4[33]),
    .b(sum_3[33]),
    .c(cout_4[32]),
    .cout(cout_4[33]),
    .sum(sum_4[33]));
  AL_FADD comp4_34 (
    .a(i4[34]),
    .b(sum_3[34]),
    .c(cout_4[33]),
    .cout(cout_4[34]),
    .sum(sum_4[34]));
  AL_FADD comp4_35 (
    .a(i4[35]),
    .b(sum_3[35]),
    .c(cout_4[34]),
    .cout(cout_4[35]),
    .sum(sum_4[35]));
  AL_FADD comp4_36 (
    .a(i4[36]),
    .b(sum_3[36]),
    .c(cout_4[35]),
    .cout(cout_4[36]),
    .sum(sum_4[36]));
  AL_FADD comp4_37 (
    .a(i4[37]),
    .b(sum_3[37]),
    .c(cout_4[36]),
    .cout(cout_4[37]),
    .sum(sum_4[37]));
  AL_FADD comp4_38 (
    .a(i4[38]),
    .b(sum_3[38]),
    .c(cout_4[37]),
    .cout(cout_4[38]),
    .sum(sum_4[38]));
  AL_FADD comp4_39 (
    .a(i4[39]),
    .b(sum_3[39]),
    .c(cout_4[38]),
    .cout(cout_4[39]),
    .sum(sum_4[39]));
  AL_FADD comp4_4 (
    .a(i4[4]),
    .b(sum_3[4]),
    .c(cout_4[3]),
    .cout(cout_4[4]),
    .sum(sum_4[4]));
  AL_FADD comp4_40 (
    .a(i4[40]),
    .b(sum_3[40]),
    .c(cout_4[39]),
    .cout(cout_4[40]),
    .sum(sum_4[40]));
  AL_FADD comp4_41 (
    .a(i4[41]),
    .b(sum_3[41]),
    .c(cout_4[40]),
    .cout(cout_4[41]),
    .sum(sum_4[41]));
  AL_FADD comp4_42 (
    .a(i4[42]),
    .b(sum_3[42]),
    .c(cout_4[41]),
    .cout(cout_4[42]),
    .sum(sum_4[42]));
  AL_FADD comp4_43 (
    .a(i4[43]),
    .b(sum_3[43]),
    .c(cout_4[42]),
    .cout(cout_4[43]),
    .sum(sum_4[43]));
  AL_FADD comp4_44 (
    .a(i4[44]),
    .b(sum_3[44]),
    .c(cout_4[43]),
    .cout(cout_4[44]),
    .sum(sum_4[44]));
  AL_FADD comp4_45 (
    .a(i4[45]),
    .b(sum_3[45]),
    .c(cout_4[44]),
    .cout(cout_4[45]),
    .sum(sum_4[45]));
  AL_FADD comp4_46 (
    .a(i4[46]),
    .b(sum_3[46]),
    .c(cout_4[45]),
    .cout(cout_4[46]),
    .sum(sum_4[46]));
  AL_FADD comp4_47 (
    .a(i4[47]),
    .b(sum_3[47]),
    .c(cout_4[46]),
    .cout(cout_4[47]),
    .sum(sum_4[47]));
  AL_FADD comp4_48 (
    .a(i4[48]),
    .b(sum_3[48]),
    .c(cout_4[47]),
    .cout(cout_4[48]),
    .sum(sum_4[48]));
  AL_FADD comp4_49 (
    .a(i4[49]),
    .b(sum_3[49]),
    .c(cout_4[48]),
    .cout(cout_4[49]),
    .sum(sum_4[49]));
  AL_FADD comp4_5 (
    .a(i4[5]),
    .b(sum_3[5]),
    .c(cout_4[4]),
    .cout(cout_4[5]),
    .sum(sum_4[5]));
  AL_FADD comp4_50 (
    .a(i4[50]),
    .b(sum_3[50]),
    .c(cout_4[49]),
    .cout(cout_4[50]),
    .sum(sum_4[50]));
  AL_FADD comp4_51 (
    .a(i4[51]),
    .b(sum_3[51]),
    .c(cout_4[50]),
    .cout(cout_4[51]),
    .sum(sum_4[51]));
  AL_FADD comp4_52 (
    .a(i4[52]),
    .b(sum_3[52]),
    .c(cout_4[51]),
    .cout(cout_4[52]),
    .sum(sum_4[52]));
  AL_FADD comp4_53 (
    .a(i4[53]),
    .b(sum_3[53]),
    .c(cout_4[52]),
    .cout(cout_4[53]),
    .sum(sum_4[53]));
  AL_FADD comp4_54 (
    .a(i4[54]),
    .b(sum_3[54]),
    .c(cout_4[53]),
    .cout(cout_4[54]),
    .sum(sum_4[54]));
  AL_FADD comp4_55 (
    .a(i4[55]),
    .b(sum_3[55]),
    .c(cout_4[54]),
    .cout(cout_4[55]),
    .sum(sum_4[55]));
  AL_FADD comp4_56 (
    .a(i4[56]),
    .b(sum_3[56]),
    .c(cout_4[55]),
    .cout(cout_4[56]),
    .sum(sum_4[56]));
  AL_FADD comp4_57 (
    .a(i4[57]),
    .b(sum_3[57]),
    .c(cout_4[56]),
    .cout(cout_4[57]),
    .sum(sum_4[57]));
  AL_FADD comp4_58 (
    .a(i4[58]),
    .b(sum_3[58]),
    .c(cout_4[57]),
    .cout(cout_4[58]),
    .sum(sum_4[58]));
  AL_FADD comp4_59 (
    .a(1'b0),
    .b(sum_3[59]),
    .c(cout_4[58]),
    .cout(cout_4[59]),
    .sum(sum_4[59]));
  AL_FADD comp4_6 (
    .a(i4[6]),
    .b(sum_3[6]),
    .c(cout_4[5]),
    .cout(cout_4[6]),
    .sum(sum_4[6]));
  AL_FADD comp4_60 (
    .a(1'b0),
    .b(sum_3[60]),
    .c(cout_4[59]),
    .cout(cout_4[60]),
    .sum(sum_4[60]));
  AL_FADD comp4_61 (
    .a(1'b0),
    .b(sum_3[61]),
    .c(cout_4[60]),
    .cout(cout_4[61]),
    .sum(sum_4[61]));
  AL_FADD comp4_62 (
    .a(1'b0),
    .b(sum_3[62]),
    .c(cout_4[61]),
    .cout(cout_4[62]),
    .sum(sum_4[62]));
  AL_FADD comp4_63 (
    .a(1'b0),
    .b(sum_3[63]),
    .c(cout_4[62]),
    .cout(cout_4[63]),
    .sum(sum_4[63]));
  AL_FADD comp4_7 (
    .a(i4[7]),
    .b(sum_3[7]),
    .c(cout_4[6]),
    .cout(cout_4[7]),
    .sum(sum_4[7]));
  AL_FADD comp4_8 (
    .a(i4[8]),
    .b(sum_3[8]),
    .c(cout_4[7]),
    .cout(cout_4[8]),
    .sum(sum_4[8]));
  AL_FADD comp4_9 (
    .a(i4[9]),
    .b(sum_3[9]),
    .c(cout_4[8]),
    .cout(cout_4[9]),
    .sum(sum_4[9]));
  AL_FADD comp5_0 (
    .a(i5[0]),
    .b(sum_4[0]),
    .c(1'b0),
    .cout(cout_5[0]),
    .sum(sum_5[0]));
  AL_FADD comp5_1 (
    .a(i5[1]),
    .b(sum_4[1]),
    .c(cout_5[0]),
    .cout(cout_5[1]),
    .sum(sum_5[1]));
  AL_FADD comp5_10 (
    .a(i5[10]),
    .b(sum_4[10]),
    .c(cout_5[9]),
    .cout(cout_5[10]),
    .sum(sum_5[10]));
  AL_FADD comp5_11 (
    .a(i5[11]),
    .b(sum_4[11]),
    .c(cout_5[10]),
    .cout(cout_5[11]),
    .sum(sum_5[11]));
  AL_FADD comp5_12 (
    .a(i5[12]),
    .b(sum_4[12]),
    .c(cout_5[11]),
    .cout(cout_5[12]),
    .sum(sum_5[12]));
  AL_FADD comp5_13 (
    .a(i5[13]),
    .b(sum_4[13]),
    .c(cout_5[12]),
    .cout(cout_5[13]),
    .sum(sum_5[13]));
  AL_FADD comp5_14 (
    .a(i5[14]),
    .b(sum_4[14]),
    .c(cout_5[13]),
    .cout(cout_5[14]),
    .sum(sum_5[14]));
  AL_FADD comp5_15 (
    .a(i5[15]),
    .b(sum_4[15]),
    .c(cout_5[14]),
    .cout(cout_5[15]),
    .sum(sum_5[15]));
  AL_FADD comp5_16 (
    .a(i5[16]),
    .b(sum_4[16]),
    .c(cout_5[15]),
    .cout(cout_5[16]),
    .sum(sum_5[16]));
  AL_FADD comp5_17 (
    .a(i5[17]),
    .b(sum_4[17]),
    .c(cout_5[16]),
    .cout(cout_5[17]),
    .sum(sum_5[17]));
  AL_FADD comp5_18 (
    .a(i5[18]),
    .b(sum_4[18]),
    .c(cout_5[17]),
    .cout(cout_5[18]),
    .sum(sum_5[18]));
  AL_FADD comp5_19 (
    .a(i5[19]),
    .b(sum_4[19]),
    .c(cout_5[18]),
    .cout(cout_5[19]),
    .sum(sum_5[19]));
  AL_FADD comp5_2 (
    .a(i5[2]),
    .b(sum_4[2]),
    .c(cout_5[1]),
    .cout(cout_5[2]),
    .sum(sum_5[2]));
  AL_FADD comp5_20 (
    .a(i5[20]),
    .b(sum_4[20]),
    .c(cout_5[19]),
    .cout(cout_5[20]),
    .sum(sum_5[20]));
  AL_FADD comp5_21 (
    .a(i5[21]),
    .b(sum_4[21]),
    .c(cout_5[20]),
    .cout(cout_5[21]),
    .sum(sum_5[21]));
  AL_FADD comp5_22 (
    .a(i5[22]),
    .b(sum_4[22]),
    .c(cout_5[21]),
    .cout(cout_5[22]),
    .sum(sum_5[22]));
  AL_FADD comp5_23 (
    .a(i5[23]),
    .b(sum_4[23]),
    .c(cout_5[22]),
    .cout(cout_5[23]),
    .sum(sum_5[23]));
  AL_FADD comp5_24 (
    .a(i5[24]),
    .b(sum_4[24]),
    .c(cout_5[23]),
    .cout(cout_5[24]),
    .sum(sum_5[24]));
  AL_FADD comp5_25 (
    .a(i5[25]),
    .b(sum_4[25]),
    .c(cout_5[24]),
    .cout(cout_5[25]),
    .sum(sum_5[25]));
  AL_FADD comp5_26 (
    .a(i5[26]),
    .b(sum_4[26]),
    .c(cout_5[25]),
    .cout(cout_5[26]),
    .sum(sum_5[26]));
  AL_FADD comp5_27 (
    .a(i5[27]),
    .b(sum_4[27]),
    .c(cout_5[26]),
    .cout(cout_5[27]),
    .sum(sum_5[27]));
  AL_FADD comp5_28 (
    .a(i5[28]),
    .b(sum_4[28]),
    .c(cout_5[27]),
    .cout(cout_5[28]),
    .sum(sum_5[28]));
  AL_FADD comp5_29 (
    .a(i5[29]),
    .b(sum_4[29]),
    .c(cout_5[28]),
    .cout(cout_5[29]),
    .sum(sum_5[29]));
  AL_FADD comp5_3 (
    .a(i5[3]),
    .b(sum_4[3]),
    .c(cout_5[2]),
    .cout(cout_5[3]),
    .sum(sum_5[3]));
  AL_FADD comp5_30 (
    .a(i5[30]),
    .b(sum_4[30]),
    .c(cout_5[29]),
    .cout(cout_5[30]),
    .sum(sum_5[30]));
  AL_FADD comp5_31 (
    .a(i5[31]),
    .b(sum_4[31]),
    .c(cout_5[30]),
    .cout(cout_5[31]),
    .sum(sum_5[31]));
  AL_FADD comp5_32 (
    .a(i5[32]),
    .b(sum_4[32]),
    .c(cout_5[31]),
    .cout(cout_5[32]),
    .sum(sum_5[32]));
  AL_FADD comp5_33 (
    .a(i5[33]),
    .b(sum_4[33]),
    .c(cout_5[32]),
    .cout(cout_5[33]),
    .sum(sum_5[33]));
  AL_FADD comp5_34 (
    .a(i5[34]),
    .b(sum_4[34]),
    .c(cout_5[33]),
    .cout(cout_5[34]),
    .sum(sum_5[34]));
  AL_FADD comp5_35 (
    .a(i5[35]),
    .b(sum_4[35]),
    .c(cout_5[34]),
    .cout(cout_5[35]),
    .sum(sum_5[35]));
  AL_FADD comp5_36 (
    .a(i5[36]),
    .b(sum_4[36]),
    .c(cout_5[35]),
    .cout(cout_5[36]),
    .sum(sum_5[36]));
  AL_FADD comp5_37 (
    .a(i5[37]),
    .b(sum_4[37]),
    .c(cout_5[36]),
    .cout(cout_5[37]),
    .sum(sum_5[37]));
  AL_FADD comp5_38 (
    .a(i5[38]),
    .b(sum_4[38]),
    .c(cout_5[37]),
    .cout(cout_5[38]),
    .sum(sum_5[38]));
  AL_FADD comp5_39 (
    .a(i5[39]),
    .b(sum_4[39]),
    .c(cout_5[38]),
    .cout(cout_5[39]),
    .sum(sum_5[39]));
  AL_FADD comp5_4 (
    .a(i5[4]),
    .b(sum_4[4]),
    .c(cout_5[3]),
    .cout(cout_5[4]),
    .sum(sum_5[4]));
  AL_FADD comp5_40 (
    .a(i5[40]),
    .b(sum_4[40]),
    .c(cout_5[39]),
    .cout(cout_5[40]),
    .sum(sum_5[40]));
  AL_FADD comp5_41 (
    .a(i5[41]),
    .b(sum_4[41]),
    .c(cout_5[40]),
    .cout(cout_5[41]),
    .sum(sum_5[41]));
  AL_FADD comp5_42 (
    .a(i5[42]),
    .b(sum_4[42]),
    .c(cout_5[41]),
    .cout(cout_5[42]),
    .sum(sum_5[42]));
  AL_FADD comp5_43 (
    .a(i5[43]),
    .b(sum_4[43]),
    .c(cout_5[42]),
    .cout(cout_5[43]),
    .sum(sum_5[43]));
  AL_FADD comp5_44 (
    .a(i5[44]),
    .b(sum_4[44]),
    .c(cout_5[43]),
    .cout(cout_5[44]),
    .sum(sum_5[44]));
  AL_FADD comp5_45 (
    .a(i5[45]),
    .b(sum_4[45]),
    .c(cout_5[44]),
    .cout(cout_5[45]),
    .sum(sum_5[45]));
  AL_FADD comp5_46 (
    .a(i5[46]),
    .b(sum_4[46]),
    .c(cout_5[45]),
    .cout(cout_5[46]),
    .sum(sum_5[46]));
  AL_FADD comp5_47 (
    .a(i5[47]),
    .b(sum_4[47]),
    .c(cout_5[46]),
    .cout(cout_5[47]),
    .sum(sum_5[47]));
  AL_FADD comp5_48 (
    .a(i5[48]),
    .b(sum_4[48]),
    .c(cout_5[47]),
    .cout(cout_5[48]),
    .sum(sum_5[48]));
  AL_FADD comp5_49 (
    .a(i5[49]),
    .b(sum_4[49]),
    .c(cout_5[48]),
    .cout(cout_5[49]),
    .sum(sum_5[49]));
  AL_FADD comp5_5 (
    .a(i5[5]),
    .b(sum_4[5]),
    .c(cout_5[4]),
    .cout(cout_5[5]),
    .sum(sum_5[5]));
  AL_FADD comp5_50 (
    .a(i5[50]),
    .b(sum_4[50]),
    .c(cout_5[49]),
    .cout(cout_5[50]),
    .sum(sum_5[50]));
  AL_FADD comp5_51 (
    .a(i5[51]),
    .b(sum_4[51]),
    .c(cout_5[50]),
    .cout(cout_5[51]),
    .sum(sum_5[51]));
  AL_FADD comp5_52 (
    .a(i5[52]),
    .b(sum_4[52]),
    .c(cout_5[51]),
    .cout(cout_5[52]),
    .sum(sum_5[52]));
  AL_FADD comp5_53 (
    .a(i5[53]),
    .b(sum_4[53]),
    .c(cout_5[52]),
    .cout(cout_5[53]),
    .sum(sum_5[53]));
  AL_FADD comp5_54 (
    .a(i5[54]),
    .b(sum_4[54]),
    .c(cout_5[53]),
    .cout(cout_5[54]),
    .sum(sum_5[54]));
  AL_FADD comp5_55 (
    .a(i5[55]),
    .b(sum_4[55]),
    .c(cout_5[54]),
    .cout(cout_5[55]),
    .sum(sum_5[55]));
  AL_FADD comp5_56 (
    .a(i5[56]),
    .b(sum_4[56]),
    .c(cout_5[55]),
    .cout(cout_5[56]),
    .sum(sum_5[56]));
  AL_FADD comp5_57 (
    .a(i5[57]),
    .b(sum_4[57]),
    .c(cout_5[56]),
    .cout(cout_5[57]),
    .sum(sum_5[57]));
  AL_FADD comp5_58 (
    .a(1'b0),
    .b(sum_4[58]),
    .c(cout_5[57]),
    .cout(cout_5[58]),
    .sum(sum_5[58]));
  AL_FADD comp5_59 (
    .a(1'b0),
    .b(sum_4[59]),
    .c(cout_5[58]),
    .cout(cout_5[59]),
    .sum(sum_5[59]));
  AL_FADD comp5_6 (
    .a(i5[6]),
    .b(sum_4[6]),
    .c(cout_5[5]),
    .cout(cout_5[6]),
    .sum(sum_5[6]));
  AL_FADD comp5_60 (
    .a(1'b0),
    .b(sum_4[60]),
    .c(cout_5[59]),
    .cout(cout_5[60]),
    .sum(sum_5[60]));
  AL_FADD comp5_61 (
    .a(1'b0),
    .b(sum_4[61]),
    .c(cout_5[60]),
    .cout(cout_5[61]),
    .sum(sum_5[61]));
  AL_FADD comp5_62 (
    .a(1'b0),
    .b(sum_4[62]),
    .c(cout_5[61]),
    .cout(cout_5[62]),
    .sum(sum_5[62]));
  AL_FADD comp5_63 (
    .a(1'b0),
    .b(sum_4[63]),
    .c(cout_5[62]),
    .cout(cout_5[63]),
    .sum(sum_5[63]));
  AL_FADD comp5_7 (
    .a(i5[7]),
    .b(sum_4[7]),
    .c(cout_5[6]),
    .cout(cout_5[7]),
    .sum(sum_5[7]));
  AL_FADD comp5_8 (
    .a(i5[8]),
    .b(sum_4[8]),
    .c(cout_5[7]),
    .cout(cout_5[8]),
    .sum(sum_5[8]));
  AL_FADD comp5_9 (
    .a(i5[9]),
    .b(sum_4[9]),
    .c(cout_5[8]),
    .cout(cout_5[9]),
    .sum(sum_5[9]));
  AL_FADD comp6_0 (
    .a(i6[0]),
    .b(sum_5[0]),
    .c(1'b0),
    .cout(cout_6[0]),
    .sum(sum_6[0]));
  AL_FADD comp6_1 (
    .a(i6[1]),
    .b(sum_5[1]),
    .c(cout_6[0]),
    .cout(cout_6[1]),
    .sum(sum_6[1]));
  AL_FADD comp6_10 (
    .a(i6[10]),
    .b(sum_5[10]),
    .c(cout_6[9]),
    .cout(cout_6[10]),
    .sum(sum_6[10]));
  AL_FADD comp6_11 (
    .a(i6[11]),
    .b(sum_5[11]),
    .c(cout_6[10]),
    .cout(cout_6[11]),
    .sum(sum_6[11]));
  AL_FADD comp6_12 (
    .a(i6[12]),
    .b(sum_5[12]),
    .c(cout_6[11]),
    .cout(cout_6[12]),
    .sum(sum_6[12]));
  AL_FADD comp6_13 (
    .a(i6[13]),
    .b(sum_5[13]),
    .c(cout_6[12]),
    .cout(cout_6[13]),
    .sum(sum_6[13]));
  AL_FADD comp6_14 (
    .a(i6[14]),
    .b(sum_5[14]),
    .c(cout_6[13]),
    .cout(cout_6[14]),
    .sum(sum_6[14]));
  AL_FADD comp6_15 (
    .a(i6[15]),
    .b(sum_5[15]),
    .c(cout_6[14]),
    .cout(cout_6[15]),
    .sum(sum_6[15]));
  AL_FADD comp6_16 (
    .a(i6[16]),
    .b(sum_5[16]),
    .c(cout_6[15]),
    .cout(cout_6[16]),
    .sum(sum_6[16]));
  AL_FADD comp6_17 (
    .a(i6[17]),
    .b(sum_5[17]),
    .c(cout_6[16]),
    .cout(cout_6[17]),
    .sum(sum_6[17]));
  AL_FADD comp6_18 (
    .a(i6[18]),
    .b(sum_5[18]),
    .c(cout_6[17]),
    .cout(cout_6[18]),
    .sum(sum_6[18]));
  AL_FADD comp6_19 (
    .a(i6[19]),
    .b(sum_5[19]),
    .c(cout_6[18]),
    .cout(cout_6[19]),
    .sum(sum_6[19]));
  AL_FADD comp6_2 (
    .a(i6[2]),
    .b(sum_5[2]),
    .c(cout_6[1]),
    .cout(cout_6[2]),
    .sum(sum_6[2]));
  AL_FADD comp6_20 (
    .a(i6[20]),
    .b(sum_5[20]),
    .c(cout_6[19]),
    .cout(cout_6[20]),
    .sum(sum_6[20]));
  AL_FADD comp6_21 (
    .a(i6[21]),
    .b(sum_5[21]),
    .c(cout_6[20]),
    .cout(cout_6[21]),
    .sum(sum_6[21]));
  AL_FADD comp6_22 (
    .a(i6[22]),
    .b(sum_5[22]),
    .c(cout_6[21]),
    .cout(cout_6[22]),
    .sum(sum_6[22]));
  AL_FADD comp6_23 (
    .a(i6[23]),
    .b(sum_5[23]),
    .c(cout_6[22]),
    .cout(cout_6[23]),
    .sum(sum_6[23]));
  AL_FADD comp6_24 (
    .a(i6[24]),
    .b(sum_5[24]),
    .c(cout_6[23]),
    .cout(cout_6[24]),
    .sum(sum_6[24]));
  AL_FADD comp6_25 (
    .a(i6[25]),
    .b(sum_5[25]),
    .c(cout_6[24]),
    .cout(cout_6[25]),
    .sum(sum_6[25]));
  AL_FADD comp6_26 (
    .a(i6[26]),
    .b(sum_5[26]),
    .c(cout_6[25]),
    .cout(cout_6[26]),
    .sum(sum_6[26]));
  AL_FADD comp6_27 (
    .a(i6[27]),
    .b(sum_5[27]),
    .c(cout_6[26]),
    .cout(cout_6[27]),
    .sum(sum_6[27]));
  AL_FADD comp6_28 (
    .a(i6[28]),
    .b(sum_5[28]),
    .c(cout_6[27]),
    .cout(cout_6[28]),
    .sum(sum_6[28]));
  AL_FADD comp6_29 (
    .a(i6[29]),
    .b(sum_5[29]),
    .c(cout_6[28]),
    .cout(cout_6[29]),
    .sum(sum_6[29]));
  AL_FADD comp6_3 (
    .a(i6[3]),
    .b(sum_5[3]),
    .c(cout_6[2]),
    .cout(cout_6[3]),
    .sum(sum_6[3]));
  AL_FADD comp6_30 (
    .a(i6[30]),
    .b(sum_5[30]),
    .c(cout_6[29]),
    .cout(cout_6[30]),
    .sum(sum_6[30]));
  AL_FADD comp6_31 (
    .a(i6[31]),
    .b(sum_5[31]),
    .c(cout_6[30]),
    .cout(cout_6[31]),
    .sum(sum_6[31]));
  AL_FADD comp6_32 (
    .a(i6[32]),
    .b(sum_5[32]),
    .c(cout_6[31]),
    .cout(cout_6[32]),
    .sum(sum_6[32]));
  AL_FADD comp6_33 (
    .a(i6[33]),
    .b(sum_5[33]),
    .c(cout_6[32]),
    .cout(cout_6[33]),
    .sum(sum_6[33]));
  AL_FADD comp6_34 (
    .a(i6[34]),
    .b(sum_5[34]),
    .c(cout_6[33]),
    .cout(cout_6[34]),
    .sum(sum_6[34]));
  AL_FADD comp6_35 (
    .a(i6[35]),
    .b(sum_5[35]),
    .c(cout_6[34]),
    .cout(cout_6[35]),
    .sum(sum_6[35]));
  AL_FADD comp6_36 (
    .a(i6[36]),
    .b(sum_5[36]),
    .c(cout_6[35]),
    .cout(cout_6[36]),
    .sum(sum_6[36]));
  AL_FADD comp6_37 (
    .a(i6[37]),
    .b(sum_5[37]),
    .c(cout_6[36]),
    .cout(cout_6[37]),
    .sum(sum_6[37]));
  AL_FADD comp6_38 (
    .a(i6[38]),
    .b(sum_5[38]),
    .c(cout_6[37]),
    .cout(cout_6[38]),
    .sum(sum_6[38]));
  AL_FADD comp6_39 (
    .a(i6[39]),
    .b(sum_5[39]),
    .c(cout_6[38]),
    .cout(cout_6[39]),
    .sum(sum_6[39]));
  AL_FADD comp6_4 (
    .a(i6[4]),
    .b(sum_5[4]),
    .c(cout_6[3]),
    .cout(cout_6[4]),
    .sum(sum_6[4]));
  AL_FADD comp6_40 (
    .a(i6[40]),
    .b(sum_5[40]),
    .c(cout_6[39]),
    .cout(cout_6[40]),
    .sum(sum_6[40]));
  AL_FADD comp6_41 (
    .a(i6[41]),
    .b(sum_5[41]),
    .c(cout_6[40]),
    .cout(cout_6[41]),
    .sum(sum_6[41]));
  AL_FADD comp6_42 (
    .a(i6[42]),
    .b(sum_5[42]),
    .c(cout_6[41]),
    .cout(cout_6[42]),
    .sum(sum_6[42]));
  AL_FADD comp6_43 (
    .a(i6[43]),
    .b(sum_5[43]),
    .c(cout_6[42]),
    .cout(cout_6[43]),
    .sum(sum_6[43]));
  AL_FADD comp6_44 (
    .a(i6[44]),
    .b(sum_5[44]),
    .c(cout_6[43]),
    .cout(cout_6[44]),
    .sum(sum_6[44]));
  AL_FADD comp6_45 (
    .a(i6[45]),
    .b(sum_5[45]),
    .c(cout_6[44]),
    .cout(cout_6[45]),
    .sum(sum_6[45]));
  AL_FADD comp6_46 (
    .a(i6[46]),
    .b(sum_5[46]),
    .c(cout_6[45]),
    .cout(cout_6[46]),
    .sum(sum_6[46]));
  AL_FADD comp6_47 (
    .a(i6[47]),
    .b(sum_5[47]),
    .c(cout_6[46]),
    .cout(cout_6[47]),
    .sum(sum_6[47]));
  AL_FADD comp6_48 (
    .a(i6[48]),
    .b(sum_5[48]),
    .c(cout_6[47]),
    .cout(cout_6[48]),
    .sum(sum_6[48]));
  AL_FADD comp6_49 (
    .a(i6[49]),
    .b(sum_5[49]),
    .c(cout_6[48]),
    .cout(cout_6[49]),
    .sum(sum_6[49]));
  AL_FADD comp6_5 (
    .a(i6[5]),
    .b(sum_5[5]),
    .c(cout_6[4]),
    .cout(cout_6[5]),
    .sum(sum_6[5]));
  AL_FADD comp6_50 (
    .a(i6[50]),
    .b(sum_5[50]),
    .c(cout_6[49]),
    .cout(cout_6[50]),
    .sum(sum_6[50]));
  AL_FADD comp6_51 (
    .a(i6[51]),
    .b(sum_5[51]),
    .c(cout_6[50]),
    .cout(cout_6[51]),
    .sum(sum_6[51]));
  AL_FADD comp6_52 (
    .a(i6[52]),
    .b(sum_5[52]),
    .c(cout_6[51]),
    .cout(cout_6[52]),
    .sum(sum_6[52]));
  AL_FADD comp6_53 (
    .a(i6[53]),
    .b(sum_5[53]),
    .c(cout_6[52]),
    .cout(cout_6[53]),
    .sum(sum_6[53]));
  AL_FADD comp6_54 (
    .a(i6[54]),
    .b(sum_5[54]),
    .c(cout_6[53]),
    .cout(cout_6[54]),
    .sum(sum_6[54]));
  AL_FADD comp6_55 (
    .a(i6[55]),
    .b(sum_5[55]),
    .c(cout_6[54]),
    .cout(cout_6[55]),
    .sum(sum_6[55]));
  AL_FADD comp6_56 (
    .a(i6[56]),
    .b(sum_5[56]),
    .c(cout_6[55]),
    .cout(cout_6[56]),
    .sum(sum_6[56]));
  AL_FADD comp6_57 (
    .a(1'b0),
    .b(sum_5[57]),
    .c(cout_6[56]),
    .cout(cout_6[57]),
    .sum(sum_6[57]));
  AL_FADD comp6_58 (
    .a(1'b0),
    .b(sum_5[58]),
    .c(cout_6[57]),
    .cout(cout_6[58]),
    .sum(sum_6[58]));
  AL_FADD comp6_59 (
    .a(1'b0),
    .b(sum_5[59]),
    .c(cout_6[58]),
    .cout(cout_6[59]),
    .sum(sum_6[59]));
  AL_FADD comp6_6 (
    .a(i6[6]),
    .b(sum_5[6]),
    .c(cout_6[5]),
    .cout(cout_6[6]),
    .sum(sum_6[6]));
  AL_FADD comp6_60 (
    .a(1'b0),
    .b(sum_5[60]),
    .c(cout_6[59]),
    .cout(cout_6[60]),
    .sum(sum_6[60]));
  AL_FADD comp6_61 (
    .a(1'b0),
    .b(sum_5[61]),
    .c(cout_6[60]),
    .cout(cout_6[61]),
    .sum(sum_6[61]));
  AL_FADD comp6_62 (
    .a(1'b0),
    .b(sum_5[62]),
    .c(cout_6[61]),
    .cout(cout_6[62]),
    .sum(sum_6[62]));
  AL_FADD comp6_63 (
    .a(1'b0),
    .b(sum_5[63]),
    .c(cout_6[62]),
    .cout(cout_6[63]),
    .sum(sum_6[63]));
  AL_FADD comp6_7 (
    .a(i6[7]),
    .b(sum_5[7]),
    .c(cout_6[6]),
    .cout(cout_6[7]),
    .sum(sum_6[7]));
  AL_FADD comp6_8 (
    .a(i6[8]),
    .b(sum_5[8]),
    .c(cout_6[7]),
    .cout(cout_6[8]),
    .sum(sum_6[8]));
  AL_FADD comp6_9 (
    .a(i6[9]),
    .b(sum_5[9]),
    .c(cout_6[8]),
    .cout(cout_6[9]),
    .sum(sum_6[9]));
  AL_FADD comp7_0 (
    .a(i7[0]),
    .b(sum_6[0]),
    .c(1'b0),
    .cout(cout_7[0]),
    .sum(sum_7[0]));
  AL_FADD comp7_1 (
    .a(i7[1]),
    .b(sum_6[1]),
    .c(cout_7[0]),
    .cout(cout_7[1]),
    .sum(sum_7[1]));
  AL_FADD comp7_10 (
    .a(i7[10]),
    .b(sum_6[10]),
    .c(cout_7[9]),
    .cout(cout_7[10]),
    .sum(sum_7[10]));
  AL_FADD comp7_11 (
    .a(i7[11]),
    .b(sum_6[11]),
    .c(cout_7[10]),
    .cout(cout_7[11]),
    .sum(sum_7[11]));
  AL_FADD comp7_12 (
    .a(i7[12]),
    .b(sum_6[12]),
    .c(cout_7[11]),
    .cout(cout_7[12]),
    .sum(sum_7[12]));
  AL_FADD comp7_13 (
    .a(i7[13]),
    .b(sum_6[13]),
    .c(cout_7[12]),
    .cout(cout_7[13]),
    .sum(sum_7[13]));
  AL_FADD comp7_14 (
    .a(i7[14]),
    .b(sum_6[14]),
    .c(cout_7[13]),
    .cout(cout_7[14]),
    .sum(sum_7[14]));
  AL_FADD comp7_15 (
    .a(i7[15]),
    .b(sum_6[15]),
    .c(cout_7[14]),
    .cout(cout_7[15]),
    .sum(sum_7[15]));
  AL_FADD comp7_16 (
    .a(i7[16]),
    .b(sum_6[16]),
    .c(cout_7[15]),
    .cout(cout_7[16]),
    .sum(sum_7[16]));
  AL_FADD comp7_17 (
    .a(i7[17]),
    .b(sum_6[17]),
    .c(cout_7[16]),
    .cout(cout_7[17]),
    .sum(sum_7[17]));
  AL_FADD comp7_18 (
    .a(i7[18]),
    .b(sum_6[18]),
    .c(cout_7[17]),
    .cout(cout_7[18]),
    .sum(sum_7[18]));
  AL_FADD comp7_19 (
    .a(i7[19]),
    .b(sum_6[19]),
    .c(cout_7[18]),
    .cout(cout_7[19]),
    .sum(sum_7[19]));
  AL_FADD comp7_2 (
    .a(i7[2]),
    .b(sum_6[2]),
    .c(cout_7[1]),
    .cout(cout_7[2]),
    .sum(sum_7[2]));
  AL_FADD comp7_20 (
    .a(i7[20]),
    .b(sum_6[20]),
    .c(cout_7[19]),
    .cout(cout_7[20]),
    .sum(sum_7[20]));
  AL_FADD comp7_21 (
    .a(i7[21]),
    .b(sum_6[21]),
    .c(cout_7[20]),
    .cout(cout_7[21]),
    .sum(sum_7[21]));
  AL_FADD comp7_22 (
    .a(i7[22]),
    .b(sum_6[22]),
    .c(cout_7[21]),
    .cout(cout_7[22]),
    .sum(sum_7[22]));
  AL_FADD comp7_23 (
    .a(i7[23]),
    .b(sum_6[23]),
    .c(cout_7[22]),
    .cout(cout_7[23]),
    .sum(sum_7[23]));
  AL_FADD comp7_24 (
    .a(i7[24]),
    .b(sum_6[24]),
    .c(cout_7[23]),
    .cout(cout_7[24]),
    .sum(sum_7[24]));
  AL_FADD comp7_25 (
    .a(i7[25]),
    .b(sum_6[25]),
    .c(cout_7[24]),
    .cout(cout_7[25]),
    .sum(sum_7[25]));
  AL_FADD comp7_26 (
    .a(i7[26]),
    .b(sum_6[26]),
    .c(cout_7[25]),
    .cout(cout_7[26]),
    .sum(sum_7[26]));
  AL_FADD comp7_27 (
    .a(i7[27]),
    .b(sum_6[27]),
    .c(cout_7[26]),
    .cout(cout_7[27]),
    .sum(sum_7[27]));
  AL_FADD comp7_28 (
    .a(i7[28]),
    .b(sum_6[28]),
    .c(cout_7[27]),
    .cout(cout_7[28]),
    .sum(sum_7[28]));
  AL_FADD comp7_29 (
    .a(i7[29]),
    .b(sum_6[29]),
    .c(cout_7[28]),
    .cout(cout_7[29]),
    .sum(sum_7[29]));
  AL_FADD comp7_3 (
    .a(i7[3]),
    .b(sum_6[3]),
    .c(cout_7[2]),
    .cout(cout_7[3]),
    .sum(sum_7[3]));
  AL_FADD comp7_30 (
    .a(i7[30]),
    .b(sum_6[30]),
    .c(cout_7[29]),
    .cout(cout_7[30]),
    .sum(sum_7[30]));
  AL_FADD comp7_31 (
    .a(i7[31]),
    .b(sum_6[31]),
    .c(cout_7[30]),
    .cout(cout_7[31]),
    .sum(sum_7[31]));
  AL_FADD comp7_32 (
    .a(i7[32]),
    .b(sum_6[32]),
    .c(cout_7[31]),
    .cout(cout_7[32]),
    .sum(sum_7[32]));
  AL_FADD comp7_33 (
    .a(i7[33]),
    .b(sum_6[33]),
    .c(cout_7[32]),
    .cout(cout_7[33]),
    .sum(sum_7[33]));
  AL_FADD comp7_34 (
    .a(i7[34]),
    .b(sum_6[34]),
    .c(cout_7[33]),
    .cout(cout_7[34]),
    .sum(sum_7[34]));
  AL_FADD comp7_35 (
    .a(i7[35]),
    .b(sum_6[35]),
    .c(cout_7[34]),
    .cout(cout_7[35]),
    .sum(sum_7[35]));
  AL_FADD comp7_36 (
    .a(i7[36]),
    .b(sum_6[36]),
    .c(cout_7[35]),
    .cout(cout_7[36]),
    .sum(sum_7[36]));
  AL_FADD comp7_37 (
    .a(i7[37]),
    .b(sum_6[37]),
    .c(cout_7[36]),
    .cout(cout_7[37]),
    .sum(sum_7[37]));
  AL_FADD comp7_38 (
    .a(i7[38]),
    .b(sum_6[38]),
    .c(cout_7[37]),
    .cout(cout_7[38]),
    .sum(sum_7[38]));
  AL_FADD comp7_39 (
    .a(i7[39]),
    .b(sum_6[39]),
    .c(cout_7[38]),
    .cout(cout_7[39]),
    .sum(sum_7[39]));
  AL_FADD comp7_4 (
    .a(i7[4]),
    .b(sum_6[4]),
    .c(cout_7[3]),
    .cout(cout_7[4]),
    .sum(sum_7[4]));
  AL_FADD comp7_40 (
    .a(i7[40]),
    .b(sum_6[40]),
    .c(cout_7[39]),
    .cout(cout_7[40]),
    .sum(sum_7[40]));
  AL_FADD comp7_41 (
    .a(i7[41]),
    .b(sum_6[41]),
    .c(cout_7[40]),
    .cout(cout_7[41]),
    .sum(sum_7[41]));
  AL_FADD comp7_42 (
    .a(i7[42]),
    .b(sum_6[42]),
    .c(cout_7[41]),
    .cout(cout_7[42]),
    .sum(sum_7[42]));
  AL_FADD comp7_43 (
    .a(i7[43]),
    .b(sum_6[43]),
    .c(cout_7[42]),
    .cout(cout_7[43]),
    .sum(sum_7[43]));
  AL_FADD comp7_44 (
    .a(i7[44]),
    .b(sum_6[44]),
    .c(cout_7[43]),
    .cout(cout_7[44]),
    .sum(sum_7[44]));
  AL_FADD comp7_45 (
    .a(i7[45]),
    .b(sum_6[45]),
    .c(cout_7[44]),
    .cout(cout_7[45]),
    .sum(sum_7[45]));
  AL_FADD comp7_46 (
    .a(i7[46]),
    .b(sum_6[46]),
    .c(cout_7[45]),
    .cout(cout_7[46]),
    .sum(sum_7[46]));
  AL_FADD comp7_47 (
    .a(i7[47]),
    .b(sum_6[47]),
    .c(cout_7[46]),
    .cout(cout_7[47]),
    .sum(sum_7[47]));
  AL_FADD comp7_48 (
    .a(i7[48]),
    .b(sum_6[48]),
    .c(cout_7[47]),
    .cout(cout_7[48]),
    .sum(sum_7[48]));
  AL_FADD comp7_49 (
    .a(i7[49]),
    .b(sum_6[49]),
    .c(cout_7[48]),
    .cout(cout_7[49]),
    .sum(sum_7[49]));
  AL_FADD comp7_5 (
    .a(i7[5]),
    .b(sum_6[5]),
    .c(cout_7[4]),
    .cout(cout_7[5]),
    .sum(sum_7[5]));
  AL_FADD comp7_50 (
    .a(i7[50]),
    .b(sum_6[50]),
    .c(cout_7[49]),
    .cout(cout_7[50]),
    .sum(sum_7[50]));
  AL_FADD comp7_51 (
    .a(i7[51]),
    .b(sum_6[51]),
    .c(cout_7[50]),
    .cout(cout_7[51]),
    .sum(sum_7[51]));
  AL_FADD comp7_52 (
    .a(i7[52]),
    .b(sum_6[52]),
    .c(cout_7[51]),
    .cout(cout_7[52]),
    .sum(sum_7[52]));
  AL_FADD comp7_53 (
    .a(i7[53]),
    .b(sum_6[53]),
    .c(cout_7[52]),
    .cout(cout_7[53]),
    .sum(sum_7[53]));
  AL_FADD comp7_54 (
    .a(i7[54]),
    .b(sum_6[54]),
    .c(cout_7[53]),
    .cout(cout_7[54]),
    .sum(sum_7[54]));
  AL_FADD comp7_55 (
    .a(i7[55]),
    .b(sum_6[55]),
    .c(cout_7[54]),
    .cout(cout_7[55]),
    .sum(sum_7[55]));
  AL_FADD comp7_56 (
    .a(1'b0),
    .b(sum_6[56]),
    .c(cout_7[55]),
    .cout(cout_7[56]),
    .sum(sum_7[56]));
  AL_FADD comp7_57 (
    .a(1'b0),
    .b(sum_6[57]),
    .c(cout_7[56]),
    .cout(cout_7[57]),
    .sum(sum_7[57]));
  AL_FADD comp7_58 (
    .a(1'b0),
    .b(sum_6[58]),
    .c(cout_7[57]),
    .cout(cout_7[58]),
    .sum(sum_7[58]));
  AL_FADD comp7_59 (
    .a(1'b0),
    .b(sum_6[59]),
    .c(cout_7[58]),
    .cout(cout_7[59]),
    .sum(sum_7[59]));
  AL_FADD comp7_6 (
    .a(i7[6]),
    .b(sum_6[6]),
    .c(cout_7[5]),
    .cout(cout_7[6]),
    .sum(sum_7[6]));
  AL_FADD comp7_60 (
    .a(1'b0),
    .b(sum_6[60]),
    .c(cout_7[59]),
    .cout(cout_7[60]),
    .sum(sum_7[60]));
  AL_FADD comp7_61 (
    .a(1'b0),
    .b(sum_6[61]),
    .c(cout_7[60]),
    .cout(cout_7[61]),
    .sum(sum_7[61]));
  AL_FADD comp7_62 (
    .a(1'b0),
    .b(sum_6[62]),
    .c(cout_7[61]),
    .cout(cout_7[62]),
    .sum(sum_7[62]));
  AL_FADD comp7_63 (
    .a(1'b0),
    .b(sum_6[63]),
    .c(cout_7[62]),
    .cout(cout_7[63]),
    .sum(sum_7[63]));
  AL_FADD comp7_7 (
    .a(i7[7]),
    .b(sum_6[7]),
    .c(cout_7[6]),
    .cout(cout_7[7]),
    .sum(sum_7[7]));
  AL_FADD comp7_8 (
    .a(i7[8]),
    .b(sum_6[8]),
    .c(cout_7[7]),
    .cout(cout_7[8]),
    .sum(sum_7[8]));
  AL_FADD comp7_9 (
    .a(i7[9]),
    .b(sum_6[9]),
    .c(cout_7[8]),
    .cout(cout_7[9]),
    .sum(sum_7[9]));
  AL_FADD comp8_0 (
    .a(i8[0]),
    .b(sum_7[0]),
    .c(1'b0),
    .cout(cout_8[0]),
    .sum(sum_8[0]));
  AL_FADD comp8_1 (
    .a(i8[1]),
    .b(sum_7[1]),
    .c(cout_8[0]),
    .cout(cout_8[1]),
    .sum(sum_8[1]));
  AL_FADD comp8_10 (
    .a(i8[10]),
    .b(sum_7[10]),
    .c(cout_8[9]),
    .cout(cout_8[10]),
    .sum(sum_8[10]));
  AL_FADD comp8_11 (
    .a(i8[11]),
    .b(sum_7[11]),
    .c(cout_8[10]),
    .cout(cout_8[11]),
    .sum(sum_8[11]));
  AL_FADD comp8_12 (
    .a(i8[12]),
    .b(sum_7[12]),
    .c(cout_8[11]),
    .cout(cout_8[12]),
    .sum(sum_8[12]));
  AL_FADD comp8_13 (
    .a(i8[13]),
    .b(sum_7[13]),
    .c(cout_8[12]),
    .cout(cout_8[13]),
    .sum(sum_8[13]));
  AL_FADD comp8_14 (
    .a(i8[14]),
    .b(sum_7[14]),
    .c(cout_8[13]),
    .cout(cout_8[14]),
    .sum(sum_8[14]));
  AL_FADD comp8_15 (
    .a(i8[15]),
    .b(sum_7[15]),
    .c(cout_8[14]),
    .cout(cout_8[15]),
    .sum(sum_8[15]));
  AL_FADD comp8_16 (
    .a(i8[16]),
    .b(sum_7[16]),
    .c(cout_8[15]),
    .cout(cout_8[16]),
    .sum(sum_8[16]));
  AL_FADD comp8_17 (
    .a(i8[17]),
    .b(sum_7[17]),
    .c(cout_8[16]),
    .cout(cout_8[17]),
    .sum(sum_8[17]));
  AL_FADD comp8_18 (
    .a(i8[18]),
    .b(sum_7[18]),
    .c(cout_8[17]),
    .cout(cout_8[18]),
    .sum(sum_8[18]));
  AL_FADD comp8_19 (
    .a(i8[19]),
    .b(sum_7[19]),
    .c(cout_8[18]),
    .cout(cout_8[19]),
    .sum(sum_8[19]));
  AL_FADD comp8_2 (
    .a(i8[2]),
    .b(sum_7[2]),
    .c(cout_8[1]),
    .cout(cout_8[2]),
    .sum(sum_8[2]));
  AL_FADD comp8_20 (
    .a(i8[20]),
    .b(sum_7[20]),
    .c(cout_8[19]),
    .cout(cout_8[20]),
    .sum(sum_8[20]));
  AL_FADD comp8_21 (
    .a(i8[21]),
    .b(sum_7[21]),
    .c(cout_8[20]),
    .cout(cout_8[21]),
    .sum(sum_8[21]));
  AL_FADD comp8_22 (
    .a(i8[22]),
    .b(sum_7[22]),
    .c(cout_8[21]),
    .cout(cout_8[22]),
    .sum(sum_8[22]));
  AL_FADD comp8_23 (
    .a(i8[23]),
    .b(sum_7[23]),
    .c(cout_8[22]),
    .cout(cout_8[23]),
    .sum(sum_8[23]));
  AL_FADD comp8_24 (
    .a(i8[24]),
    .b(sum_7[24]),
    .c(cout_8[23]),
    .cout(cout_8[24]),
    .sum(sum_8[24]));
  AL_FADD comp8_25 (
    .a(i8[25]),
    .b(sum_7[25]),
    .c(cout_8[24]),
    .cout(cout_8[25]),
    .sum(sum_8[25]));
  AL_FADD comp8_26 (
    .a(i8[26]),
    .b(sum_7[26]),
    .c(cout_8[25]),
    .cout(cout_8[26]),
    .sum(sum_8[26]));
  AL_FADD comp8_27 (
    .a(i8[27]),
    .b(sum_7[27]),
    .c(cout_8[26]),
    .cout(cout_8[27]),
    .sum(sum_8[27]));
  AL_FADD comp8_28 (
    .a(i8[28]),
    .b(sum_7[28]),
    .c(cout_8[27]),
    .cout(cout_8[28]),
    .sum(sum_8[28]));
  AL_FADD comp8_29 (
    .a(i8[29]),
    .b(sum_7[29]),
    .c(cout_8[28]),
    .cout(cout_8[29]),
    .sum(sum_8[29]));
  AL_FADD comp8_3 (
    .a(i8[3]),
    .b(sum_7[3]),
    .c(cout_8[2]),
    .cout(cout_8[3]),
    .sum(sum_8[3]));
  AL_FADD comp8_30 (
    .a(i8[30]),
    .b(sum_7[30]),
    .c(cout_8[29]),
    .cout(cout_8[30]),
    .sum(sum_8[30]));
  AL_FADD comp8_31 (
    .a(i8[31]),
    .b(sum_7[31]),
    .c(cout_8[30]),
    .cout(cout_8[31]),
    .sum(sum_8[31]));
  AL_FADD comp8_32 (
    .a(i8[32]),
    .b(sum_7[32]),
    .c(cout_8[31]),
    .cout(cout_8[32]),
    .sum(sum_8[32]));
  AL_FADD comp8_33 (
    .a(i8[33]),
    .b(sum_7[33]),
    .c(cout_8[32]),
    .cout(cout_8[33]),
    .sum(sum_8[33]));
  AL_FADD comp8_34 (
    .a(i8[34]),
    .b(sum_7[34]),
    .c(cout_8[33]),
    .cout(cout_8[34]),
    .sum(sum_8[34]));
  AL_FADD comp8_35 (
    .a(i8[35]),
    .b(sum_7[35]),
    .c(cout_8[34]),
    .cout(cout_8[35]),
    .sum(sum_8[35]));
  AL_FADD comp8_36 (
    .a(i8[36]),
    .b(sum_7[36]),
    .c(cout_8[35]),
    .cout(cout_8[36]),
    .sum(sum_8[36]));
  AL_FADD comp8_37 (
    .a(i8[37]),
    .b(sum_7[37]),
    .c(cout_8[36]),
    .cout(cout_8[37]),
    .sum(sum_8[37]));
  AL_FADD comp8_38 (
    .a(i8[38]),
    .b(sum_7[38]),
    .c(cout_8[37]),
    .cout(cout_8[38]),
    .sum(sum_8[38]));
  AL_FADD comp8_39 (
    .a(i8[39]),
    .b(sum_7[39]),
    .c(cout_8[38]),
    .cout(cout_8[39]),
    .sum(sum_8[39]));
  AL_FADD comp8_4 (
    .a(i8[4]),
    .b(sum_7[4]),
    .c(cout_8[3]),
    .cout(cout_8[4]),
    .sum(sum_8[4]));
  AL_FADD comp8_40 (
    .a(i8[40]),
    .b(sum_7[40]),
    .c(cout_8[39]),
    .cout(cout_8[40]),
    .sum(sum_8[40]));
  AL_FADD comp8_41 (
    .a(i8[41]),
    .b(sum_7[41]),
    .c(cout_8[40]),
    .cout(cout_8[41]),
    .sum(sum_8[41]));
  AL_FADD comp8_42 (
    .a(i8[42]),
    .b(sum_7[42]),
    .c(cout_8[41]),
    .cout(cout_8[42]),
    .sum(sum_8[42]));
  AL_FADD comp8_43 (
    .a(i8[43]),
    .b(sum_7[43]),
    .c(cout_8[42]),
    .cout(cout_8[43]),
    .sum(sum_8[43]));
  AL_FADD comp8_44 (
    .a(i8[44]),
    .b(sum_7[44]),
    .c(cout_8[43]),
    .cout(cout_8[44]),
    .sum(sum_8[44]));
  AL_FADD comp8_45 (
    .a(i8[45]),
    .b(sum_7[45]),
    .c(cout_8[44]),
    .cout(cout_8[45]),
    .sum(sum_8[45]));
  AL_FADD comp8_46 (
    .a(i8[46]),
    .b(sum_7[46]),
    .c(cout_8[45]),
    .cout(cout_8[46]),
    .sum(sum_8[46]));
  AL_FADD comp8_47 (
    .a(i8[47]),
    .b(sum_7[47]),
    .c(cout_8[46]),
    .cout(cout_8[47]),
    .sum(sum_8[47]));
  AL_FADD comp8_48 (
    .a(i8[48]),
    .b(sum_7[48]),
    .c(cout_8[47]),
    .cout(cout_8[48]),
    .sum(sum_8[48]));
  AL_FADD comp8_49 (
    .a(i8[49]),
    .b(sum_7[49]),
    .c(cout_8[48]),
    .cout(cout_8[49]),
    .sum(sum_8[49]));
  AL_FADD comp8_5 (
    .a(i8[5]),
    .b(sum_7[5]),
    .c(cout_8[4]),
    .cout(cout_8[5]),
    .sum(sum_8[5]));
  AL_FADD comp8_50 (
    .a(i8[50]),
    .b(sum_7[50]),
    .c(cout_8[49]),
    .cout(cout_8[50]),
    .sum(sum_8[50]));
  AL_FADD comp8_51 (
    .a(i8[51]),
    .b(sum_7[51]),
    .c(cout_8[50]),
    .cout(cout_8[51]),
    .sum(sum_8[51]));
  AL_FADD comp8_52 (
    .a(i8[52]),
    .b(sum_7[52]),
    .c(cout_8[51]),
    .cout(cout_8[52]),
    .sum(sum_8[52]));
  AL_FADD comp8_53 (
    .a(i8[53]),
    .b(sum_7[53]),
    .c(cout_8[52]),
    .cout(cout_8[53]),
    .sum(sum_8[53]));
  AL_FADD comp8_54 (
    .a(i8[54]),
    .b(sum_7[54]),
    .c(cout_8[53]),
    .cout(cout_8[54]),
    .sum(sum_8[54]));
  AL_FADD comp8_55 (
    .a(1'b0),
    .b(sum_7[55]),
    .c(cout_8[54]),
    .cout(cout_8[55]),
    .sum(sum_8[55]));
  AL_FADD comp8_56 (
    .a(1'b0),
    .b(sum_7[56]),
    .c(cout_8[55]),
    .cout(cout_8[56]),
    .sum(sum_8[56]));
  AL_FADD comp8_57 (
    .a(1'b0),
    .b(sum_7[57]),
    .c(cout_8[56]),
    .cout(cout_8[57]),
    .sum(sum_8[57]));
  AL_FADD comp8_58 (
    .a(1'b0),
    .b(sum_7[58]),
    .c(cout_8[57]),
    .cout(cout_8[58]),
    .sum(sum_8[58]));
  AL_FADD comp8_59 (
    .a(1'b0),
    .b(sum_7[59]),
    .c(cout_8[58]),
    .cout(cout_8[59]),
    .sum(sum_8[59]));
  AL_FADD comp8_6 (
    .a(i8[6]),
    .b(sum_7[6]),
    .c(cout_8[5]),
    .cout(cout_8[6]),
    .sum(sum_8[6]));
  AL_FADD comp8_60 (
    .a(1'b0),
    .b(sum_7[60]),
    .c(cout_8[59]),
    .cout(cout_8[60]),
    .sum(sum_8[60]));
  AL_FADD comp8_61 (
    .a(1'b0),
    .b(sum_7[61]),
    .c(cout_8[60]),
    .cout(cout_8[61]),
    .sum(sum_8[61]));
  AL_FADD comp8_62 (
    .a(1'b0),
    .b(sum_7[62]),
    .c(cout_8[61]),
    .cout(cout_8[62]),
    .sum(sum_8[62]));
  AL_FADD comp8_63 (
    .a(1'b0),
    .b(sum_7[63]),
    .c(cout_8[62]),
    .cout(cout_8[63]),
    .sum(sum_8[63]));
  AL_FADD comp8_7 (
    .a(i8[7]),
    .b(sum_7[7]),
    .c(cout_8[6]),
    .cout(cout_8[7]),
    .sum(sum_8[7]));
  AL_FADD comp8_8 (
    .a(i8[8]),
    .b(sum_7[8]),
    .c(cout_8[7]),
    .cout(cout_8[8]),
    .sum(sum_8[8]));
  AL_FADD comp8_9 (
    .a(i8[9]),
    .b(sum_7[9]),
    .c(cout_8[8]),
    .cout(cout_8[9]),
    .sum(sum_8[9]));
  AL_FADD comp9_0 (
    .a(i9[0]),
    .b(sum_8[0]),
    .c(1'b0),
    .cout(cout_9[0]),
    .sum(sum_9[0]));
  AL_FADD comp9_1 (
    .a(i9[1]),
    .b(sum_8[1]),
    .c(cout_9[0]),
    .cout(cout_9[1]),
    .sum(sum_9[1]));
  AL_FADD comp9_10 (
    .a(i9[10]),
    .b(sum_8[10]),
    .c(cout_9[9]),
    .cout(cout_9[10]),
    .sum(sum_9[10]));
  AL_FADD comp9_11 (
    .a(i9[11]),
    .b(sum_8[11]),
    .c(cout_9[10]),
    .cout(cout_9[11]),
    .sum(sum_9[11]));
  AL_FADD comp9_12 (
    .a(i9[12]),
    .b(sum_8[12]),
    .c(cout_9[11]),
    .cout(cout_9[12]),
    .sum(sum_9[12]));
  AL_FADD comp9_13 (
    .a(i9[13]),
    .b(sum_8[13]),
    .c(cout_9[12]),
    .cout(cout_9[13]),
    .sum(sum_9[13]));
  AL_FADD comp9_14 (
    .a(i9[14]),
    .b(sum_8[14]),
    .c(cout_9[13]),
    .cout(cout_9[14]),
    .sum(sum_9[14]));
  AL_FADD comp9_15 (
    .a(i9[15]),
    .b(sum_8[15]),
    .c(cout_9[14]),
    .cout(cout_9[15]),
    .sum(sum_9[15]));
  AL_FADD comp9_16 (
    .a(i9[16]),
    .b(sum_8[16]),
    .c(cout_9[15]),
    .cout(cout_9[16]),
    .sum(sum_9[16]));
  AL_FADD comp9_17 (
    .a(i9[17]),
    .b(sum_8[17]),
    .c(cout_9[16]),
    .cout(cout_9[17]),
    .sum(sum_9[17]));
  AL_FADD comp9_18 (
    .a(i9[18]),
    .b(sum_8[18]),
    .c(cout_9[17]),
    .cout(cout_9[18]),
    .sum(sum_9[18]));
  AL_FADD comp9_19 (
    .a(i9[19]),
    .b(sum_8[19]),
    .c(cout_9[18]),
    .cout(cout_9[19]),
    .sum(sum_9[19]));
  AL_FADD comp9_2 (
    .a(i9[2]),
    .b(sum_8[2]),
    .c(cout_9[1]),
    .cout(cout_9[2]),
    .sum(sum_9[2]));
  AL_FADD comp9_20 (
    .a(i9[20]),
    .b(sum_8[20]),
    .c(cout_9[19]),
    .cout(cout_9[20]),
    .sum(sum_9[20]));
  AL_FADD comp9_21 (
    .a(i9[21]),
    .b(sum_8[21]),
    .c(cout_9[20]),
    .cout(cout_9[21]),
    .sum(sum_9[21]));
  AL_FADD comp9_22 (
    .a(i9[22]),
    .b(sum_8[22]),
    .c(cout_9[21]),
    .cout(cout_9[22]),
    .sum(sum_9[22]));
  AL_FADD comp9_23 (
    .a(i9[23]),
    .b(sum_8[23]),
    .c(cout_9[22]),
    .cout(cout_9[23]),
    .sum(sum_9[23]));
  AL_FADD comp9_24 (
    .a(i9[24]),
    .b(sum_8[24]),
    .c(cout_9[23]),
    .cout(cout_9[24]),
    .sum(sum_9[24]));
  AL_FADD comp9_25 (
    .a(i9[25]),
    .b(sum_8[25]),
    .c(cout_9[24]),
    .cout(cout_9[25]),
    .sum(sum_9[25]));
  AL_FADD comp9_26 (
    .a(i9[26]),
    .b(sum_8[26]),
    .c(cout_9[25]),
    .cout(cout_9[26]),
    .sum(sum_9[26]));
  AL_FADD comp9_27 (
    .a(i9[27]),
    .b(sum_8[27]),
    .c(cout_9[26]),
    .cout(cout_9[27]),
    .sum(sum_9[27]));
  AL_FADD comp9_28 (
    .a(i9[28]),
    .b(sum_8[28]),
    .c(cout_9[27]),
    .cout(cout_9[28]),
    .sum(sum_9[28]));
  AL_FADD comp9_29 (
    .a(i9[29]),
    .b(sum_8[29]),
    .c(cout_9[28]),
    .cout(cout_9[29]),
    .sum(sum_9[29]));
  AL_FADD comp9_3 (
    .a(i9[3]),
    .b(sum_8[3]),
    .c(cout_9[2]),
    .cout(cout_9[3]),
    .sum(sum_9[3]));
  AL_FADD comp9_30 (
    .a(i9[30]),
    .b(sum_8[30]),
    .c(cout_9[29]),
    .cout(cout_9[30]),
    .sum(sum_9[30]));
  AL_FADD comp9_31 (
    .a(i9[31]),
    .b(sum_8[31]),
    .c(cout_9[30]),
    .cout(cout_9[31]),
    .sum(sum_9[31]));
  AL_FADD comp9_32 (
    .a(i9[32]),
    .b(sum_8[32]),
    .c(cout_9[31]),
    .cout(cout_9[32]),
    .sum(sum_9[32]));
  AL_FADD comp9_33 (
    .a(i9[33]),
    .b(sum_8[33]),
    .c(cout_9[32]),
    .cout(cout_9[33]),
    .sum(sum_9[33]));
  AL_FADD comp9_34 (
    .a(i9[34]),
    .b(sum_8[34]),
    .c(cout_9[33]),
    .cout(cout_9[34]),
    .sum(sum_9[34]));
  AL_FADD comp9_35 (
    .a(i9[35]),
    .b(sum_8[35]),
    .c(cout_9[34]),
    .cout(cout_9[35]),
    .sum(sum_9[35]));
  AL_FADD comp9_36 (
    .a(i9[36]),
    .b(sum_8[36]),
    .c(cout_9[35]),
    .cout(cout_9[36]),
    .sum(sum_9[36]));
  AL_FADD comp9_37 (
    .a(i9[37]),
    .b(sum_8[37]),
    .c(cout_9[36]),
    .cout(cout_9[37]),
    .sum(sum_9[37]));
  AL_FADD comp9_38 (
    .a(i9[38]),
    .b(sum_8[38]),
    .c(cout_9[37]),
    .cout(cout_9[38]),
    .sum(sum_9[38]));
  AL_FADD comp9_39 (
    .a(i9[39]),
    .b(sum_8[39]),
    .c(cout_9[38]),
    .cout(cout_9[39]),
    .sum(sum_9[39]));
  AL_FADD comp9_4 (
    .a(i9[4]),
    .b(sum_8[4]),
    .c(cout_9[3]),
    .cout(cout_9[4]),
    .sum(sum_9[4]));
  AL_FADD comp9_40 (
    .a(i9[40]),
    .b(sum_8[40]),
    .c(cout_9[39]),
    .cout(cout_9[40]),
    .sum(sum_9[40]));
  AL_FADD comp9_41 (
    .a(i9[41]),
    .b(sum_8[41]),
    .c(cout_9[40]),
    .cout(cout_9[41]),
    .sum(sum_9[41]));
  AL_FADD comp9_42 (
    .a(i9[42]),
    .b(sum_8[42]),
    .c(cout_9[41]),
    .cout(cout_9[42]),
    .sum(sum_9[42]));
  AL_FADD comp9_43 (
    .a(i9[43]),
    .b(sum_8[43]),
    .c(cout_9[42]),
    .cout(cout_9[43]),
    .sum(sum_9[43]));
  AL_FADD comp9_44 (
    .a(i9[44]),
    .b(sum_8[44]),
    .c(cout_9[43]),
    .cout(cout_9[44]),
    .sum(sum_9[44]));
  AL_FADD comp9_45 (
    .a(i9[45]),
    .b(sum_8[45]),
    .c(cout_9[44]),
    .cout(cout_9[45]),
    .sum(sum_9[45]));
  AL_FADD comp9_46 (
    .a(i9[46]),
    .b(sum_8[46]),
    .c(cout_9[45]),
    .cout(cout_9[46]),
    .sum(sum_9[46]));
  AL_FADD comp9_47 (
    .a(i9[47]),
    .b(sum_8[47]),
    .c(cout_9[46]),
    .cout(cout_9[47]),
    .sum(sum_9[47]));
  AL_FADD comp9_48 (
    .a(i9[48]),
    .b(sum_8[48]),
    .c(cout_9[47]),
    .cout(cout_9[48]),
    .sum(sum_9[48]));
  AL_FADD comp9_49 (
    .a(i9[49]),
    .b(sum_8[49]),
    .c(cout_9[48]),
    .cout(cout_9[49]),
    .sum(sum_9[49]));
  AL_FADD comp9_5 (
    .a(i9[5]),
    .b(sum_8[5]),
    .c(cout_9[4]),
    .cout(cout_9[5]),
    .sum(sum_9[5]));
  AL_FADD comp9_50 (
    .a(i9[50]),
    .b(sum_8[50]),
    .c(cout_9[49]),
    .cout(cout_9[50]),
    .sum(sum_9[50]));
  AL_FADD comp9_51 (
    .a(i9[51]),
    .b(sum_8[51]),
    .c(cout_9[50]),
    .cout(cout_9[51]),
    .sum(sum_9[51]));
  AL_FADD comp9_52 (
    .a(i9[52]),
    .b(sum_8[52]),
    .c(cout_9[51]),
    .cout(cout_9[52]),
    .sum(sum_9[52]));
  AL_FADD comp9_53 (
    .a(i9[53]),
    .b(sum_8[53]),
    .c(cout_9[52]),
    .cout(cout_9[53]),
    .sum(sum_9[53]));
  AL_FADD comp9_54 (
    .a(1'b0),
    .b(sum_8[54]),
    .c(cout_9[53]),
    .cout(cout_9[54]),
    .sum(sum_9[54]));
  AL_FADD comp9_55 (
    .a(1'b0),
    .b(sum_8[55]),
    .c(cout_9[54]),
    .cout(cout_9[55]),
    .sum(sum_9[55]));
  AL_FADD comp9_56 (
    .a(1'b0),
    .b(sum_8[56]),
    .c(cout_9[55]),
    .cout(cout_9[56]),
    .sum(sum_9[56]));
  AL_FADD comp9_57 (
    .a(1'b0),
    .b(sum_8[57]),
    .c(cout_9[56]),
    .cout(cout_9[57]),
    .sum(sum_9[57]));
  AL_FADD comp9_58 (
    .a(1'b0),
    .b(sum_8[58]),
    .c(cout_9[57]),
    .cout(cout_9[58]),
    .sum(sum_9[58]));
  AL_FADD comp9_59 (
    .a(1'b0),
    .b(sum_8[59]),
    .c(cout_9[58]),
    .cout(cout_9[59]),
    .sum(sum_9[59]));
  AL_FADD comp9_6 (
    .a(i9[6]),
    .b(sum_8[6]),
    .c(cout_9[5]),
    .cout(cout_9[6]),
    .sum(sum_9[6]));
  AL_FADD comp9_60 (
    .a(1'b0),
    .b(sum_8[60]),
    .c(cout_9[59]),
    .cout(cout_9[60]),
    .sum(sum_9[60]));
  AL_FADD comp9_61 (
    .a(1'b0),
    .b(sum_8[61]),
    .c(cout_9[60]),
    .cout(cout_9[61]),
    .sum(sum_9[61]));
  AL_FADD comp9_62 (
    .a(1'b0),
    .b(sum_8[62]),
    .c(cout_9[61]),
    .cout(cout_9[62]),
    .sum(sum_9[62]));
  AL_FADD comp9_63 (
    .a(1'b0),
    .b(sum_8[63]),
    .c(cout_9[62]),
    .cout(cout_9[63]),
    .sum(sum_9[63]));
  AL_FADD comp9_7 (
    .a(i9[7]),
    .b(sum_8[7]),
    .c(cout_9[6]),
    .cout(cout_9[7]),
    .sum(sum_9[7]));
  AL_FADD comp9_8 (
    .a(i9[8]),
    .b(sum_8[8]),
    .c(cout_9[7]),
    .cout(cout_9[8]),
    .sum(sum_9[8]));
  AL_FADD comp9_9 (
    .a(i9[9]),
    .b(sum_8[9]),
    .c(cout_9[8]),
    .cout(cout_9[9]),
    .sum(sum_9[9]));

endmodule 

module add_pu64_pu61_pu60_pu59_pu58_pu57_pu56_pu55_pu54_pu53_pu52_pu51_pu50_pu49_pu48_pu47_pu46_pu45_pu44_pu43_pu42_pu41_pu40_pu39_pu38_pu37_pu36_pu35_pu34_pu33_pu32_mu63_mu63_o64
  (
  i0,
  i1,
  i10,
  i11,
  i12,
  i13,
  i14,
  i15,
  i16,
  i17,
  i18,
  i19,
  i2,
  i20,
  i21,
  i22,
  i23,
  i24,
  i25,
  i26,
  i27,
  i28,
  i29,
  i3,
  i30,
  i31,
  i32,
  i4,
  i5,
  i6,
  i7,
  i8,
  i9,
  o
  );

  input [63:0] i0;
  input [60:0] i1;
  input [51:0] i10;
  input [50:0] i11;
  input [49:0] i12;
  input [48:0] i13;
  input [47:0] i14;
  input [46:0] i15;
  input [45:0] i16;
  input [44:0] i17;
  input [43:0] i18;
  input [42:0] i19;
  input [59:0] i2;
  input [41:0] i20;
  input [40:0] i21;
  input [39:0] i22;
  input [38:0] i23;
  input [37:0] i24;
  input [36:0] i25;
  input [35:0] i26;
  input [34:0] i27;
  input [33:0] i28;
  input [32:0] i29;
  input [58:0] i3;
  input [31:0] i30;
  input [62:0] i31;
  input [62:0] i32;
  input [57:0] i4;
  input [56:0] i5;
  input [55:0] i6;
  input [54:0] i7;
  input [53:0] i8;
  input [52:0] i9;
  output [63:0] o;

  wire [63:0] cout_1;
  wire [63:0] cout_10;
  wire [63:0] cout_11;
  wire [63:0] cout_12;
  wire [63:0] cout_13;
  wire [63:0] cout_14;
  wire [63:0] cout_15;
  wire [63:0] cout_16;
  wire [63:0] cout_17;
  wire [63:0] cout_18;
  wire [63:0] cout_19;
  wire [63:0] cout_2;
  wire [63:0] cout_20;
  wire [63:0] cout_21;
  wire [63:0] cout_22;
  wire [63:0] cout_23;
  wire [63:0] cout_24;
  wire [63:0] cout_25;
  wire [63:0] cout_26;
  wire [63:0] cout_27;
  wire [63:0] cout_28;
  wire [63:0] cout_29;
  wire [63:0] cout_3;
  wire [63:0] cout_30;
  wire [63:0] cout_31;
  wire [63:0] cout_32;
  wire [63:0] cout_4;
  wire [63:0] cout_5;
  wire [63:0] cout_6;
  wire [63:0] cout_7;
  wire [63:0] cout_8;
  wire [63:0] cout_9;
  wire [63:0] sum_1;
  wire [63:0] sum_10;
  wire [63:0] sum_11;
  wire [63:0] sum_12;
  wire [63:0] sum_13;
  wire [63:0] sum_14;
  wire [63:0] sum_15;
  wire [63:0] sum_16;
  wire [63:0] sum_17;
  wire [63:0] sum_18;
  wire [63:0] sum_19;
  wire [63:0] sum_2;
  wire [63:0] sum_20;
  wire [63:0] sum_21;
  wire [63:0] sum_22;
  wire [63:0] sum_23;
  wire [63:0] sum_24;
  wire [63:0] sum_25;
  wire [63:0] sum_26;
  wire [63:0] sum_27;
  wire [63:0] sum_28;
  wire [63:0] sum_29;
  wire [63:0] sum_3;
  wire [63:0] sum_30;
  wire [63:0] sum_31;
  wire [63:0] sum_32;
  wire [63:0] sum_4;
  wire [63:0] sum_5;
  wire [63:0] sum_6;
  wire [63:0] sum_7;
  wire [63:0] sum_8;
  wire [63:0] sum_9;
  wire net_nb31_0;
  wire net_nb31_1;
  wire net_nb31_10;
  wire net_nb31_11;
  wire net_nb31_12;
  wire net_nb31_13;
  wire net_nb31_14;
  wire net_nb31_15;
  wire net_nb31_16;
  wire net_nb31_17;
  wire net_nb31_18;
  wire net_nb31_19;
  wire net_nb31_2;
  wire net_nb31_20;
  wire net_nb31_21;
  wire net_nb31_22;
  wire net_nb31_23;
  wire net_nb31_24;
  wire net_nb31_25;
  wire net_nb31_26;
  wire net_nb31_27;
  wire net_nb31_28;
  wire net_nb31_29;
  wire net_nb31_3;
  wire net_nb31_30;
  wire net_nb31_31;
  wire net_nb31_32;
  wire net_nb31_33;
  wire net_nb31_34;
  wire net_nb31_35;
  wire net_nb31_36;
  wire net_nb31_37;
  wire net_nb31_38;
  wire net_nb31_39;
  wire net_nb31_4;
  wire net_nb31_40;
  wire net_nb31_41;
  wire net_nb31_42;
  wire net_nb31_43;
  wire net_nb31_44;
  wire net_nb31_45;
  wire net_nb31_46;
  wire net_nb31_47;
  wire net_nb31_48;
  wire net_nb31_49;
  wire net_nb31_5;
  wire net_nb31_50;
  wire net_nb31_51;
  wire net_nb31_52;
  wire net_nb31_53;
  wire net_nb31_54;
  wire net_nb31_55;
  wire net_nb31_56;
  wire net_nb31_57;
  wire net_nb31_58;
  wire net_nb31_59;
  wire net_nb31_6;
  wire net_nb31_60;
  wire net_nb31_61;
  wire net_nb31_62;
  wire net_nb31_63;
  wire net_nb31_7;
  wire net_nb31_8;
  wire net_nb31_9;
  wire net_nb32_0;
  wire net_nb32_1;
  wire net_nb32_10;
  wire net_nb32_11;
  wire net_nb32_12;
  wire net_nb32_13;
  wire net_nb32_14;
  wire net_nb32_15;
  wire net_nb32_16;
  wire net_nb32_17;
  wire net_nb32_18;
  wire net_nb32_19;
  wire net_nb32_2;
  wire net_nb32_20;
  wire net_nb32_21;
  wire net_nb32_22;
  wire net_nb32_23;
  wire net_nb32_24;
  wire net_nb32_25;
  wire net_nb32_26;
  wire net_nb32_27;
  wire net_nb32_28;
  wire net_nb32_29;
  wire net_nb32_3;
  wire net_nb32_30;
  wire net_nb32_31;
  wire net_nb32_32;
  wire net_nb32_33;
  wire net_nb32_34;
  wire net_nb32_35;
  wire net_nb32_36;
  wire net_nb32_37;
  wire net_nb32_38;
  wire net_nb32_39;
  wire net_nb32_4;
  wire net_nb32_40;
  wire net_nb32_41;
  wire net_nb32_42;
  wire net_nb32_43;
  wire net_nb32_44;
  wire net_nb32_45;
  wire net_nb32_46;
  wire net_nb32_47;
  wire net_nb32_48;
  wire net_nb32_49;
  wire net_nb32_5;
  wire net_nb32_50;
  wire net_nb32_51;
  wire net_nb32_52;
  wire net_nb32_53;
  wire net_nb32_54;
  wire net_nb32_55;
  wire net_nb32_56;
  wire net_nb32_57;
  wire net_nb32_58;
  wire net_nb32_59;
  wire net_nb32_6;
  wire net_nb32_60;
  wire net_nb32_61;
  wire net_nb32_62;
  wire net_nb32_63;
  wire net_nb32_7;
  wire net_nb32_8;
  wire net_nb32_9;
  wire net_ncout31_63;
  wire net_ncout32_63;

  assign o[63] = sum_32[63];
  assign o[62] = sum_32[62];
  assign o[61] = sum_32[61];
  assign o[60] = sum_32[60];
  assign o[59] = sum_32[59];
  assign o[58] = sum_32[58];
  assign o[57] = sum_32[57];
  assign o[56] = sum_32[56];
  assign o[55] = sum_32[55];
  assign o[54] = sum_32[54];
  assign o[53] = sum_32[53];
  assign o[52] = sum_32[52];
  assign o[51] = sum_32[51];
  assign o[50] = sum_32[50];
  assign o[49] = sum_32[49];
  assign o[48] = sum_32[48];
  assign o[47] = sum_32[47];
  assign o[46] = sum_32[46];
  assign o[45] = sum_32[45];
  assign o[44] = sum_32[44];
  assign o[43] = sum_32[43];
  assign o[42] = sum_32[42];
  assign o[41] = sum_32[41];
  assign o[40] = sum_32[40];
  assign o[39] = sum_32[39];
  assign o[38] = sum_32[38];
  assign o[37] = sum_32[37];
  assign o[36] = sum_32[36];
  assign o[35] = sum_32[35];
  assign o[34] = sum_32[34];
  assign o[33] = sum_32[33];
  assign o[32] = sum_32[32];
  assign o[31] = sum_32[31];
  assign o[30] = sum_32[30];
  assign o[29] = sum_32[29];
  assign o[28] = sum_32[28];
  assign o[27] = sum_32[27];
  assign o[26] = sum_32[26];
  assign o[25] = sum_32[25];
  assign o[24] = sum_32[24];
  assign o[23] = sum_32[23];
  assign o[22] = sum_32[22];
  assign o[21] = sum_32[21];
  assign o[20] = sum_32[20];
  assign o[19] = sum_32[19];
  assign o[18] = sum_32[18];
  assign o[17] = sum_32[17];
  assign o[16] = sum_32[16];
  assign o[15] = sum_32[15];
  assign o[14] = sum_32[14];
  assign o[13] = sum_32[13];
  assign o[12] = sum_32[12];
  assign o[11] = sum_32[11];
  assign o[10] = sum_32[10];
  assign o[9] = sum_32[9];
  assign o[8] = sum_32[8];
  assign o[7] = sum_32[7];
  assign o[6] = sum_32[6];
  assign o[5] = sum_32[5];
  assign o[4] = sum_32[4];
  assign o[3] = sum_32[3];
  assign o[2] = sum_32[2];
  assign o[1] = sum_32[1];
  assign o[0] = sum_32[0];
  AL_FADD comp10_0 (
    .a(i10[0]),
    .b(sum_9[0]),
    .c(1'b0),
    .cout(cout_10[0]),
    .sum(sum_10[0]));
  AL_FADD comp10_1 (
    .a(i10[1]),
    .b(sum_9[1]),
    .c(cout_10[0]),
    .cout(cout_10[1]),
    .sum(sum_10[1]));
  AL_FADD comp10_10 (
    .a(i10[10]),
    .b(sum_9[10]),
    .c(cout_10[9]),
    .cout(cout_10[10]),
    .sum(sum_10[10]));
  AL_FADD comp10_11 (
    .a(i10[11]),
    .b(sum_9[11]),
    .c(cout_10[10]),
    .cout(cout_10[11]),
    .sum(sum_10[11]));
  AL_FADD comp10_12 (
    .a(i10[12]),
    .b(sum_9[12]),
    .c(cout_10[11]),
    .cout(cout_10[12]),
    .sum(sum_10[12]));
  AL_FADD comp10_13 (
    .a(i10[13]),
    .b(sum_9[13]),
    .c(cout_10[12]),
    .cout(cout_10[13]),
    .sum(sum_10[13]));
  AL_FADD comp10_14 (
    .a(i10[14]),
    .b(sum_9[14]),
    .c(cout_10[13]),
    .cout(cout_10[14]),
    .sum(sum_10[14]));
  AL_FADD comp10_15 (
    .a(i10[15]),
    .b(sum_9[15]),
    .c(cout_10[14]),
    .cout(cout_10[15]),
    .sum(sum_10[15]));
  AL_FADD comp10_16 (
    .a(i10[16]),
    .b(sum_9[16]),
    .c(cout_10[15]),
    .cout(cout_10[16]),
    .sum(sum_10[16]));
  AL_FADD comp10_17 (
    .a(i10[17]),
    .b(sum_9[17]),
    .c(cout_10[16]),
    .cout(cout_10[17]),
    .sum(sum_10[17]));
  AL_FADD comp10_18 (
    .a(i10[18]),
    .b(sum_9[18]),
    .c(cout_10[17]),
    .cout(cout_10[18]),
    .sum(sum_10[18]));
  AL_FADD comp10_19 (
    .a(i10[19]),
    .b(sum_9[19]),
    .c(cout_10[18]),
    .cout(cout_10[19]),
    .sum(sum_10[19]));
  AL_FADD comp10_2 (
    .a(i10[2]),
    .b(sum_9[2]),
    .c(cout_10[1]),
    .cout(cout_10[2]),
    .sum(sum_10[2]));
  AL_FADD comp10_20 (
    .a(i10[20]),
    .b(sum_9[20]),
    .c(cout_10[19]),
    .cout(cout_10[20]),
    .sum(sum_10[20]));
  AL_FADD comp10_21 (
    .a(i10[21]),
    .b(sum_9[21]),
    .c(cout_10[20]),
    .cout(cout_10[21]),
    .sum(sum_10[21]));
  AL_FADD comp10_22 (
    .a(i10[22]),
    .b(sum_9[22]),
    .c(cout_10[21]),
    .cout(cout_10[22]),
    .sum(sum_10[22]));
  AL_FADD comp10_23 (
    .a(i10[23]),
    .b(sum_9[23]),
    .c(cout_10[22]),
    .cout(cout_10[23]),
    .sum(sum_10[23]));
  AL_FADD comp10_24 (
    .a(i10[24]),
    .b(sum_9[24]),
    .c(cout_10[23]),
    .cout(cout_10[24]),
    .sum(sum_10[24]));
  AL_FADD comp10_25 (
    .a(i10[25]),
    .b(sum_9[25]),
    .c(cout_10[24]),
    .cout(cout_10[25]),
    .sum(sum_10[25]));
  AL_FADD comp10_26 (
    .a(i10[26]),
    .b(sum_9[26]),
    .c(cout_10[25]),
    .cout(cout_10[26]),
    .sum(sum_10[26]));
  AL_FADD comp10_27 (
    .a(i10[27]),
    .b(sum_9[27]),
    .c(cout_10[26]),
    .cout(cout_10[27]),
    .sum(sum_10[27]));
  AL_FADD comp10_28 (
    .a(i10[28]),
    .b(sum_9[28]),
    .c(cout_10[27]),
    .cout(cout_10[28]),
    .sum(sum_10[28]));
  AL_FADD comp10_29 (
    .a(i10[29]),
    .b(sum_9[29]),
    .c(cout_10[28]),
    .cout(cout_10[29]),
    .sum(sum_10[29]));
  AL_FADD comp10_3 (
    .a(i10[3]),
    .b(sum_9[3]),
    .c(cout_10[2]),
    .cout(cout_10[3]),
    .sum(sum_10[3]));
  AL_FADD comp10_30 (
    .a(i10[30]),
    .b(sum_9[30]),
    .c(cout_10[29]),
    .cout(cout_10[30]),
    .sum(sum_10[30]));
  AL_FADD comp10_31 (
    .a(i10[31]),
    .b(sum_9[31]),
    .c(cout_10[30]),
    .cout(cout_10[31]),
    .sum(sum_10[31]));
  AL_FADD comp10_32 (
    .a(i10[32]),
    .b(sum_9[32]),
    .c(cout_10[31]),
    .cout(cout_10[32]),
    .sum(sum_10[32]));
  AL_FADD comp10_33 (
    .a(i10[33]),
    .b(sum_9[33]),
    .c(cout_10[32]),
    .cout(cout_10[33]),
    .sum(sum_10[33]));
  AL_FADD comp10_34 (
    .a(i10[34]),
    .b(sum_9[34]),
    .c(cout_10[33]),
    .cout(cout_10[34]),
    .sum(sum_10[34]));
  AL_FADD comp10_35 (
    .a(i10[35]),
    .b(sum_9[35]),
    .c(cout_10[34]),
    .cout(cout_10[35]),
    .sum(sum_10[35]));
  AL_FADD comp10_36 (
    .a(i10[36]),
    .b(sum_9[36]),
    .c(cout_10[35]),
    .cout(cout_10[36]),
    .sum(sum_10[36]));
  AL_FADD comp10_37 (
    .a(i10[37]),
    .b(sum_9[37]),
    .c(cout_10[36]),
    .cout(cout_10[37]),
    .sum(sum_10[37]));
  AL_FADD comp10_38 (
    .a(i10[38]),
    .b(sum_9[38]),
    .c(cout_10[37]),
    .cout(cout_10[38]),
    .sum(sum_10[38]));
  AL_FADD comp10_39 (
    .a(i10[39]),
    .b(sum_9[39]),
    .c(cout_10[38]),
    .cout(cout_10[39]),
    .sum(sum_10[39]));
  AL_FADD comp10_4 (
    .a(i10[4]),
    .b(sum_9[4]),
    .c(cout_10[3]),
    .cout(cout_10[4]),
    .sum(sum_10[4]));
  AL_FADD comp10_40 (
    .a(i10[40]),
    .b(sum_9[40]),
    .c(cout_10[39]),
    .cout(cout_10[40]),
    .sum(sum_10[40]));
  AL_FADD comp10_41 (
    .a(i10[41]),
    .b(sum_9[41]),
    .c(cout_10[40]),
    .cout(cout_10[41]),
    .sum(sum_10[41]));
  AL_FADD comp10_42 (
    .a(i10[42]),
    .b(sum_9[42]),
    .c(cout_10[41]),
    .cout(cout_10[42]),
    .sum(sum_10[42]));
  AL_FADD comp10_43 (
    .a(i10[43]),
    .b(sum_9[43]),
    .c(cout_10[42]),
    .cout(cout_10[43]),
    .sum(sum_10[43]));
  AL_FADD comp10_44 (
    .a(i10[44]),
    .b(sum_9[44]),
    .c(cout_10[43]),
    .cout(cout_10[44]),
    .sum(sum_10[44]));
  AL_FADD comp10_45 (
    .a(i10[45]),
    .b(sum_9[45]),
    .c(cout_10[44]),
    .cout(cout_10[45]),
    .sum(sum_10[45]));
  AL_FADD comp10_46 (
    .a(i10[46]),
    .b(sum_9[46]),
    .c(cout_10[45]),
    .cout(cout_10[46]),
    .sum(sum_10[46]));
  AL_FADD comp10_47 (
    .a(i10[47]),
    .b(sum_9[47]),
    .c(cout_10[46]),
    .cout(cout_10[47]),
    .sum(sum_10[47]));
  AL_FADD comp10_48 (
    .a(i10[48]),
    .b(sum_9[48]),
    .c(cout_10[47]),
    .cout(cout_10[48]),
    .sum(sum_10[48]));
  AL_FADD comp10_49 (
    .a(i10[49]),
    .b(sum_9[49]),
    .c(cout_10[48]),
    .cout(cout_10[49]),
    .sum(sum_10[49]));
  AL_FADD comp10_5 (
    .a(i10[5]),
    .b(sum_9[5]),
    .c(cout_10[4]),
    .cout(cout_10[5]),
    .sum(sum_10[5]));
  AL_FADD comp10_50 (
    .a(i10[50]),
    .b(sum_9[50]),
    .c(cout_10[49]),
    .cout(cout_10[50]),
    .sum(sum_10[50]));
  AL_FADD comp10_51 (
    .a(i10[51]),
    .b(sum_9[51]),
    .c(cout_10[50]),
    .cout(cout_10[51]),
    .sum(sum_10[51]));
  AL_FADD comp10_52 (
    .a(1'b0),
    .b(sum_9[52]),
    .c(cout_10[51]),
    .cout(cout_10[52]),
    .sum(sum_10[52]));
  AL_FADD comp10_53 (
    .a(1'b0),
    .b(sum_9[53]),
    .c(cout_10[52]),
    .cout(cout_10[53]),
    .sum(sum_10[53]));
  AL_FADD comp10_54 (
    .a(1'b0),
    .b(sum_9[54]),
    .c(cout_10[53]),
    .cout(cout_10[54]),
    .sum(sum_10[54]));
  AL_FADD comp10_55 (
    .a(1'b0),
    .b(sum_9[55]),
    .c(cout_10[54]),
    .cout(cout_10[55]),
    .sum(sum_10[55]));
  AL_FADD comp10_56 (
    .a(1'b0),
    .b(sum_9[56]),
    .c(cout_10[55]),
    .cout(cout_10[56]),
    .sum(sum_10[56]));
  AL_FADD comp10_57 (
    .a(1'b0),
    .b(sum_9[57]),
    .c(cout_10[56]),
    .cout(cout_10[57]),
    .sum(sum_10[57]));
  AL_FADD comp10_58 (
    .a(1'b0),
    .b(sum_9[58]),
    .c(cout_10[57]),
    .cout(cout_10[58]),
    .sum(sum_10[58]));
  AL_FADD comp10_59 (
    .a(1'b0),
    .b(sum_9[59]),
    .c(cout_10[58]),
    .cout(cout_10[59]),
    .sum(sum_10[59]));
  AL_FADD comp10_6 (
    .a(i10[6]),
    .b(sum_9[6]),
    .c(cout_10[5]),
    .cout(cout_10[6]),
    .sum(sum_10[6]));
  AL_FADD comp10_60 (
    .a(1'b0),
    .b(sum_9[60]),
    .c(cout_10[59]),
    .cout(cout_10[60]),
    .sum(sum_10[60]));
  AL_FADD comp10_61 (
    .a(1'b0),
    .b(sum_9[61]),
    .c(cout_10[60]),
    .cout(cout_10[61]),
    .sum(sum_10[61]));
  AL_FADD comp10_62 (
    .a(1'b0),
    .b(sum_9[62]),
    .c(cout_10[61]),
    .cout(cout_10[62]),
    .sum(sum_10[62]));
  AL_FADD comp10_63 (
    .a(1'b0),
    .b(sum_9[63]),
    .c(cout_10[62]),
    .cout(cout_10[63]),
    .sum(sum_10[63]));
  AL_FADD comp10_7 (
    .a(i10[7]),
    .b(sum_9[7]),
    .c(cout_10[6]),
    .cout(cout_10[7]),
    .sum(sum_10[7]));
  AL_FADD comp10_8 (
    .a(i10[8]),
    .b(sum_9[8]),
    .c(cout_10[7]),
    .cout(cout_10[8]),
    .sum(sum_10[8]));
  AL_FADD comp10_9 (
    .a(i10[9]),
    .b(sum_9[9]),
    .c(cout_10[8]),
    .cout(cout_10[9]),
    .sum(sum_10[9]));
  AL_FADD comp11_0 (
    .a(i11[0]),
    .b(sum_10[0]),
    .c(1'b0),
    .cout(cout_11[0]),
    .sum(sum_11[0]));
  AL_FADD comp11_1 (
    .a(i11[1]),
    .b(sum_10[1]),
    .c(cout_11[0]),
    .cout(cout_11[1]),
    .sum(sum_11[1]));
  AL_FADD comp11_10 (
    .a(i11[10]),
    .b(sum_10[10]),
    .c(cout_11[9]),
    .cout(cout_11[10]),
    .sum(sum_11[10]));
  AL_FADD comp11_11 (
    .a(i11[11]),
    .b(sum_10[11]),
    .c(cout_11[10]),
    .cout(cout_11[11]),
    .sum(sum_11[11]));
  AL_FADD comp11_12 (
    .a(i11[12]),
    .b(sum_10[12]),
    .c(cout_11[11]),
    .cout(cout_11[12]),
    .sum(sum_11[12]));
  AL_FADD comp11_13 (
    .a(i11[13]),
    .b(sum_10[13]),
    .c(cout_11[12]),
    .cout(cout_11[13]),
    .sum(sum_11[13]));
  AL_FADD comp11_14 (
    .a(i11[14]),
    .b(sum_10[14]),
    .c(cout_11[13]),
    .cout(cout_11[14]),
    .sum(sum_11[14]));
  AL_FADD comp11_15 (
    .a(i11[15]),
    .b(sum_10[15]),
    .c(cout_11[14]),
    .cout(cout_11[15]),
    .sum(sum_11[15]));
  AL_FADD comp11_16 (
    .a(i11[16]),
    .b(sum_10[16]),
    .c(cout_11[15]),
    .cout(cout_11[16]),
    .sum(sum_11[16]));
  AL_FADD comp11_17 (
    .a(i11[17]),
    .b(sum_10[17]),
    .c(cout_11[16]),
    .cout(cout_11[17]),
    .sum(sum_11[17]));
  AL_FADD comp11_18 (
    .a(i11[18]),
    .b(sum_10[18]),
    .c(cout_11[17]),
    .cout(cout_11[18]),
    .sum(sum_11[18]));
  AL_FADD comp11_19 (
    .a(i11[19]),
    .b(sum_10[19]),
    .c(cout_11[18]),
    .cout(cout_11[19]),
    .sum(sum_11[19]));
  AL_FADD comp11_2 (
    .a(i11[2]),
    .b(sum_10[2]),
    .c(cout_11[1]),
    .cout(cout_11[2]),
    .sum(sum_11[2]));
  AL_FADD comp11_20 (
    .a(i11[20]),
    .b(sum_10[20]),
    .c(cout_11[19]),
    .cout(cout_11[20]),
    .sum(sum_11[20]));
  AL_FADD comp11_21 (
    .a(i11[21]),
    .b(sum_10[21]),
    .c(cout_11[20]),
    .cout(cout_11[21]),
    .sum(sum_11[21]));
  AL_FADD comp11_22 (
    .a(i11[22]),
    .b(sum_10[22]),
    .c(cout_11[21]),
    .cout(cout_11[22]),
    .sum(sum_11[22]));
  AL_FADD comp11_23 (
    .a(i11[23]),
    .b(sum_10[23]),
    .c(cout_11[22]),
    .cout(cout_11[23]),
    .sum(sum_11[23]));
  AL_FADD comp11_24 (
    .a(i11[24]),
    .b(sum_10[24]),
    .c(cout_11[23]),
    .cout(cout_11[24]),
    .sum(sum_11[24]));
  AL_FADD comp11_25 (
    .a(i11[25]),
    .b(sum_10[25]),
    .c(cout_11[24]),
    .cout(cout_11[25]),
    .sum(sum_11[25]));
  AL_FADD comp11_26 (
    .a(i11[26]),
    .b(sum_10[26]),
    .c(cout_11[25]),
    .cout(cout_11[26]),
    .sum(sum_11[26]));
  AL_FADD comp11_27 (
    .a(i11[27]),
    .b(sum_10[27]),
    .c(cout_11[26]),
    .cout(cout_11[27]),
    .sum(sum_11[27]));
  AL_FADD comp11_28 (
    .a(i11[28]),
    .b(sum_10[28]),
    .c(cout_11[27]),
    .cout(cout_11[28]),
    .sum(sum_11[28]));
  AL_FADD comp11_29 (
    .a(i11[29]),
    .b(sum_10[29]),
    .c(cout_11[28]),
    .cout(cout_11[29]),
    .sum(sum_11[29]));
  AL_FADD comp11_3 (
    .a(i11[3]),
    .b(sum_10[3]),
    .c(cout_11[2]),
    .cout(cout_11[3]),
    .sum(sum_11[3]));
  AL_FADD comp11_30 (
    .a(i11[30]),
    .b(sum_10[30]),
    .c(cout_11[29]),
    .cout(cout_11[30]),
    .sum(sum_11[30]));
  AL_FADD comp11_31 (
    .a(i11[31]),
    .b(sum_10[31]),
    .c(cout_11[30]),
    .cout(cout_11[31]),
    .sum(sum_11[31]));
  AL_FADD comp11_32 (
    .a(i11[32]),
    .b(sum_10[32]),
    .c(cout_11[31]),
    .cout(cout_11[32]),
    .sum(sum_11[32]));
  AL_FADD comp11_33 (
    .a(i11[33]),
    .b(sum_10[33]),
    .c(cout_11[32]),
    .cout(cout_11[33]),
    .sum(sum_11[33]));
  AL_FADD comp11_34 (
    .a(i11[34]),
    .b(sum_10[34]),
    .c(cout_11[33]),
    .cout(cout_11[34]),
    .sum(sum_11[34]));
  AL_FADD comp11_35 (
    .a(i11[35]),
    .b(sum_10[35]),
    .c(cout_11[34]),
    .cout(cout_11[35]),
    .sum(sum_11[35]));
  AL_FADD comp11_36 (
    .a(i11[36]),
    .b(sum_10[36]),
    .c(cout_11[35]),
    .cout(cout_11[36]),
    .sum(sum_11[36]));
  AL_FADD comp11_37 (
    .a(i11[37]),
    .b(sum_10[37]),
    .c(cout_11[36]),
    .cout(cout_11[37]),
    .sum(sum_11[37]));
  AL_FADD comp11_38 (
    .a(i11[38]),
    .b(sum_10[38]),
    .c(cout_11[37]),
    .cout(cout_11[38]),
    .sum(sum_11[38]));
  AL_FADD comp11_39 (
    .a(i11[39]),
    .b(sum_10[39]),
    .c(cout_11[38]),
    .cout(cout_11[39]),
    .sum(sum_11[39]));
  AL_FADD comp11_4 (
    .a(i11[4]),
    .b(sum_10[4]),
    .c(cout_11[3]),
    .cout(cout_11[4]),
    .sum(sum_11[4]));
  AL_FADD comp11_40 (
    .a(i11[40]),
    .b(sum_10[40]),
    .c(cout_11[39]),
    .cout(cout_11[40]),
    .sum(sum_11[40]));
  AL_FADD comp11_41 (
    .a(i11[41]),
    .b(sum_10[41]),
    .c(cout_11[40]),
    .cout(cout_11[41]),
    .sum(sum_11[41]));
  AL_FADD comp11_42 (
    .a(i11[42]),
    .b(sum_10[42]),
    .c(cout_11[41]),
    .cout(cout_11[42]),
    .sum(sum_11[42]));
  AL_FADD comp11_43 (
    .a(i11[43]),
    .b(sum_10[43]),
    .c(cout_11[42]),
    .cout(cout_11[43]),
    .sum(sum_11[43]));
  AL_FADD comp11_44 (
    .a(i11[44]),
    .b(sum_10[44]),
    .c(cout_11[43]),
    .cout(cout_11[44]),
    .sum(sum_11[44]));
  AL_FADD comp11_45 (
    .a(i11[45]),
    .b(sum_10[45]),
    .c(cout_11[44]),
    .cout(cout_11[45]),
    .sum(sum_11[45]));
  AL_FADD comp11_46 (
    .a(i11[46]),
    .b(sum_10[46]),
    .c(cout_11[45]),
    .cout(cout_11[46]),
    .sum(sum_11[46]));
  AL_FADD comp11_47 (
    .a(i11[47]),
    .b(sum_10[47]),
    .c(cout_11[46]),
    .cout(cout_11[47]),
    .sum(sum_11[47]));
  AL_FADD comp11_48 (
    .a(i11[48]),
    .b(sum_10[48]),
    .c(cout_11[47]),
    .cout(cout_11[48]),
    .sum(sum_11[48]));
  AL_FADD comp11_49 (
    .a(i11[49]),
    .b(sum_10[49]),
    .c(cout_11[48]),
    .cout(cout_11[49]),
    .sum(sum_11[49]));
  AL_FADD comp11_5 (
    .a(i11[5]),
    .b(sum_10[5]),
    .c(cout_11[4]),
    .cout(cout_11[5]),
    .sum(sum_11[5]));
  AL_FADD comp11_50 (
    .a(i11[50]),
    .b(sum_10[50]),
    .c(cout_11[49]),
    .cout(cout_11[50]),
    .sum(sum_11[50]));
  AL_FADD comp11_51 (
    .a(1'b0),
    .b(sum_10[51]),
    .c(cout_11[50]),
    .cout(cout_11[51]),
    .sum(sum_11[51]));
  AL_FADD comp11_52 (
    .a(1'b0),
    .b(sum_10[52]),
    .c(cout_11[51]),
    .cout(cout_11[52]),
    .sum(sum_11[52]));
  AL_FADD comp11_53 (
    .a(1'b0),
    .b(sum_10[53]),
    .c(cout_11[52]),
    .cout(cout_11[53]),
    .sum(sum_11[53]));
  AL_FADD comp11_54 (
    .a(1'b0),
    .b(sum_10[54]),
    .c(cout_11[53]),
    .cout(cout_11[54]),
    .sum(sum_11[54]));
  AL_FADD comp11_55 (
    .a(1'b0),
    .b(sum_10[55]),
    .c(cout_11[54]),
    .cout(cout_11[55]),
    .sum(sum_11[55]));
  AL_FADD comp11_56 (
    .a(1'b0),
    .b(sum_10[56]),
    .c(cout_11[55]),
    .cout(cout_11[56]),
    .sum(sum_11[56]));
  AL_FADD comp11_57 (
    .a(1'b0),
    .b(sum_10[57]),
    .c(cout_11[56]),
    .cout(cout_11[57]),
    .sum(sum_11[57]));
  AL_FADD comp11_58 (
    .a(1'b0),
    .b(sum_10[58]),
    .c(cout_11[57]),
    .cout(cout_11[58]),
    .sum(sum_11[58]));
  AL_FADD comp11_59 (
    .a(1'b0),
    .b(sum_10[59]),
    .c(cout_11[58]),
    .cout(cout_11[59]),
    .sum(sum_11[59]));
  AL_FADD comp11_6 (
    .a(i11[6]),
    .b(sum_10[6]),
    .c(cout_11[5]),
    .cout(cout_11[6]),
    .sum(sum_11[6]));
  AL_FADD comp11_60 (
    .a(1'b0),
    .b(sum_10[60]),
    .c(cout_11[59]),
    .cout(cout_11[60]),
    .sum(sum_11[60]));
  AL_FADD comp11_61 (
    .a(1'b0),
    .b(sum_10[61]),
    .c(cout_11[60]),
    .cout(cout_11[61]),
    .sum(sum_11[61]));
  AL_FADD comp11_62 (
    .a(1'b0),
    .b(sum_10[62]),
    .c(cout_11[61]),
    .cout(cout_11[62]),
    .sum(sum_11[62]));
  AL_FADD comp11_63 (
    .a(1'b0),
    .b(sum_10[63]),
    .c(cout_11[62]),
    .cout(cout_11[63]),
    .sum(sum_11[63]));
  AL_FADD comp11_7 (
    .a(i11[7]),
    .b(sum_10[7]),
    .c(cout_11[6]),
    .cout(cout_11[7]),
    .sum(sum_11[7]));
  AL_FADD comp11_8 (
    .a(i11[8]),
    .b(sum_10[8]),
    .c(cout_11[7]),
    .cout(cout_11[8]),
    .sum(sum_11[8]));
  AL_FADD comp11_9 (
    .a(i11[9]),
    .b(sum_10[9]),
    .c(cout_11[8]),
    .cout(cout_11[9]),
    .sum(sum_11[9]));
  AL_FADD comp12_0 (
    .a(i12[0]),
    .b(sum_11[0]),
    .c(1'b0),
    .cout(cout_12[0]),
    .sum(sum_12[0]));
  AL_FADD comp12_1 (
    .a(i12[1]),
    .b(sum_11[1]),
    .c(cout_12[0]),
    .cout(cout_12[1]),
    .sum(sum_12[1]));
  AL_FADD comp12_10 (
    .a(i12[10]),
    .b(sum_11[10]),
    .c(cout_12[9]),
    .cout(cout_12[10]),
    .sum(sum_12[10]));
  AL_FADD comp12_11 (
    .a(i12[11]),
    .b(sum_11[11]),
    .c(cout_12[10]),
    .cout(cout_12[11]),
    .sum(sum_12[11]));
  AL_FADD comp12_12 (
    .a(i12[12]),
    .b(sum_11[12]),
    .c(cout_12[11]),
    .cout(cout_12[12]),
    .sum(sum_12[12]));
  AL_FADD comp12_13 (
    .a(i12[13]),
    .b(sum_11[13]),
    .c(cout_12[12]),
    .cout(cout_12[13]),
    .sum(sum_12[13]));
  AL_FADD comp12_14 (
    .a(i12[14]),
    .b(sum_11[14]),
    .c(cout_12[13]),
    .cout(cout_12[14]),
    .sum(sum_12[14]));
  AL_FADD comp12_15 (
    .a(i12[15]),
    .b(sum_11[15]),
    .c(cout_12[14]),
    .cout(cout_12[15]),
    .sum(sum_12[15]));
  AL_FADD comp12_16 (
    .a(i12[16]),
    .b(sum_11[16]),
    .c(cout_12[15]),
    .cout(cout_12[16]),
    .sum(sum_12[16]));
  AL_FADD comp12_17 (
    .a(i12[17]),
    .b(sum_11[17]),
    .c(cout_12[16]),
    .cout(cout_12[17]),
    .sum(sum_12[17]));
  AL_FADD comp12_18 (
    .a(i12[18]),
    .b(sum_11[18]),
    .c(cout_12[17]),
    .cout(cout_12[18]),
    .sum(sum_12[18]));
  AL_FADD comp12_19 (
    .a(i12[19]),
    .b(sum_11[19]),
    .c(cout_12[18]),
    .cout(cout_12[19]),
    .sum(sum_12[19]));
  AL_FADD comp12_2 (
    .a(i12[2]),
    .b(sum_11[2]),
    .c(cout_12[1]),
    .cout(cout_12[2]),
    .sum(sum_12[2]));
  AL_FADD comp12_20 (
    .a(i12[20]),
    .b(sum_11[20]),
    .c(cout_12[19]),
    .cout(cout_12[20]),
    .sum(sum_12[20]));
  AL_FADD comp12_21 (
    .a(i12[21]),
    .b(sum_11[21]),
    .c(cout_12[20]),
    .cout(cout_12[21]),
    .sum(sum_12[21]));
  AL_FADD comp12_22 (
    .a(i12[22]),
    .b(sum_11[22]),
    .c(cout_12[21]),
    .cout(cout_12[22]),
    .sum(sum_12[22]));
  AL_FADD comp12_23 (
    .a(i12[23]),
    .b(sum_11[23]),
    .c(cout_12[22]),
    .cout(cout_12[23]),
    .sum(sum_12[23]));
  AL_FADD comp12_24 (
    .a(i12[24]),
    .b(sum_11[24]),
    .c(cout_12[23]),
    .cout(cout_12[24]),
    .sum(sum_12[24]));
  AL_FADD comp12_25 (
    .a(i12[25]),
    .b(sum_11[25]),
    .c(cout_12[24]),
    .cout(cout_12[25]),
    .sum(sum_12[25]));
  AL_FADD comp12_26 (
    .a(i12[26]),
    .b(sum_11[26]),
    .c(cout_12[25]),
    .cout(cout_12[26]),
    .sum(sum_12[26]));
  AL_FADD comp12_27 (
    .a(i12[27]),
    .b(sum_11[27]),
    .c(cout_12[26]),
    .cout(cout_12[27]),
    .sum(sum_12[27]));
  AL_FADD comp12_28 (
    .a(i12[28]),
    .b(sum_11[28]),
    .c(cout_12[27]),
    .cout(cout_12[28]),
    .sum(sum_12[28]));
  AL_FADD comp12_29 (
    .a(i12[29]),
    .b(sum_11[29]),
    .c(cout_12[28]),
    .cout(cout_12[29]),
    .sum(sum_12[29]));
  AL_FADD comp12_3 (
    .a(i12[3]),
    .b(sum_11[3]),
    .c(cout_12[2]),
    .cout(cout_12[3]),
    .sum(sum_12[3]));
  AL_FADD comp12_30 (
    .a(i12[30]),
    .b(sum_11[30]),
    .c(cout_12[29]),
    .cout(cout_12[30]),
    .sum(sum_12[30]));
  AL_FADD comp12_31 (
    .a(i12[31]),
    .b(sum_11[31]),
    .c(cout_12[30]),
    .cout(cout_12[31]),
    .sum(sum_12[31]));
  AL_FADD comp12_32 (
    .a(i12[32]),
    .b(sum_11[32]),
    .c(cout_12[31]),
    .cout(cout_12[32]),
    .sum(sum_12[32]));
  AL_FADD comp12_33 (
    .a(i12[33]),
    .b(sum_11[33]),
    .c(cout_12[32]),
    .cout(cout_12[33]),
    .sum(sum_12[33]));
  AL_FADD comp12_34 (
    .a(i12[34]),
    .b(sum_11[34]),
    .c(cout_12[33]),
    .cout(cout_12[34]),
    .sum(sum_12[34]));
  AL_FADD comp12_35 (
    .a(i12[35]),
    .b(sum_11[35]),
    .c(cout_12[34]),
    .cout(cout_12[35]),
    .sum(sum_12[35]));
  AL_FADD comp12_36 (
    .a(i12[36]),
    .b(sum_11[36]),
    .c(cout_12[35]),
    .cout(cout_12[36]),
    .sum(sum_12[36]));
  AL_FADD comp12_37 (
    .a(i12[37]),
    .b(sum_11[37]),
    .c(cout_12[36]),
    .cout(cout_12[37]),
    .sum(sum_12[37]));
  AL_FADD comp12_38 (
    .a(i12[38]),
    .b(sum_11[38]),
    .c(cout_12[37]),
    .cout(cout_12[38]),
    .sum(sum_12[38]));
  AL_FADD comp12_39 (
    .a(i12[39]),
    .b(sum_11[39]),
    .c(cout_12[38]),
    .cout(cout_12[39]),
    .sum(sum_12[39]));
  AL_FADD comp12_4 (
    .a(i12[4]),
    .b(sum_11[4]),
    .c(cout_12[3]),
    .cout(cout_12[4]),
    .sum(sum_12[4]));
  AL_FADD comp12_40 (
    .a(i12[40]),
    .b(sum_11[40]),
    .c(cout_12[39]),
    .cout(cout_12[40]),
    .sum(sum_12[40]));
  AL_FADD comp12_41 (
    .a(i12[41]),
    .b(sum_11[41]),
    .c(cout_12[40]),
    .cout(cout_12[41]),
    .sum(sum_12[41]));
  AL_FADD comp12_42 (
    .a(i12[42]),
    .b(sum_11[42]),
    .c(cout_12[41]),
    .cout(cout_12[42]),
    .sum(sum_12[42]));
  AL_FADD comp12_43 (
    .a(i12[43]),
    .b(sum_11[43]),
    .c(cout_12[42]),
    .cout(cout_12[43]),
    .sum(sum_12[43]));
  AL_FADD comp12_44 (
    .a(i12[44]),
    .b(sum_11[44]),
    .c(cout_12[43]),
    .cout(cout_12[44]),
    .sum(sum_12[44]));
  AL_FADD comp12_45 (
    .a(i12[45]),
    .b(sum_11[45]),
    .c(cout_12[44]),
    .cout(cout_12[45]),
    .sum(sum_12[45]));
  AL_FADD comp12_46 (
    .a(i12[46]),
    .b(sum_11[46]),
    .c(cout_12[45]),
    .cout(cout_12[46]),
    .sum(sum_12[46]));
  AL_FADD comp12_47 (
    .a(i12[47]),
    .b(sum_11[47]),
    .c(cout_12[46]),
    .cout(cout_12[47]),
    .sum(sum_12[47]));
  AL_FADD comp12_48 (
    .a(i12[48]),
    .b(sum_11[48]),
    .c(cout_12[47]),
    .cout(cout_12[48]),
    .sum(sum_12[48]));
  AL_FADD comp12_49 (
    .a(i12[49]),
    .b(sum_11[49]),
    .c(cout_12[48]),
    .cout(cout_12[49]),
    .sum(sum_12[49]));
  AL_FADD comp12_5 (
    .a(i12[5]),
    .b(sum_11[5]),
    .c(cout_12[4]),
    .cout(cout_12[5]),
    .sum(sum_12[5]));
  AL_FADD comp12_50 (
    .a(1'b0),
    .b(sum_11[50]),
    .c(cout_12[49]),
    .cout(cout_12[50]),
    .sum(sum_12[50]));
  AL_FADD comp12_51 (
    .a(1'b0),
    .b(sum_11[51]),
    .c(cout_12[50]),
    .cout(cout_12[51]),
    .sum(sum_12[51]));
  AL_FADD comp12_52 (
    .a(1'b0),
    .b(sum_11[52]),
    .c(cout_12[51]),
    .cout(cout_12[52]),
    .sum(sum_12[52]));
  AL_FADD comp12_53 (
    .a(1'b0),
    .b(sum_11[53]),
    .c(cout_12[52]),
    .cout(cout_12[53]),
    .sum(sum_12[53]));
  AL_FADD comp12_54 (
    .a(1'b0),
    .b(sum_11[54]),
    .c(cout_12[53]),
    .cout(cout_12[54]),
    .sum(sum_12[54]));
  AL_FADD comp12_55 (
    .a(1'b0),
    .b(sum_11[55]),
    .c(cout_12[54]),
    .cout(cout_12[55]),
    .sum(sum_12[55]));
  AL_FADD comp12_56 (
    .a(1'b0),
    .b(sum_11[56]),
    .c(cout_12[55]),
    .cout(cout_12[56]),
    .sum(sum_12[56]));
  AL_FADD comp12_57 (
    .a(1'b0),
    .b(sum_11[57]),
    .c(cout_12[56]),
    .cout(cout_12[57]),
    .sum(sum_12[57]));
  AL_FADD comp12_58 (
    .a(1'b0),
    .b(sum_11[58]),
    .c(cout_12[57]),
    .cout(cout_12[58]),
    .sum(sum_12[58]));
  AL_FADD comp12_59 (
    .a(1'b0),
    .b(sum_11[59]),
    .c(cout_12[58]),
    .cout(cout_12[59]),
    .sum(sum_12[59]));
  AL_FADD comp12_6 (
    .a(i12[6]),
    .b(sum_11[6]),
    .c(cout_12[5]),
    .cout(cout_12[6]),
    .sum(sum_12[6]));
  AL_FADD comp12_60 (
    .a(1'b0),
    .b(sum_11[60]),
    .c(cout_12[59]),
    .cout(cout_12[60]),
    .sum(sum_12[60]));
  AL_FADD comp12_61 (
    .a(1'b0),
    .b(sum_11[61]),
    .c(cout_12[60]),
    .cout(cout_12[61]),
    .sum(sum_12[61]));
  AL_FADD comp12_62 (
    .a(1'b0),
    .b(sum_11[62]),
    .c(cout_12[61]),
    .cout(cout_12[62]),
    .sum(sum_12[62]));
  AL_FADD comp12_63 (
    .a(1'b0),
    .b(sum_11[63]),
    .c(cout_12[62]),
    .cout(cout_12[63]),
    .sum(sum_12[63]));
  AL_FADD comp12_7 (
    .a(i12[7]),
    .b(sum_11[7]),
    .c(cout_12[6]),
    .cout(cout_12[7]),
    .sum(sum_12[7]));
  AL_FADD comp12_8 (
    .a(i12[8]),
    .b(sum_11[8]),
    .c(cout_12[7]),
    .cout(cout_12[8]),
    .sum(sum_12[8]));
  AL_FADD comp12_9 (
    .a(i12[9]),
    .b(sum_11[9]),
    .c(cout_12[8]),
    .cout(cout_12[9]),
    .sum(sum_12[9]));
  AL_FADD comp13_0 (
    .a(i13[0]),
    .b(sum_12[0]),
    .c(1'b0),
    .cout(cout_13[0]),
    .sum(sum_13[0]));
  AL_FADD comp13_1 (
    .a(i13[1]),
    .b(sum_12[1]),
    .c(cout_13[0]),
    .cout(cout_13[1]),
    .sum(sum_13[1]));
  AL_FADD comp13_10 (
    .a(i13[10]),
    .b(sum_12[10]),
    .c(cout_13[9]),
    .cout(cout_13[10]),
    .sum(sum_13[10]));
  AL_FADD comp13_11 (
    .a(i13[11]),
    .b(sum_12[11]),
    .c(cout_13[10]),
    .cout(cout_13[11]),
    .sum(sum_13[11]));
  AL_FADD comp13_12 (
    .a(i13[12]),
    .b(sum_12[12]),
    .c(cout_13[11]),
    .cout(cout_13[12]),
    .sum(sum_13[12]));
  AL_FADD comp13_13 (
    .a(i13[13]),
    .b(sum_12[13]),
    .c(cout_13[12]),
    .cout(cout_13[13]),
    .sum(sum_13[13]));
  AL_FADD comp13_14 (
    .a(i13[14]),
    .b(sum_12[14]),
    .c(cout_13[13]),
    .cout(cout_13[14]),
    .sum(sum_13[14]));
  AL_FADD comp13_15 (
    .a(i13[15]),
    .b(sum_12[15]),
    .c(cout_13[14]),
    .cout(cout_13[15]),
    .sum(sum_13[15]));
  AL_FADD comp13_16 (
    .a(i13[16]),
    .b(sum_12[16]),
    .c(cout_13[15]),
    .cout(cout_13[16]),
    .sum(sum_13[16]));
  AL_FADD comp13_17 (
    .a(i13[17]),
    .b(sum_12[17]),
    .c(cout_13[16]),
    .cout(cout_13[17]),
    .sum(sum_13[17]));
  AL_FADD comp13_18 (
    .a(i13[18]),
    .b(sum_12[18]),
    .c(cout_13[17]),
    .cout(cout_13[18]),
    .sum(sum_13[18]));
  AL_FADD comp13_19 (
    .a(i13[19]),
    .b(sum_12[19]),
    .c(cout_13[18]),
    .cout(cout_13[19]),
    .sum(sum_13[19]));
  AL_FADD comp13_2 (
    .a(i13[2]),
    .b(sum_12[2]),
    .c(cout_13[1]),
    .cout(cout_13[2]),
    .sum(sum_13[2]));
  AL_FADD comp13_20 (
    .a(i13[20]),
    .b(sum_12[20]),
    .c(cout_13[19]),
    .cout(cout_13[20]),
    .sum(sum_13[20]));
  AL_FADD comp13_21 (
    .a(i13[21]),
    .b(sum_12[21]),
    .c(cout_13[20]),
    .cout(cout_13[21]),
    .sum(sum_13[21]));
  AL_FADD comp13_22 (
    .a(i13[22]),
    .b(sum_12[22]),
    .c(cout_13[21]),
    .cout(cout_13[22]),
    .sum(sum_13[22]));
  AL_FADD comp13_23 (
    .a(i13[23]),
    .b(sum_12[23]),
    .c(cout_13[22]),
    .cout(cout_13[23]),
    .sum(sum_13[23]));
  AL_FADD comp13_24 (
    .a(i13[24]),
    .b(sum_12[24]),
    .c(cout_13[23]),
    .cout(cout_13[24]),
    .sum(sum_13[24]));
  AL_FADD comp13_25 (
    .a(i13[25]),
    .b(sum_12[25]),
    .c(cout_13[24]),
    .cout(cout_13[25]),
    .sum(sum_13[25]));
  AL_FADD comp13_26 (
    .a(i13[26]),
    .b(sum_12[26]),
    .c(cout_13[25]),
    .cout(cout_13[26]),
    .sum(sum_13[26]));
  AL_FADD comp13_27 (
    .a(i13[27]),
    .b(sum_12[27]),
    .c(cout_13[26]),
    .cout(cout_13[27]),
    .sum(sum_13[27]));
  AL_FADD comp13_28 (
    .a(i13[28]),
    .b(sum_12[28]),
    .c(cout_13[27]),
    .cout(cout_13[28]),
    .sum(sum_13[28]));
  AL_FADD comp13_29 (
    .a(i13[29]),
    .b(sum_12[29]),
    .c(cout_13[28]),
    .cout(cout_13[29]),
    .sum(sum_13[29]));
  AL_FADD comp13_3 (
    .a(i13[3]),
    .b(sum_12[3]),
    .c(cout_13[2]),
    .cout(cout_13[3]),
    .sum(sum_13[3]));
  AL_FADD comp13_30 (
    .a(i13[30]),
    .b(sum_12[30]),
    .c(cout_13[29]),
    .cout(cout_13[30]),
    .sum(sum_13[30]));
  AL_FADD comp13_31 (
    .a(i13[31]),
    .b(sum_12[31]),
    .c(cout_13[30]),
    .cout(cout_13[31]),
    .sum(sum_13[31]));
  AL_FADD comp13_32 (
    .a(i13[32]),
    .b(sum_12[32]),
    .c(cout_13[31]),
    .cout(cout_13[32]),
    .sum(sum_13[32]));
  AL_FADD comp13_33 (
    .a(i13[33]),
    .b(sum_12[33]),
    .c(cout_13[32]),
    .cout(cout_13[33]),
    .sum(sum_13[33]));
  AL_FADD comp13_34 (
    .a(i13[34]),
    .b(sum_12[34]),
    .c(cout_13[33]),
    .cout(cout_13[34]),
    .sum(sum_13[34]));
  AL_FADD comp13_35 (
    .a(i13[35]),
    .b(sum_12[35]),
    .c(cout_13[34]),
    .cout(cout_13[35]),
    .sum(sum_13[35]));
  AL_FADD comp13_36 (
    .a(i13[36]),
    .b(sum_12[36]),
    .c(cout_13[35]),
    .cout(cout_13[36]),
    .sum(sum_13[36]));
  AL_FADD comp13_37 (
    .a(i13[37]),
    .b(sum_12[37]),
    .c(cout_13[36]),
    .cout(cout_13[37]),
    .sum(sum_13[37]));
  AL_FADD comp13_38 (
    .a(i13[38]),
    .b(sum_12[38]),
    .c(cout_13[37]),
    .cout(cout_13[38]),
    .sum(sum_13[38]));
  AL_FADD comp13_39 (
    .a(i13[39]),
    .b(sum_12[39]),
    .c(cout_13[38]),
    .cout(cout_13[39]),
    .sum(sum_13[39]));
  AL_FADD comp13_4 (
    .a(i13[4]),
    .b(sum_12[4]),
    .c(cout_13[3]),
    .cout(cout_13[4]),
    .sum(sum_13[4]));
  AL_FADD comp13_40 (
    .a(i13[40]),
    .b(sum_12[40]),
    .c(cout_13[39]),
    .cout(cout_13[40]),
    .sum(sum_13[40]));
  AL_FADD comp13_41 (
    .a(i13[41]),
    .b(sum_12[41]),
    .c(cout_13[40]),
    .cout(cout_13[41]),
    .sum(sum_13[41]));
  AL_FADD comp13_42 (
    .a(i13[42]),
    .b(sum_12[42]),
    .c(cout_13[41]),
    .cout(cout_13[42]),
    .sum(sum_13[42]));
  AL_FADD comp13_43 (
    .a(i13[43]),
    .b(sum_12[43]),
    .c(cout_13[42]),
    .cout(cout_13[43]),
    .sum(sum_13[43]));
  AL_FADD comp13_44 (
    .a(i13[44]),
    .b(sum_12[44]),
    .c(cout_13[43]),
    .cout(cout_13[44]),
    .sum(sum_13[44]));
  AL_FADD comp13_45 (
    .a(i13[45]),
    .b(sum_12[45]),
    .c(cout_13[44]),
    .cout(cout_13[45]),
    .sum(sum_13[45]));
  AL_FADD comp13_46 (
    .a(i13[46]),
    .b(sum_12[46]),
    .c(cout_13[45]),
    .cout(cout_13[46]),
    .sum(sum_13[46]));
  AL_FADD comp13_47 (
    .a(i13[47]),
    .b(sum_12[47]),
    .c(cout_13[46]),
    .cout(cout_13[47]),
    .sum(sum_13[47]));
  AL_FADD comp13_48 (
    .a(i13[48]),
    .b(sum_12[48]),
    .c(cout_13[47]),
    .cout(cout_13[48]),
    .sum(sum_13[48]));
  AL_FADD comp13_49 (
    .a(1'b0),
    .b(sum_12[49]),
    .c(cout_13[48]),
    .cout(cout_13[49]),
    .sum(sum_13[49]));
  AL_FADD comp13_5 (
    .a(i13[5]),
    .b(sum_12[5]),
    .c(cout_13[4]),
    .cout(cout_13[5]),
    .sum(sum_13[5]));
  AL_FADD comp13_50 (
    .a(1'b0),
    .b(sum_12[50]),
    .c(cout_13[49]),
    .cout(cout_13[50]),
    .sum(sum_13[50]));
  AL_FADD comp13_51 (
    .a(1'b0),
    .b(sum_12[51]),
    .c(cout_13[50]),
    .cout(cout_13[51]),
    .sum(sum_13[51]));
  AL_FADD comp13_52 (
    .a(1'b0),
    .b(sum_12[52]),
    .c(cout_13[51]),
    .cout(cout_13[52]),
    .sum(sum_13[52]));
  AL_FADD comp13_53 (
    .a(1'b0),
    .b(sum_12[53]),
    .c(cout_13[52]),
    .cout(cout_13[53]),
    .sum(sum_13[53]));
  AL_FADD comp13_54 (
    .a(1'b0),
    .b(sum_12[54]),
    .c(cout_13[53]),
    .cout(cout_13[54]),
    .sum(sum_13[54]));
  AL_FADD comp13_55 (
    .a(1'b0),
    .b(sum_12[55]),
    .c(cout_13[54]),
    .cout(cout_13[55]),
    .sum(sum_13[55]));
  AL_FADD comp13_56 (
    .a(1'b0),
    .b(sum_12[56]),
    .c(cout_13[55]),
    .cout(cout_13[56]),
    .sum(sum_13[56]));
  AL_FADD comp13_57 (
    .a(1'b0),
    .b(sum_12[57]),
    .c(cout_13[56]),
    .cout(cout_13[57]),
    .sum(sum_13[57]));
  AL_FADD comp13_58 (
    .a(1'b0),
    .b(sum_12[58]),
    .c(cout_13[57]),
    .cout(cout_13[58]),
    .sum(sum_13[58]));
  AL_FADD comp13_59 (
    .a(1'b0),
    .b(sum_12[59]),
    .c(cout_13[58]),
    .cout(cout_13[59]),
    .sum(sum_13[59]));
  AL_FADD comp13_6 (
    .a(i13[6]),
    .b(sum_12[6]),
    .c(cout_13[5]),
    .cout(cout_13[6]),
    .sum(sum_13[6]));
  AL_FADD comp13_60 (
    .a(1'b0),
    .b(sum_12[60]),
    .c(cout_13[59]),
    .cout(cout_13[60]),
    .sum(sum_13[60]));
  AL_FADD comp13_61 (
    .a(1'b0),
    .b(sum_12[61]),
    .c(cout_13[60]),
    .cout(cout_13[61]),
    .sum(sum_13[61]));
  AL_FADD comp13_62 (
    .a(1'b0),
    .b(sum_12[62]),
    .c(cout_13[61]),
    .cout(cout_13[62]),
    .sum(sum_13[62]));
  AL_FADD comp13_63 (
    .a(1'b0),
    .b(sum_12[63]),
    .c(cout_13[62]),
    .cout(cout_13[63]),
    .sum(sum_13[63]));
  AL_FADD comp13_7 (
    .a(i13[7]),
    .b(sum_12[7]),
    .c(cout_13[6]),
    .cout(cout_13[7]),
    .sum(sum_13[7]));
  AL_FADD comp13_8 (
    .a(i13[8]),
    .b(sum_12[8]),
    .c(cout_13[7]),
    .cout(cout_13[8]),
    .sum(sum_13[8]));
  AL_FADD comp13_9 (
    .a(i13[9]),
    .b(sum_12[9]),
    .c(cout_13[8]),
    .cout(cout_13[9]),
    .sum(sum_13[9]));
  AL_FADD comp14_0 (
    .a(i14[0]),
    .b(sum_13[0]),
    .c(1'b0),
    .cout(cout_14[0]),
    .sum(sum_14[0]));
  AL_FADD comp14_1 (
    .a(i14[1]),
    .b(sum_13[1]),
    .c(cout_14[0]),
    .cout(cout_14[1]),
    .sum(sum_14[1]));
  AL_FADD comp14_10 (
    .a(i14[10]),
    .b(sum_13[10]),
    .c(cout_14[9]),
    .cout(cout_14[10]),
    .sum(sum_14[10]));
  AL_FADD comp14_11 (
    .a(i14[11]),
    .b(sum_13[11]),
    .c(cout_14[10]),
    .cout(cout_14[11]),
    .sum(sum_14[11]));
  AL_FADD comp14_12 (
    .a(i14[12]),
    .b(sum_13[12]),
    .c(cout_14[11]),
    .cout(cout_14[12]),
    .sum(sum_14[12]));
  AL_FADD comp14_13 (
    .a(i14[13]),
    .b(sum_13[13]),
    .c(cout_14[12]),
    .cout(cout_14[13]),
    .sum(sum_14[13]));
  AL_FADD comp14_14 (
    .a(i14[14]),
    .b(sum_13[14]),
    .c(cout_14[13]),
    .cout(cout_14[14]),
    .sum(sum_14[14]));
  AL_FADD comp14_15 (
    .a(i14[15]),
    .b(sum_13[15]),
    .c(cout_14[14]),
    .cout(cout_14[15]),
    .sum(sum_14[15]));
  AL_FADD comp14_16 (
    .a(i14[16]),
    .b(sum_13[16]),
    .c(cout_14[15]),
    .cout(cout_14[16]),
    .sum(sum_14[16]));
  AL_FADD comp14_17 (
    .a(i14[17]),
    .b(sum_13[17]),
    .c(cout_14[16]),
    .cout(cout_14[17]),
    .sum(sum_14[17]));
  AL_FADD comp14_18 (
    .a(i14[18]),
    .b(sum_13[18]),
    .c(cout_14[17]),
    .cout(cout_14[18]),
    .sum(sum_14[18]));
  AL_FADD comp14_19 (
    .a(i14[19]),
    .b(sum_13[19]),
    .c(cout_14[18]),
    .cout(cout_14[19]),
    .sum(sum_14[19]));
  AL_FADD comp14_2 (
    .a(i14[2]),
    .b(sum_13[2]),
    .c(cout_14[1]),
    .cout(cout_14[2]),
    .sum(sum_14[2]));
  AL_FADD comp14_20 (
    .a(i14[20]),
    .b(sum_13[20]),
    .c(cout_14[19]),
    .cout(cout_14[20]),
    .sum(sum_14[20]));
  AL_FADD comp14_21 (
    .a(i14[21]),
    .b(sum_13[21]),
    .c(cout_14[20]),
    .cout(cout_14[21]),
    .sum(sum_14[21]));
  AL_FADD comp14_22 (
    .a(i14[22]),
    .b(sum_13[22]),
    .c(cout_14[21]),
    .cout(cout_14[22]),
    .sum(sum_14[22]));
  AL_FADD comp14_23 (
    .a(i14[23]),
    .b(sum_13[23]),
    .c(cout_14[22]),
    .cout(cout_14[23]),
    .sum(sum_14[23]));
  AL_FADD comp14_24 (
    .a(i14[24]),
    .b(sum_13[24]),
    .c(cout_14[23]),
    .cout(cout_14[24]),
    .sum(sum_14[24]));
  AL_FADD comp14_25 (
    .a(i14[25]),
    .b(sum_13[25]),
    .c(cout_14[24]),
    .cout(cout_14[25]),
    .sum(sum_14[25]));
  AL_FADD comp14_26 (
    .a(i14[26]),
    .b(sum_13[26]),
    .c(cout_14[25]),
    .cout(cout_14[26]),
    .sum(sum_14[26]));
  AL_FADD comp14_27 (
    .a(i14[27]),
    .b(sum_13[27]),
    .c(cout_14[26]),
    .cout(cout_14[27]),
    .sum(sum_14[27]));
  AL_FADD comp14_28 (
    .a(i14[28]),
    .b(sum_13[28]),
    .c(cout_14[27]),
    .cout(cout_14[28]),
    .sum(sum_14[28]));
  AL_FADD comp14_29 (
    .a(i14[29]),
    .b(sum_13[29]),
    .c(cout_14[28]),
    .cout(cout_14[29]),
    .sum(sum_14[29]));
  AL_FADD comp14_3 (
    .a(i14[3]),
    .b(sum_13[3]),
    .c(cout_14[2]),
    .cout(cout_14[3]),
    .sum(sum_14[3]));
  AL_FADD comp14_30 (
    .a(i14[30]),
    .b(sum_13[30]),
    .c(cout_14[29]),
    .cout(cout_14[30]),
    .sum(sum_14[30]));
  AL_FADD comp14_31 (
    .a(i14[31]),
    .b(sum_13[31]),
    .c(cout_14[30]),
    .cout(cout_14[31]),
    .sum(sum_14[31]));
  AL_FADD comp14_32 (
    .a(i14[32]),
    .b(sum_13[32]),
    .c(cout_14[31]),
    .cout(cout_14[32]),
    .sum(sum_14[32]));
  AL_FADD comp14_33 (
    .a(i14[33]),
    .b(sum_13[33]),
    .c(cout_14[32]),
    .cout(cout_14[33]),
    .sum(sum_14[33]));
  AL_FADD comp14_34 (
    .a(i14[34]),
    .b(sum_13[34]),
    .c(cout_14[33]),
    .cout(cout_14[34]),
    .sum(sum_14[34]));
  AL_FADD comp14_35 (
    .a(i14[35]),
    .b(sum_13[35]),
    .c(cout_14[34]),
    .cout(cout_14[35]),
    .sum(sum_14[35]));
  AL_FADD comp14_36 (
    .a(i14[36]),
    .b(sum_13[36]),
    .c(cout_14[35]),
    .cout(cout_14[36]),
    .sum(sum_14[36]));
  AL_FADD comp14_37 (
    .a(i14[37]),
    .b(sum_13[37]),
    .c(cout_14[36]),
    .cout(cout_14[37]),
    .sum(sum_14[37]));
  AL_FADD comp14_38 (
    .a(i14[38]),
    .b(sum_13[38]),
    .c(cout_14[37]),
    .cout(cout_14[38]),
    .sum(sum_14[38]));
  AL_FADD comp14_39 (
    .a(i14[39]),
    .b(sum_13[39]),
    .c(cout_14[38]),
    .cout(cout_14[39]),
    .sum(sum_14[39]));
  AL_FADD comp14_4 (
    .a(i14[4]),
    .b(sum_13[4]),
    .c(cout_14[3]),
    .cout(cout_14[4]),
    .sum(sum_14[4]));
  AL_FADD comp14_40 (
    .a(i14[40]),
    .b(sum_13[40]),
    .c(cout_14[39]),
    .cout(cout_14[40]),
    .sum(sum_14[40]));
  AL_FADD comp14_41 (
    .a(i14[41]),
    .b(sum_13[41]),
    .c(cout_14[40]),
    .cout(cout_14[41]),
    .sum(sum_14[41]));
  AL_FADD comp14_42 (
    .a(i14[42]),
    .b(sum_13[42]),
    .c(cout_14[41]),
    .cout(cout_14[42]),
    .sum(sum_14[42]));
  AL_FADD comp14_43 (
    .a(i14[43]),
    .b(sum_13[43]),
    .c(cout_14[42]),
    .cout(cout_14[43]),
    .sum(sum_14[43]));
  AL_FADD comp14_44 (
    .a(i14[44]),
    .b(sum_13[44]),
    .c(cout_14[43]),
    .cout(cout_14[44]),
    .sum(sum_14[44]));
  AL_FADD comp14_45 (
    .a(i14[45]),
    .b(sum_13[45]),
    .c(cout_14[44]),
    .cout(cout_14[45]),
    .sum(sum_14[45]));
  AL_FADD comp14_46 (
    .a(i14[46]),
    .b(sum_13[46]),
    .c(cout_14[45]),
    .cout(cout_14[46]),
    .sum(sum_14[46]));
  AL_FADD comp14_47 (
    .a(i14[47]),
    .b(sum_13[47]),
    .c(cout_14[46]),
    .cout(cout_14[47]),
    .sum(sum_14[47]));
  AL_FADD comp14_48 (
    .a(1'b0),
    .b(sum_13[48]),
    .c(cout_14[47]),
    .cout(cout_14[48]),
    .sum(sum_14[48]));
  AL_FADD comp14_49 (
    .a(1'b0),
    .b(sum_13[49]),
    .c(cout_14[48]),
    .cout(cout_14[49]),
    .sum(sum_14[49]));
  AL_FADD comp14_5 (
    .a(i14[5]),
    .b(sum_13[5]),
    .c(cout_14[4]),
    .cout(cout_14[5]),
    .sum(sum_14[5]));
  AL_FADD comp14_50 (
    .a(1'b0),
    .b(sum_13[50]),
    .c(cout_14[49]),
    .cout(cout_14[50]),
    .sum(sum_14[50]));
  AL_FADD comp14_51 (
    .a(1'b0),
    .b(sum_13[51]),
    .c(cout_14[50]),
    .cout(cout_14[51]),
    .sum(sum_14[51]));
  AL_FADD comp14_52 (
    .a(1'b0),
    .b(sum_13[52]),
    .c(cout_14[51]),
    .cout(cout_14[52]),
    .sum(sum_14[52]));
  AL_FADD comp14_53 (
    .a(1'b0),
    .b(sum_13[53]),
    .c(cout_14[52]),
    .cout(cout_14[53]),
    .sum(sum_14[53]));
  AL_FADD comp14_54 (
    .a(1'b0),
    .b(sum_13[54]),
    .c(cout_14[53]),
    .cout(cout_14[54]),
    .sum(sum_14[54]));
  AL_FADD comp14_55 (
    .a(1'b0),
    .b(sum_13[55]),
    .c(cout_14[54]),
    .cout(cout_14[55]),
    .sum(sum_14[55]));
  AL_FADD comp14_56 (
    .a(1'b0),
    .b(sum_13[56]),
    .c(cout_14[55]),
    .cout(cout_14[56]),
    .sum(sum_14[56]));
  AL_FADD comp14_57 (
    .a(1'b0),
    .b(sum_13[57]),
    .c(cout_14[56]),
    .cout(cout_14[57]),
    .sum(sum_14[57]));
  AL_FADD comp14_58 (
    .a(1'b0),
    .b(sum_13[58]),
    .c(cout_14[57]),
    .cout(cout_14[58]),
    .sum(sum_14[58]));
  AL_FADD comp14_59 (
    .a(1'b0),
    .b(sum_13[59]),
    .c(cout_14[58]),
    .cout(cout_14[59]),
    .sum(sum_14[59]));
  AL_FADD comp14_6 (
    .a(i14[6]),
    .b(sum_13[6]),
    .c(cout_14[5]),
    .cout(cout_14[6]),
    .sum(sum_14[6]));
  AL_FADD comp14_60 (
    .a(1'b0),
    .b(sum_13[60]),
    .c(cout_14[59]),
    .cout(cout_14[60]),
    .sum(sum_14[60]));
  AL_FADD comp14_61 (
    .a(1'b0),
    .b(sum_13[61]),
    .c(cout_14[60]),
    .cout(cout_14[61]),
    .sum(sum_14[61]));
  AL_FADD comp14_62 (
    .a(1'b0),
    .b(sum_13[62]),
    .c(cout_14[61]),
    .cout(cout_14[62]),
    .sum(sum_14[62]));
  AL_FADD comp14_63 (
    .a(1'b0),
    .b(sum_13[63]),
    .c(cout_14[62]),
    .cout(cout_14[63]),
    .sum(sum_14[63]));
  AL_FADD comp14_7 (
    .a(i14[7]),
    .b(sum_13[7]),
    .c(cout_14[6]),
    .cout(cout_14[7]),
    .sum(sum_14[7]));
  AL_FADD comp14_8 (
    .a(i14[8]),
    .b(sum_13[8]),
    .c(cout_14[7]),
    .cout(cout_14[8]),
    .sum(sum_14[8]));
  AL_FADD comp14_9 (
    .a(i14[9]),
    .b(sum_13[9]),
    .c(cout_14[8]),
    .cout(cout_14[9]),
    .sum(sum_14[9]));
  AL_FADD comp15_0 (
    .a(i15[0]),
    .b(sum_14[0]),
    .c(1'b0),
    .cout(cout_15[0]),
    .sum(sum_15[0]));
  AL_FADD comp15_1 (
    .a(i15[1]),
    .b(sum_14[1]),
    .c(cout_15[0]),
    .cout(cout_15[1]),
    .sum(sum_15[1]));
  AL_FADD comp15_10 (
    .a(i15[10]),
    .b(sum_14[10]),
    .c(cout_15[9]),
    .cout(cout_15[10]),
    .sum(sum_15[10]));
  AL_FADD comp15_11 (
    .a(i15[11]),
    .b(sum_14[11]),
    .c(cout_15[10]),
    .cout(cout_15[11]),
    .sum(sum_15[11]));
  AL_FADD comp15_12 (
    .a(i15[12]),
    .b(sum_14[12]),
    .c(cout_15[11]),
    .cout(cout_15[12]),
    .sum(sum_15[12]));
  AL_FADD comp15_13 (
    .a(i15[13]),
    .b(sum_14[13]),
    .c(cout_15[12]),
    .cout(cout_15[13]),
    .sum(sum_15[13]));
  AL_FADD comp15_14 (
    .a(i15[14]),
    .b(sum_14[14]),
    .c(cout_15[13]),
    .cout(cout_15[14]),
    .sum(sum_15[14]));
  AL_FADD comp15_15 (
    .a(i15[15]),
    .b(sum_14[15]),
    .c(cout_15[14]),
    .cout(cout_15[15]),
    .sum(sum_15[15]));
  AL_FADD comp15_16 (
    .a(i15[16]),
    .b(sum_14[16]),
    .c(cout_15[15]),
    .cout(cout_15[16]),
    .sum(sum_15[16]));
  AL_FADD comp15_17 (
    .a(i15[17]),
    .b(sum_14[17]),
    .c(cout_15[16]),
    .cout(cout_15[17]),
    .sum(sum_15[17]));
  AL_FADD comp15_18 (
    .a(i15[18]),
    .b(sum_14[18]),
    .c(cout_15[17]),
    .cout(cout_15[18]),
    .sum(sum_15[18]));
  AL_FADD comp15_19 (
    .a(i15[19]),
    .b(sum_14[19]),
    .c(cout_15[18]),
    .cout(cout_15[19]),
    .sum(sum_15[19]));
  AL_FADD comp15_2 (
    .a(i15[2]),
    .b(sum_14[2]),
    .c(cout_15[1]),
    .cout(cout_15[2]),
    .sum(sum_15[2]));
  AL_FADD comp15_20 (
    .a(i15[20]),
    .b(sum_14[20]),
    .c(cout_15[19]),
    .cout(cout_15[20]),
    .sum(sum_15[20]));
  AL_FADD comp15_21 (
    .a(i15[21]),
    .b(sum_14[21]),
    .c(cout_15[20]),
    .cout(cout_15[21]),
    .sum(sum_15[21]));
  AL_FADD comp15_22 (
    .a(i15[22]),
    .b(sum_14[22]),
    .c(cout_15[21]),
    .cout(cout_15[22]),
    .sum(sum_15[22]));
  AL_FADD comp15_23 (
    .a(i15[23]),
    .b(sum_14[23]),
    .c(cout_15[22]),
    .cout(cout_15[23]),
    .sum(sum_15[23]));
  AL_FADD comp15_24 (
    .a(i15[24]),
    .b(sum_14[24]),
    .c(cout_15[23]),
    .cout(cout_15[24]),
    .sum(sum_15[24]));
  AL_FADD comp15_25 (
    .a(i15[25]),
    .b(sum_14[25]),
    .c(cout_15[24]),
    .cout(cout_15[25]),
    .sum(sum_15[25]));
  AL_FADD comp15_26 (
    .a(i15[26]),
    .b(sum_14[26]),
    .c(cout_15[25]),
    .cout(cout_15[26]),
    .sum(sum_15[26]));
  AL_FADD comp15_27 (
    .a(i15[27]),
    .b(sum_14[27]),
    .c(cout_15[26]),
    .cout(cout_15[27]),
    .sum(sum_15[27]));
  AL_FADD comp15_28 (
    .a(i15[28]),
    .b(sum_14[28]),
    .c(cout_15[27]),
    .cout(cout_15[28]),
    .sum(sum_15[28]));
  AL_FADD comp15_29 (
    .a(i15[29]),
    .b(sum_14[29]),
    .c(cout_15[28]),
    .cout(cout_15[29]),
    .sum(sum_15[29]));
  AL_FADD comp15_3 (
    .a(i15[3]),
    .b(sum_14[3]),
    .c(cout_15[2]),
    .cout(cout_15[3]),
    .sum(sum_15[3]));
  AL_FADD comp15_30 (
    .a(i15[30]),
    .b(sum_14[30]),
    .c(cout_15[29]),
    .cout(cout_15[30]),
    .sum(sum_15[30]));
  AL_FADD comp15_31 (
    .a(i15[31]),
    .b(sum_14[31]),
    .c(cout_15[30]),
    .cout(cout_15[31]),
    .sum(sum_15[31]));
  AL_FADD comp15_32 (
    .a(i15[32]),
    .b(sum_14[32]),
    .c(cout_15[31]),
    .cout(cout_15[32]),
    .sum(sum_15[32]));
  AL_FADD comp15_33 (
    .a(i15[33]),
    .b(sum_14[33]),
    .c(cout_15[32]),
    .cout(cout_15[33]),
    .sum(sum_15[33]));
  AL_FADD comp15_34 (
    .a(i15[34]),
    .b(sum_14[34]),
    .c(cout_15[33]),
    .cout(cout_15[34]),
    .sum(sum_15[34]));
  AL_FADD comp15_35 (
    .a(i15[35]),
    .b(sum_14[35]),
    .c(cout_15[34]),
    .cout(cout_15[35]),
    .sum(sum_15[35]));
  AL_FADD comp15_36 (
    .a(i15[36]),
    .b(sum_14[36]),
    .c(cout_15[35]),
    .cout(cout_15[36]),
    .sum(sum_15[36]));
  AL_FADD comp15_37 (
    .a(i15[37]),
    .b(sum_14[37]),
    .c(cout_15[36]),
    .cout(cout_15[37]),
    .sum(sum_15[37]));
  AL_FADD comp15_38 (
    .a(i15[38]),
    .b(sum_14[38]),
    .c(cout_15[37]),
    .cout(cout_15[38]),
    .sum(sum_15[38]));
  AL_FADD comp15_39 (
    .a(i15[39]),
    .b(sum_14[39]),
    .c(cout_15[38]),
    .cout(cout_15[39]),
    .sum(sum_15[39]));
  AL_FADD comp15_4 (
    .a(i15[4]),
    .b(sum_14[4]),
    .c(cout_15[3]),
    .cout(cout_15[4]),
    .sum(sum_15[4]));
  AL_FADD comp15_40 (
    .a(i15[40]),
    .b(sum_14[40]),
    .c(cout_15[39]),
    .cout(cout_15[40]),
    .sum(sum_15[40]));
  AL_FADD comp15_41 (
    .a(i15[41]),
    .b(sum_14[41]),
    .c(cout_15[40]),
    .cout(cout_15[41]),
    .sum(sum_15[41]));
  AL_FADD comp15_42 (
    .a(i15[42]),
    .b(sum_14[42]),
    .c(cout_15[41]),
    .cout(cout_15[42]),
    .sum(sum_15[42]));
  AL_FADD comp15_43 (
    .a(i15[43]),
    .b(sum_14[43]),
    .c(cout_15[42]),
    .cout(cout_15[43]),
    .sum(sum_15[43]));
  AL_FADD comp15_44 (
    .a(i15[44]),
    .b(sum_14[44]),
    .c(cout_15[43]),
    .cout(cout_15[44]),
    .sum(sum_15[44]));
  AL_FADD comp15_45 (
    .a(i15[45]),
    .b(sum_14[45]),
    .c(cout_15[44]),
    .cout(cout_15[45]),
    .sum(sum_15[45]));
  AL_FADD comp15_46 (
    .a(i15[46]),
    .b(sum_14[46]),
    .c(cout_15[45]),
    .cout(cout_15[46]),
    .sum(sum_15[46]));
  AL_FADD comp15_47 (
    .a(1'b0),
    .b(sum_14[47]),
    .c(cout_15[46]),
    .cout(cout_15[47]),
    .sum(sum_15[47]));
  AL_FADD comp15_48 (
    .a(1'b0),
    .b(sum_14[48]),
    .c(cout_15[47]),
    .cout(cout_15[48]),
    .sum(sum_15[48]));
  AL_FADD comp15_49 (
    .a(1'b0),
    .b(sum_14[49]),
    .c(cout_15[48]),
    .cout(cout_15[49]),
    .sum(sum_15[49]));
  AL_FADD comp15_5 (
    .a(i15[5]),
    .b(sum_14[5]),
    .c(cout_15[4]),
    .cout(cout_15[5]),
    .sum(sum_15[5]));
  AL_FADD comp15_50 (
    .a(1'b0),
    .b(sum_14[50]),
    .c(cout_15[49]),
    .cout(cout_15[50]),
    .sum(sum_15[50]));
  AL_FADD comp15_51 (
    .a(1'b0),
    .b(sum_14[51]),
    .c(cout_15[50]),
    .cout(cout_15[51]),
    .sum(sum_15[51]));
  AL_FADD comp15_52 (
    .a(1'b0),
    .b(sum_14[52]),
    .c(cout_15[51]),
    .cout(cout_15[52]),
    .sum(sum_15[52]));
  AL_FADD comp15_53 (
    .a(1'b0),
    .b(sum_14[53]),
    .c(cout_15[52]),
    .cout(cout_15[53]),
    .sum(sum_15[53]));
  AL_FADD comp15_54 (
    .a(1'b0),
    .b(sum_14[54]),
    .c(cout_15[53]),
    .cout(cout_15[54]),
    .sum(sum_15[54]));
  AL_FADD comp15_55 (
    .a(1'b0),
    .b(sum_14[55]),
    .c(cout_15[54]),
    .cout(cout_15[55]),
    .sum(sum_15[55]));
  AL_FADD comp15_56 (
    .a(1'b0),
    .b(sum_14[56]),
    .c(cout_15[55]),
    .cout(cout_15[56]),
    .sum(sum_15[56]));
  AL_FADD comp15_57 (
    .a(1'b0),
    .b(sum_14[57]),
    .c(cout_15[56]),
    .cout(cout_15[57]),
    .sum(sum_15[57]));
  AL_FADD comp15_58 (
    .a(1'b0),
    .b(sum_14[58]),
    .c(cout_15[57]),
    .cout(cout_15[58]),
    .sum(sum_15[58]));
  AL_FADD comp15_59 (
    .a(1'b0),
    .b(sum_14[59]),
    .c(cout_15[58]),
    .cout(cout_15[59]),
    .sum(sum_15[59]));
  AL_FADD comp15_6 (
    .a(i15[6]),
    .b(sum_14[6]),
    .c(cout_15[5]),
    .cout(cout_15[6]),
    .sum(sum_15[6]));
  AL_FADD comp15_60 (
    .a(1'b0),
    .b(sum_14[60]),
    .c(cout_15[59]),
    .cout(cout_15[60]),
    .sum(sum_15[60]));
  AL_FADD comp15_61 (
    .a(1'b0),
    .b(sum_14[61]),
    .c(cout_15[60]),
    .cout(cout_15[61]),
    .sum(sum_15[61]));
  AL_FADD comp15_62 (
    .a(1'b0),
    .b(sum_14[62]),
    .c(cout_15[61]),
    .cout(cout_15[62]),
    .sum(sum_15[62]));
  AL_FADD comp15_63 (
    .a(1'b0),
    .b(sum_14[63]),
    .c(cout_15[62]),
    .cout(cout_15[63]),
    .sum(sum_15[63]));
  AL_FADD comp15_7 (
    .a(i15[7]),
    .b(sum_14[7]),
    .c(cout_15[6]),
    .cout(cout_15[7]),
    .sum(sum_15[7]));
  AL_FADD comp15_8 (
    .a(i15[8]),
    .b(sum_14[8]),
    .c(cout_15[7]),
    .cout(cout_15[8]),
    .sum(sum_15[8]));
  AL_FADD comp15_9 (
    .a(i15[9]),
    .b(sum_14[9]),
    .c(cout_15[8]),
    .cout(cout_15[9]),
    .sum(sum_15[9]));
  AL_FADD comp16_0 (
    .a(i16[0]),
    .b(sum_15[0]),
    .c(1'b0),
    .cout(cout_16[0]),
    .sum(sum_16[0]));
  AL_FADD comp16_1 (
    .a(i16[1]),
    .b(sum_15[1]),
    .c(cout_16[0]),
    .cout(cout_16[1]),
    .sum(sum_16[1]));
  AL_FADD comp16_10 (
    .a(i16[10]),
    .b(sum_15[10]),
    .c(cout_16[9]),
    .cout(cout_16[10]),
    .sum(sum_16[10]));
  AL_FADD comp16_11 (
    .a(i16[11]),
    .b(sum_15[11]),
    .c(cout_16[10]),
    .cout(cout_16[11]),
    .sum(sum_16[11]));
  AL_FADD comp16_12 (
    .a(i16[12]),
    .b(sum_15[12]),
    .c(cout_16[11]),
    .cout(cout_16[12]),
    .sum(sum_16[12]));
  AL_FADD comp16_13 (
    .a(i16[13]),
    .b(sum_15[13]),
    .c(cout_16[12]),
    .cout(cout_16[13]),
    .sum(sum_16[13]));
  AL_FADD comp16_14 (
    .a(i16[14]),
    .b(sum_15[14]),
    .c(cout_16[13]),
    .cout(cout_16[14]),
    .sum(sum_16[14]));
  AL_FADD comp16_15 (
    .a(i16[15]),
    .b(sum_15[15]),
    .c(cout_16[14]),
    .cout(cout_16[15]),
    .sum(sum_16[15]));
  AL_FADD comp16_16 (
    .a(i16[16]),
    .b(sum_15[16]),
    .c(cout_16[15]),
    .cout(cout_16[16]),
    .sum(sum_16[16]));
  AL_FADD comp16_17 (
    .a(i16[17]),
    .b(sum_15[17]),
    .c(cout_16[16]),
    .cout(cout_16[17]),
    .sum(sum_16[17]));
  AL_FADD comp16_18 (
    .a(i16[18]),
    .b(sum_15[18]),
    .c(cout_16[17]),
    .cout(cout_16[18]),
    .sum(sum_16[18]));
  AL_FADD comp16_19 (
    .a(i16[19]),
    .b(sum_15[19]),
    .c(cout_16[18]),
    .cout(cout_16[19]),
    .sum(sum_16[19]));
  AL_FADD comp16_2 (
    .a(i16[2]),
    .b(sum_15[2]),
    .c(cout_16[1]),
    .cout(cout_16[2]),
    .sum(sum_16[2]));
  AL_FADD comp16_20 (
    .a(i16[20]),
    .b(sum_15[20]),
    .c(cout_16[19]),
    .cout(cout_16[20]),
    .sum(sum_16[20]));
  AL_FADD comp16_21 (
    .a(i16[21]),
    .b(sum_15[21]),
    .c(cout_16[20]),
    .cout(cout_16[21]),
    .sum(sum_16[21]));
  AL_FADD comp16_22 (
    .a(i16[22]),
    .b(sum_15[22]),
    .c(cout_16[21]),
    .cout(cout_16[22]),
    .sum(sum_16[22]));
  AL_FADD comp16_23 (
    .a(i16[23]),
    .b(sum_15[23]),
    .c(cout_16[22]),
    .cout(cout_16[23]),
    .sum(sum_16[23]));
  AL_FADD comp16_24 (
    .a(i16[24]),
    .b(sum_15[24]),
    .c(cout_16[23]),
    .cout(cout_16[24]),
    .sum(sum_16[24]));
  AL_FADD comp16_25 (
    .a(i16[25]),
    .b(sum_15[25]),
    .c(cout_16[24]),
    .cout(cout_16[25]),
    .sum(sum_16[25]));
  AL_FADD comp16_26 (
    .a(i16[26]),
    .b(sum_15[26]),
    .c(cout_16[25]),
    .cout(cout_16[26]),
    .sum(sum_16[26]));
  AL_FADD comp16_27 (
    .a(i16[27]),
    .b(sum_15[27]),
    .c(cout_16[26]),
    .cout(cout_16[27]),
    .sum(sum_16[27]));
  AL_FADD comp16_28 (
    .a(i16[28]),
    .b(sum_15[28]),
    .c(cout_16[27]),
    .cout(cout_16[28]),
    .sum(sum_16[28]));
  AL_FADD comp16_29 (
    .a(i16[29]),
    .b(sum_15[29]),
    .c(cout_16[28]),
    .cout(cout_16[29]),
    .sum(sum_16[29]));
  AL_FADD comp16_3 (
    .a(i16[3]),
    .b(sum_15[3]),
    .c(cout_16[2]),
    .cout(cout_16[3]),
    .sum(sum_16[3]));
  AL_FADD comp16_30 (
    .a(i16[30]),
    .b(sum_15[30]),
    .c(cout_16[29]),
    .cout(cout_16[30]),
    .sum(sum_16[30]));
  AL_FADD comp16_31 (
    .a(i16[31]),
    .b(sum_15[31]),
    .c(cout_16[30]),
    .cout(cout_16[31]),
    .sum(sum_16[31]));
  AL_FADD comp16_32 (
    .a(i16[32]),
    .b(sum_15[32]),
    .c(cout_16[31]),
    .cout(cout_16[32]),
    .sum(sum_16[32]));
  AL_FADD comp16_33 (
    .a(i16[33]),
    .b(sum_15[33]),
    .c(cout_16[32]),
    .cout(cout_16[33]),
    .sum(sum_16[33]));
  AL_FADD comp16_34 (
    .a(i16[34]),
    .b(sum_15[34]),
    .c(cout_16[33]),
    .cout(cout_16[34]),
    .sum(sum_16[34]));
  AL_FADD comp16_35 (
    .a(i16[35]),
    .b(sum_15[35]),
    .c(cout_16[34]),
    .cout(cout_16[35]),
    .sum(sum_16[35]));
  AL_FADD comp16_36 (
    .a(i16[36]),
    .b(sum_15[36]),
    .c(cout_16[35]),
    .cout(cout_16[36]),
    .sum(sum_16[36]));
  AL_FADD comp16_37 (
    .a(i16[37]),
    .b(sum_15[37]),
    .c(cout_16[36]),
    .cout(cout_16[37]),
    .sum(sum_16[37]));
  AL_FADD comp16_38 (
    .a(i16[38]),
    .b(sum_15[38]),
    .c(cout_16[37]),
    .cout(cout_16[38]),
    .sum(sum_16[38]));
  AL_FADD comp16_39 (
    .a(i16[39]),
    .b(sum_15[39]),
    .c(cout_16[38]),
    .cout(cout_16[39]),
    .sum(sum_16[39]));
  AL_FADD comp16_4 (
    .a(i16[4]),
    .b(sum_15[4]),
    .c(cout_16[3]),
    .cout(cout_16[4]),
    .sum(sum_16[4]));
  AL_FADD comp16_40 (
    .a(i16[40]),
    .b(sum_15[40]),
    .c(cout_16[39]),
    .cout(cout_16[40]),
    .sum(sum_16[40]));
  AL_FADD comp16_41 (
    .a(i16[41]),
    .b(sum_15[41]),
    .c(cout_16[40]),
    .cout(cout_16[41]),
    .sum(sum_16[41]));
  AL_FADD comp16_42 (
    .a(i16[42]),
    .b(sum_15[42]),
    .c(cout_16[41]),
    .cout(cout_16[42]),
    .sum(sum_16[42]));
  AL_FADD comp16_43 (
    .a(i16[43]),
    .b(sum_15[43]),
    .c(cout_16[42]),
    .cout(cout_16[43]),
    .sum(sum_16[43]));
  AL_FADD comp16_44 (
    .a(i16[44]),
    .b(sum_15[44]),
    .c(cout_16[43]),
    .cout(cout_16[44]),
    .sum(sum_16[44]));
  AL_FADD comp16_45 (
    .a(i16[45]),
    .b(sum_15[45]),
    .c(cout_16[44]),
    .cout(cout_16[45]),
    .sum(sum_16[45]));
  AL_FADD comp16_46 (
    .a(1'b0),
    .b(sum_15[46]),
    .c(cout_16[45]),
    .cout(cout_16[46]),
    .sum(sum_16[46]));
  AL_FADD comp16_47 (
    .a(1'b0),
    .b(sum_15[47]),
    .c(cout_16[46]),
    .cout(cout_16[47]),
    .sum(sum_16[47]));
  AL_FADD comp16_48 (
    .a(1'b0),
    .b(sum_15[48]),
    .c(cout_16[47]),
    .cout(cout_16[48]),
    .sum(sum_16[48]));
  AL_FADD comp16_49 (
    .a(1'b0),
    .b(sum_15[49]),
    .c(cout_16[48]),
    .cout(cout_16[49]),
    .sum(sum_16[49]));
  AL_FADD comp16_5 (
    .a(i16[5]),
    .b(sum_15[5]),
    .c(cout_16[4]),
    .cout(cout_16[5]),
    .sum(sum_16[5]));
  AL_FADD comp16_50 (
    .a(1'b0),
    .b(sum_15[50]),
    .c(cout_16[49]),
    .cout(cout_16[50]),
    .sum(sum_16[50]));
  AL_FADD comp16_51 (
    .a(1'b0),
    .b(sum_15[51]),
    .c(cout_16[50]),
    .cout(cout_16[51]),
    .sum(sum_16[51]));
  AL_FADD comp16_52 (
    .a(1'b0),
    .b(sum_15[52]),
    .c(cout_16[51]),
    .cout(cout_16[52]),
    .sum(sum_16[52]));
  AL_FADD comp16_53 (
    .a(1'b0),
    .b(sum_15[53]),
    .c(cout_16[52]),
    .cout(cout_16[53]),
    .sum(sum_16[53]));
  AL_FADD comp16_54 (
    .a(1'b0),
    .b(sum_15[54]),
    .c(cout_16[53]),
    .cout(cout_16[54]),
    .sum(sum_16[54]));
  AL_FADD comp16_55 (
    .a(1'b0),
    .b(sum_15[55]),
    .c(cout_16[54]),
    .cout(cout_16[55]),
    .sum(sum_16[55]));
  AL_FADD comp16_56 (
    .a(1'b0),
    .b(sum_15[56]),
    .c(cout_16[55]),
    .cout(cout_16[56]),
    .sum(sum_16[56]));
  AL_FADD comp16_57 (
    .a(1'b0),
    .b(sum_15[57]),
    .c(cout_16[56]),
    .cout(cout_16[57]),
    .sum(sum_16[57]));
  AL_FADD comp16_58 (
    .a(1'b0),
    .b(sum_15[58]),
    .c(cout_16[57]),
    .cout(cout_16[58]),
    .sum(sum_16[58]));
  AL_FADD comp16_59 (
    .a(1'b0),
    .b(sum_15[59]),
    .c(cout_16[58]),
    .cout(cout_16[59]),
    .sum(sum_16[59]));
  AL_FADD comp16_6 (
    .a(i16[6]),
    .b(sum_15[6]),
    .c(cout_16[5]),
    .cout(cout_16[6]),
    .sum(sum_16[6]));
  AL_FADD comp16_60 (
    .a(1'b0),
    .b(sum_15[60]),
    .c(cout_16[59]),
    .cout(cout_16[60]),
    .sum(sum_16[60]));
  AL_FADD comp16_61 (
    .a(1'b0),
    .b(sum_15[61]),
    .c(cout_16[60]),
    .cout(cout_16[61]),
    .sum(sum_16[61]));
  AL_FADD comp16_62 (
    .a(1'b0),
    .b(sum_15[62]),
    .c(cout_16[61]),
    .cout(cout_16[62]),
    .sum(sum_16[62]));
  AL_FADD comp16_63 (
    .a(1'b0),
    .b(sum_15[63]),
    .c(cout_16[62]),
    .cout(cout_16[63]),
    .sum(sum_16[63]));
  AL_FADD comp16_7 (
    .a(i16[7]),
    .b(sum_15[7]),
    .c(cout_16[6]),
    .cout(cout_16[7]),
    .sum(sum_16[7]));
  AL_FADD comp16_8 (
    .a(i16[8]),
    .b(sum_15[8]),
    .c(cout_16[7]),
    .cout(cout_16[8]),
    .sum(sum_16[8]));
  AL_FADD comp16_9 (
    .a(i16[9]),
    .b(sum_15[9]),
    .c(cout_16[8]),
    .cout(cout_16[9]),
    .sum(sum_16[9]));
  AL_FADD comp17_0 (
    .a(i17[0]),
    .b(sum_16[0]),
    .c(1'b0),
    .cout(cout_17[0]),
    .sum(sum_17[0]));
  AL_FADD comp17_1 (
    .a(i17[1]),
    .b(sum_16[1]),
    .c(cout_17[0]),
    .cout(cout_17[1]),
    .sum(sum_17[1]));
  AL_FADD comp17_10 (
    .a(i17[10]),
    .b(sum_16[10]),
    .c(cout_17[9]),
    .cout(cout_17[10]),
    .sum(sum_17[10]));
  AL_FADD comp17_11 (
    .a(i17[11]),
    .b(sum_16[11]),
    .c(cout_17[10]),
    .cout(cout_17[11]),
    .sum(sum_17[11]));
  AL_FADD comp17_12 (
    .a(i17[12]),
    .b(sum_16[12]),
    .c(cout_17[11]),
    .cout(cout_17[12]),
    .sum(sum_17[12]));
  AL_FADD comp17_13 (
    .a(i17[13]),
    .b(sum_16[13]),
    .c(cout_17[12]),
    .cout(cout_17[13]),
    .sum(sum_17[13]));
  AL_FADD comp17_14 (
    .a(i17[14]),
    .b(sum_16[14]),
    .c(cout_17[13]),
    .cout(cout_17[14]),
    .sum(sum_17[14]));
  AL_FADD comp17_15 (
    .a(i17[15]),
    .b(sum_16[15]),
    .c(cout_17[14]),
    .cout(cout_17[15]),
    .sum(sum_17[15]));
  AL_FADD comp17_16 (
    .a(i17[16]),
    .b(sum_16[16]),
    .c(cout_17[15]),
    .cout(cout_17[16]),
    .sum(sum_17[16]));
  AL_FADD comp17_17 (
    .a(i17[17]),
    .b(sum_16[17]),
    .c(cout_17[16]),
    .cout(cout_17[17]),
    .sum(sum_17[17]));
  AL_FADD comp17_18 (
    .a(i17[18]),
    .b(sum_16[18]),
    .c(cout_17[17]),
    .cout(cout_17[18]),
    .sum(sum_17[18]));
  AL_FADD comp17_19 (
    .a(i17[19]),
    .b(sum_16[19]),
    .c(cout_17[18]),
    .cout(cout_17[19]),
    .sum(sum_17[19]));
  AL_FADD comp17_2 (
    .a(i17[2]),
    .b(sum_16[2]),
    .c(cout_17[1]),
    .cout(cout_17[2]),
    .sum(sum_17[2]));
  AL_FADD comp17_20 (
    .a(i17[20]),
    .b(sum_16[20]),
    .c(cout_17[19]),
    .cout(cout_17[20]),
    .sum(sum_17[20]));
  AL_FADD comp17_21 (
    .a(i17[21]),
    .b(sum_16[21]),
    .c(cout_17[20]),
    .cout(cout_17[21]),
    .sum(sum_17[21]));
  AL_FADD comp17_22 (
    .a(i17[22]),
    .b(sum_16[22]),
    .c(cout_17[21]),
    .cout(cout_17[22]),
    .sum(sum_17[22]));
  AL_FADD comp17_23 (
    .a(i17[23]),
    .b(sum_16[23]),
    .c(cout_17[22]),
    .cout(cout_17[23]),
    .sum(sum_17[23]));
  AL_FADD comp17_24 (
    .a(i17[24]),
    .b(sum_16[24]),
    .c(cout_17[23]),
    .cout(cout_17[24]),
    .sum(sum_17[24]));
  AL_FADD comp17_25 (
    .a(i17[25]),
    .b(sum_16[25]),
    .c(cout_17[24]),
    .cout(cout_17[25]),
    .sum(sum_17[25]));
  AL_FADD comp17_26 (
    .a(i17[26]),
    .b(sum_16[26]),
    .c(cout_17[25]),
    .cout(cout_17[26]),
    .sum(sum_17[26]));
  AL_FADD comp17_27 (
    .a(i17[27]),
    .b(sum_16[27]),
    .c(cout_17[26]),
    .cout(cout_17[27]),
    .sum(sum_17[27]));
  AL_FADD comp17_28 (
    .a(i17[28]),
    .b(sum_16[28]),
    .c(cout_17[27]),
    .cout(cout_17[28]),
    .sum(sum_17[28]));
  AL_FADD comp17_29 (
    .a(i17[29]),
    .b(sum_16[29]),
    .c(cout_17[28]),
    .cout(cout_17[29]),
    .sum(sum_17[29]));
  AL_FADD comp17_3 (
    .a(i17[3]),
    .b(sum_16[3]),
    .c(cout_17[2]),
    .cout(cout_17[3]),
    .sum(sum_17[3]));
  AL_FADD comp17_30 (
    .a(i17[30]),
    .b(sum_16[30]),
    .c(cout_17[29]),
    .cout(cout_17[30]),
    .sum(sum_17[30]));
  AL_FADD comp17_31 (
    .a(i17[31]),
    .b(sum_16[31]),
    .c(cout_17[30]),
    .cout(cout_17[31]),
    .sum(sum_17[31]));
  AL_FADD comp17_32 (
    .a(i17[32]),
    .b(sum_16[32]),
    .c(cout_17[31]),
    .cout(cout_17[32]),
    .sum(sum_17[32]));
  AL_FADD comp17_33 (
    .a(i17[33]),
    .b(sum_16[33]),
    .c(cout_17[32]),
    .cout(cout_17[33]),
    .sum(sum_17[33]));
  AL_FADD comp17_34 (
    .a(i17[34]),
    .b(sum_16[34]),
    .c(cout_17[33]),
    .cout(cout_17[34]),
    .sum(sum_17[34]));
  AL_FADD comp17_35 (
    .a(i17[35]),
    .b(sum_16[35]),
    .c(cout_17[34]),
    .cout(cout_17[35]),
    .sum(sum_17[35]));
  AL_FADD comp17_36 (
    .a(i17[36]),
    .b(sum_16[36]),
    .c(cout_17[35]),
    .cout(cout_17[36]),
    .sum(sum_17[36]));
  AL_FADD comp17_37 (
    .a(i17[37]),
    .b(sum_16[37]),
    .c(cout_17[36]),
    .cout(cout_17[37]),
    .sum(sum_17[37]));
  AL_FADD comp17_38 (
    .a(i17[38]),
    .b(sum_16[38]),
    .c(cout_17[37]),
    .cout(cout_17[38]),
    .sum(sum_17[38]));
  AL_FADD comp17_39 (
    .a(i17[39]),
    .b(sum_16[39]),
    .c(cout_17[38]),
    .cout(cout_17[39]),
    .sum(sum_17[39]));
  AL_FADD comp17_4 (
    .a(i17[4]),
    .b(sum_16[4]),
    .c(cout_17[3]),
    .cout(cout_17[4]),
    .sum(sum_17[4]));
  AL_FADD comp17_40 (
    .a(i17[40]),
    .b(sum_16[40]),
    .c(cout_17[39]),
    .cout(cout_17[40]),
    .sum(sum_17[40]));
  AL_FADD comp17_41 (
    .a(i17[41]),
    .b(sum_16[41]),
    .c(cout_17[40]),
    .cout(cout_17[41]),
    .sum(sum_17[41]));
  AL_FADD comp17_42 (
    .a(i17[42]),
    .b(sum_16[42]),
    .c(cout_17[41]),
    .cout(cout_17[42]),
    .sum(sum_17[42]));
  AL_FADD comp17_43 (
    .a(i17[43]),
    .b(sum_16[43]),
    .c(cout_17[42]),
    .cout(cout_17[43]),
    .sum(sum_17[43]));
  AL_FADD comp17_44 (
    .a(i17[44]),
    .b(sum_16[44]),
    .c(cout_17[43]),
    .cout(cout_17[44]),
    .sum(sum_17[44]));
  AL_FADD comp17_45 (
    .a(1'b0),
    .b(sum_16[45]),
    .c(cout_17[44]),
    .cout(cout_17[45]),
    .sum(sum_17[45]));
  AL_FADD comp17_46 (
    .a(1'b0),
    .b(sum_16[46]),
    .c(cout_17[45]),
    .cout(cout_17[46]),
    .sum(sum_17[46]));
  AL_FADD comp17_47 (
    .a(1'b0),
    .b(sum_16[47]),
    .c(cout_17[46]),
    .cout(cout_17[47]),
    .sum(sum_17[47]));
  AL_FADD comp17_48 (
    .a(1'b0),
    .b(sum_16[48]),
    .c(cout_17[47]),
    .cout(cout_17[48]),
    .sum(sum_17[48]));
  AL_FADD comp17_49 (
    .a(1'b0),
    .b(sum_16[49]),
    .c(cout_17[48]),
    .cout(cout_17[49]),
    .sum(sum_17[49]));
  AL_FADD comp17_5 (
    .a(i17[5]),
    .b(sum_16[5]),
    .c(cout_17[4]),
    .cout(cout_17[5]),
    .sum(sum_17[5]));
  AL_FADD comp17_50 (
    .a(1'b0),
    .b(sum_16[50]),
    .c(cout_17[49]),
    .cout(cout_17[50]),
    .sum(sum_17[50]));
  AL_FADD comp17_51 (
    .a(1'b0),
    .b(sum_16[51]),
    .c(cout_17[50]),
    .cout(cout_17[51]),
    .sum(sum_17[51]));
  AL_FADD comp17_52 (
    .a(1'b0),
    .b(sum_16[52]),
    .c(cout_17[51]),
    .cout(cout_17[52]),
    .sum(sum_17[52]));
  AL_FADD comp17_53 (
    .a(1'b0),
    .b(sum_16[53]),
    .c(cout_17[52]),
    .cout(cout_17[53]),
    .sum(sum_17[53]));
  AL_FADD comp17_54 (
    .a(1'b0),
    .b(sum_16[54]),
    .c(cout_17[53]),
    .cout(cout_17[54]),
    .sum(sum_17[54]));
  AL_FADD comp17_55 (
    .a(1'b0),
    .b(sum_16[55]),
    .c(cout_17[54]),
    .cout(cout_17[55]),
    .sum(sum_17[55]));
  AL_FADD comp17_56 (
    .a(1'b0),
    .b(sum_16[56]),
    .c(cout_17[55]),
    .cout(cout_17[56]),
    .sum(sum_17[56]));
  AL_FADD comp17_57 (
    .a(1'b0),
    .b(sum_16[57]),
    .c(cout_17[56]),
    .cout(cout_17[57]),
    .sum(sum_17[57]));
  AL_FADD comp17_58 (
    .a(1'b0),
    .b(sum_16[58]),
    .c(cout_17[57]),
    .cout(cout_17[58]),
    .sum(sum_17[58]));
  AL_FADD comp17_59 (
    .a(1'b0),
    .b(sum_16[59]),
    .c(cout_17[58]),
    .cout(cout_17[59]),
    .sum(sum_17[59]));
  AL_FADD comp17_6 (
    .a(i17[6]),
    .b(sum_16[6]),
    .c(cout_17[5]),
    .cout(cout_17[6]),
    .sum(sum_17[6]));
  AL_FADD comp17_60 (
    .a(1'b0),
    .b(sum_16[60]),
    .c(cout_17[59]),
    .cout(cout_17[60]),
    .sum(sum_17[60]));
  AL_FADD comp17_61 (
    .a(1'b0),
    .b(sum_16[61]),
    .c(cout_17[60]),
    .cout(cout_17[61]),
    .sum(sum_17[61]));
  AL_FADD comp17_62 (
    .a(1'b0),
    .b(sum_16[62]),
    .c(cout_17[61]),
    .cout(cout_17[62]),
    .sum(sum_17[62]));
  AL_FADD comp17_63 (
    .a(1'b0),
    .b(sum_16[63]),
    .c(cout_17[62]),
    .cout(cout_17[63]),
    .sum(sum_17[63]));
  AL_FADD comp17_7 (
    .a(i17[7]),
    .b(sum_16[7]),
    .c(cout_17[6]),
    .cout(cout_17[7]),
    .sum(sum_17[7]));
  AL_FADD comp17_8 (
    .a(i17[8]),
    .b(sum_16[8]),
    .c(cout_17[7]),
    .cout(cout_17[8]),
    .sum(sum_17[8]));
  AL_FADD comp17_9 (
    .a(i17[9]),
    .b(sum_16[9]),
    .c(cout_17[8]),
    .cout(cout_17[9]),
    .sum(sum_17[9]));
  AL_FADD comp18_0 (
    .a(i18[0]),
    .b(sum_17[0]),
    .c(1'b0),
    .cout(cout_18[0]),
    .sum(sum_18[0]));
  AL_FADD comp18_1 (
    .a(i18[1]),
    .b(sum_17[1]),
    .c(cout_18[0]),
    .cout(cout_18[1]),
    .sum(sum_18[1]));
  AL_FADD comp18_10 (
    .a(i18[10]),
    .b(sum_17[10]),
    .c(cout_18[9]),
    .cout(cout_18[10]),
    .sum(sum_18[10]));
  AL_FADD comp18_11 (
    .a(i18[11]),
    .b(sum_17[11]),
    .c(cout_18[10]),
    .cout(cout_18[11]),
    .sum(sum_18[11]));
  AL_FADD comp18_12 (
    .a(i18[12]),
    .b(sum_17[12]),
    .c(cout_18[11]),
    .cout(cout_18[12]),
    .sum(sum_18[12]));
  AL_FADD comp18_13 (
    .a(i18[13]),
    .b(sum_17[13]),
    .c(cout_18[12]),
    .cout(cout_18[13]),
    .sum(sum_18[13]));
  AL_FADD comp18_14 (
    .a(i18[14]),
    .b(sum_17[14]),
    .c(cout_18[13]),
    .cout(cout_18[14]),
    .sum(sum_18[14]));
  AL_FADD comp18_15 (
    .a(i18[15]),
    .b(sum_17[15]),
    .c(cout_18[14]),
    .cout(cout_18[15]),
    .sum(sum_18[15]));
  AL_FADD comp18_16 (
    .a(i18[16]),
    .b(sum_17[16]),
    .c(cout_18[15]),
    .cout(cout_18[16]),
    .sum(sum_18[16]));
  AL_FADD comp18_17 (
    .a(i18[17]),
    .b(sum_17[17]),
    .c(cout_18[16]),
    .cout(cout_18[17]),
    .sum(sum_18[17]));
  AL_FADD comp18_18 (
    .a(i18[18]),
    .b(sum_17[18]),
    .c(cout_18[17]),
    .cout(cout_18[18]),
    .sum(sum_18[18]));
  AL_FADD comp18_19 (
    .a(i18[19]),
    .b(sum_17[19]),
    .c(cout_18[18]),
    .cout(cout_18[19]),
    .sum(sum_18[19]));
  AL_FADD comp18_2 (
    .a(i18[2]),
    .b(sum_17[2]),
    .c(cout_18[1]),
    .cout(cout_18[2]),
    .sum(sum_18[2]));
  AL_FADD comp18_20 (
    .a(i18[20]),
    .b(sum_17[20]),
    .c(cout_18[19]),
    .cout(cout_18[20]),
    .sum(sum_18[20]));
  AL_FADD comp18_21 (
    .a(i18[21]),
    .b(sum_17[21]),
    .c(cout_18[20]),
    .cout(cout_18[21]),
    .sum(sum_18[21]));
  AL_FADD comp18_22 (
    .a(i18[22]),
    .b(sum_17[22]),
    .c(cout_18[21]),
    .cout(cout_18[22]),
    .sum(sum_18[22]));
  AL_FADD comp18_23 (
    .a(i18[23]),
    .b(sum_17[23]),
    .c(cout_18[22]),
    .cout(cout_18[23]),
    .sum(sum_18[23]));
  AL_FADD comp18_24 (
    .a(i18[24]),
    .b(sum_17[24]),
    .c(cout_18[23]),
    .cout(cout_18[24]),
    .sum(sum_18[24]));
  AL_FADD comp18_25 (
    .a(i18[25]),
    .b(sum_17[25]),
    .c(cout_18[24]),
    .cout(cout_18[25]),
    .sum(sum_18[25]));
  AL_FADD comp18_26 (
    .a(i18[26]),
    .b(sum_17[26]),
    .c(cout_18[25]),
    .cout(cout_18[26]),
    .sum(sum_18[26]));
  AL_FADD comp18_27 (
    .a(i18[27]),
    .b(sum_17[27]),
    .c(cout_18[26]),
    .cout(cout_18[27]),
    .sum(sum_18[27]));
  AL_FADD comp18_28 (
    .a(i18[28]),
    .b(sum_17[28]),
    .c(cout_18[27]),
    .cout(cout_18[28]),
    .sum(sum_18[28]));
  AL_FADD comp18_29 (
    .a(i18[29]),
    .b(sum_17[29]),
    .c(cout_18[28]),
    .cout(cout_18[29]),
    .sum(sum_18[29]));
  AL_FADD comp18_3 (
    .a(i18[3]),
    .b(sum_17[3]),
    .c(cout_18[2]),
    .cout(cout_18[3]),
    .sum(sum_18[3]));
  AL_FADD comp18_30 (
    .a(i18[30]),
    .b(sum_17[30]),
    .c(cout_18[29]),
    .cout(cout_18[30]),
    .sum(sum_18[30]));
  AL_FADD comp18_31 (
    .a(i18[31]),
    .b(sum_17[31]),
    .c(cout_18[30]),
    .cout(cout_18[31]),
    .sum(sum_18[31]));
  AL_FADD comp18_32 (
    .a(i18[32]),
    .b(sum_17[32]),
    .c(cout_18[31]),
    .cout(cout_18[32]),
    .sum(sum_18[32]));
  AL_FADD comp18_33 (
    .a(i18[33]),
    .b(sum_17[33]),
    .c(cout_18[32]),
    .cout(cout_18[33]),
    .sum(sum_18[33]));
  AL_FADD comp18_34 (
    .a(i18[34]),
    .b(sum_17[34]),
    .c(cout_18[33]),
    .cout(cout_18[34]),
    .sum(sum_18[34]));
  AL_FADD comp18_35 (
    .a(i18[35]),
    .b(sum_17[35]),
    .c(cout_18[34]),
    .cout(cout_18[35]),
    .sum(sum_18[35]));
  AL_FADD comp18_36 (
    .a(i18[36]),
    .b(sum_17[36]),
    .c(cout_18[35]),
    .cout(cout_18[36]),
    .sum(sum_18[36]));
  AL_FADD comp18_37 (
    .a(i18[37]),
    .b(sum_17[37]),
    .c(cout_18[36]),
    .cout(cout_18[37]),
    .sum(sum_18[37]));
  AL_FADD comp18_38 (
    .a(i18[38]),
    .b(sum_17[38]),
    .c(cout_18[37]),
    .cout(cout_18[38]),
    .sum(sum_18[38]));
  AL_FADD comp18_39 (
    .a(i18[39]),
    .b(sum_17[39]),
    .c(cout_18[38]),
    .cout(cout_18[39]),
    .sum(sum_18[39]));
  AL_FADD comp18_4 (
    .a(i18[4]),
    .b(sum_17[4]),
    .c(cout_18[3]),
    .cout(cout_18[4]),
    .sum(sum_18[4]));
  AL_FADD comp18_40 (
    .a(i18[40]),
    .b(sum_17[40]),
    .c(cout_18[39]),
    .cout(cout_18[40]),
    .sum(sum_18[40]));
  AL_FADD comp18_41 (
    .a(i18[41]),
    .b(sum_17[41]),
    .c(cout_18[40]),
    .cout(cout_18[41]),
    .sum(sum_18[41]));
  AL_FADD comp18_42 (
    .a(i18[42]),
    .b(sum_17[42]),
    .c(cout_18[41]),
    .cout(cout_18[42]),
    .sum(sum_18[42]));
  AL_FADD comp18_43 (
    .a(i18[43]),
    .b(sum_17[43]),
    .c(cout_18[42]),
    .cout(cout_18[43]),
    .sum(sum_18[43]));
  AL_FADD comp18_44 (
    .a(1'b0),
    .b(sum_17[44]),
    .c(cout_18[43]),
    .cout(cout_18[44]),
    .sum(sum_18[44]));
  AL_FADD comp18_45 (
    .a(1'b0),
    .b(sum_17[45]),
    .c(cout_18[44]),
    .cout(cout_18[45]),
    .sum(sum_18[45]));
  AL_FADD comp18_46 (
    .a(1'b0),
    .b(sum_17[46]),
    .c(cout_18[45]),
    .cout(cout_18[46]),
    .sum(sum_18[46]));
  AL_FADD comp18_47 (
    .a(1'b0),
    .b(sum_17[47]),
    .c(cout_18[46]),
    .cout(cout_18[47]),
    .sum(sum_18[47]));
  AL_FADD comp18_48 (
    .a(1'b0),
    .b(sum_17[48]),
    .c(cout_18[47]),
    .cout(cout_18[48]),
    .sum(sum_18[48]));
  AL_FADD comp18_49 (
    .a(1'b0),
    .b(sum_17[49]),
    .c(cout_18[48]),
    .cout(cout_18[49]),
    .sum(sum_18[49]));
  AL_FADD comp18_5 (
    .a(i18[5]),
    .b(sum_17[5]),
    .c(cout_18[4]),
    .cout(cout_18[5]),
    .sum(sum_18[5]));
  AL_FADD comp18_50 (
    .a(1'b0),
    .b(sum_17[50]),
    .c(cout_18[49]),
    .cout(cout_18[50]),
    .sum(sum_18[50]));
  AL_FADD comp18_51 (
    .a(1'b0),
    .b(sum_17[51]),
    .c(cout_18[50]),
    .cout(cout_18[51]),
    .sum(sum_18[51]));
  AL_FADD comp18_52 (
    .a(1'b0),
    .b(sum_17[52]),
    .c(cout_18[51]),
    .cout(cout_18[52]),
    .sum(sum_18[52]));
  AL_FADD comp18_53 (
    .a(1'b0),
    .b(sum_17[53]),
    .c(cout_18[52]),
    .cout(cout_18[53]),
    .sum(sum_18[53]));
  AL_FADD comp18_54 (
    .a(1'b0),
    .b(sum_17[54]),
    .c(cout_18[53]),
    .cout(cout_18[54]),
    .sum(sum_18[54]));
  AL_FADD comp18_55 (
    .a(1'b0),
    .b(sum_17[55]),
    .c(cout_18[54]),
    .cout(cout_18[55]),
    .sum(sum_18[55]));
  AL_FADD comp18_56 (
    .a(1'b0),
    .b(sum_17[56]),
    .c(cout_18[55]),
    .cout(cout_18[56]),
    .sum(sum_18[56]));
  AL_FADD comp18_57 (
    .a(1'b0),
    .b(sum_17[57]),
    .c(cout_18[56]),
    .cout(cout_18[57]),
    .sum(sum_18[57]));
  AL_FADD comp18_58 (
    .a(1'b0),
    .b(sum_17[58]),
    .c(cout_18[57]),
    .cout(cout_18[58]),
    .sum(sum_18[58]));
  AL_FADD comp18_59 (
    .a(1'b0),
    .b(sum_17[59]),
    .c(cout_18[58]),
    .cout(cout_18[59]),
    .sum(sum_18[59]));
  AL_FADD comp18_6 (
    .a(i18[6]),
    .b(sum_17[6]),
    .c(cout_18[5]),
    .cout(cout_18[6]),
    .sum(sum_18[6]));
  AL_FADD comp18_60 (
    .a(1'b0),
    .b(sum_17[60]),
    .c(cout_18[59]),
    .cout(cout_18[60]),
    .sum(sum_18[60]));
  AL_FADD comp18_61 (
    .a(1'b0),
    .b(sum_17[61]),
    .c(cout_18[60]),
    .cout(cout_18[61]),
    .sum(sum_18[61]));
  AL_FADD comp18_62 (
    .a(1'b0),
    .b(sum_17[62]),
    .c(cout_18[61]),
    .cout(cout_18[62]),
    .sum(sum_18[62]));
  AL_FADD comp18_63 (
    .a(1'b0),
    .b(sum_17[63]),
    .c(cout_18[62]),
    .cout(cout_18[63]),
    .sum(sum_18[63]));
  AL_FADD comp18_7 (
    .a(i18[7]),
    .b(sum_17[7]),
    .c(cout_18[6]),
    .cout(cout_18[7]),
    .sum(sum_18[7]));
  AL_FADD comp18_8 (
    .a(i18[8]),
    .b(sum_17[8]),
    .c(cout_18[7]),
    .cout(cout_18[8]),
    .sum(sum_18[8]));
  AL_FADD comp18_9 (
    .a(i18[9]),
    .b(sum_17[9]),
    .c(cout_18[8]),
    .cout(cout_18[9]),
    .sum(sum_18[9]));
  AL_FADD comp19_0 (
    .a(i19[0]),
    .b(sum_18[0]),
    .c(1'b0),
    .cout(cout_19[0]),
    .sum(sum_19[0]));
  AL_FADD comp19_1 (
    .a(i19[1]),
    .b(sum_18[1]),
    .c(cout_19[0]),
    .cout(cout_19[1]),
    .sum(sum_19[1]));
  AL_FADD comp19_10 (
    .a(i19[10]),
    .b(sum_18[10]),
    .c(cout_19[9]),
    .cout(cout_19[10]),
    .sum(sum_19[10]));
  AL_FADD comp19_11 (
    .a(i19[11]),
    .b(sum_18[11]),
    .c(cout_19[10]),
    .cout(cout_19[11]),
    .sum(sum_19[11]));
  AL_FADD comp19_12 (
    .a(i19[12]),
    .b(sum_18[12]),
    .c(cout_19[11]),
    .cout(cout_19[12]),
    .sum(sum_19[12]));
  AL_FADD comp19_13 (
    .a(i19[13]),
    .b(sum_18[13]),
    .c(cout_19[12]),
    .cout(cout_19[13]),
    .sum(sum_19[13]));
  AL_FADD comp19_14 (
    .a(i19[14]),
    .b(sum_18[14]),
    .c(cout_19[13]),
    .cout(cout_19[14]),
    .sum(sum_19[14]));
  AL_FADD comp19_15 (
    .a(i19[15]),
    .b(sum_18[15]),
    .c(cout_19[14]),
    .cout(cout_19[15]),
    .sum(sum_19[15]));
  AL_FADD comp19_16 (
    .a(i19[16]),
    .b(sum_18[16]),
    .c(cout_19[15]),
    .cout(cout_19[16]),
    .sum(sum_19[16]));
  AL_FADD comp19_17 (
    .a(i19[17]),
    .b(sum_18[17]),
    .c(cout_19[16]),
    .cout(cout_19[17]),
    .sum(sum_19[17]));
  AL_FADD comp19_18 (
    .a(i19[18]),
    .b(sum_18[18]),
    .c(cout_19[17]),
    .cout(cout_19[18]),
    .sum(sum_19[18]));
  AL_FADD comp19_19 (
    .a(i19[19]),
    .b(sum_18[19]),
    .c(cout_19[18]),
    .cout(cout_19[19]),
    .sum(sum_19[19]));
  AL_FADD comp19_2 (
    .a(i19[2]),
    .b(sum_18[2]),
    .c(cout_19[1]),
    .cout(cout_19[2]),
    .sum(sum_19[2]));
  AL_FADD comp19_20 (
    .a(i19[20]),
    .b(sum_18[20]),
    .c(cout_19[19]),
    .cout(cout_19[20]),
    .sum(sum_19[20]));
  AL_FADD comp19_21 (
    .a(i19[21]),
    .b(sum_18[21]),
    .c(cout_19[20]),
    .cout(cout_19[21]),
    .sum(sum_19[21]));
  AL_FADD comp19_22 (
    .a(i19[22]),
    .b(sum_18[22]),
    .c(cout_19[21]),
    .cout(cout_19[22]),
    .sum(sum_19[22]));
  AL_FADD comp19_23 (
    .a(i19[23]),
    .b(sum_18[23]),
    .c(cout_19[22]),
    .cout(cout_19[23]),
    .sum(sum_19[23]));
  AL_FADD comp19_24 (
    .a(i19[24]),
    .b(sum_18[24]),
    .c(cout_19[23]),
    .cout(cout_19[24]),
    .sum(sum_19[24]));
  AL_FADD comp19_25 (
    .a(i19[25]),
    .b(sum_18[25]),
    .c(cout_19[24]),
    .cout(cout_19[25]),
    .sum(sum_19[25]));
  AL_FADD comp19_26 (
    .a(i19[26]),
    .b(sum_18[26]),
    .c(cout_19[25]),
    .cout(cout_19[26]),
    .sum(sum_19[26]));
  AL_FADD comp19_27 (
    .a(i19[27]),
    .b(sum_18[27]),
    .c(cout_19[26]),
    .cout(cout_19[27]),
    .sum(sum_19[27]));
  AL_FADD comp19_28 (
    .a(i19[28]),
    .b(sum_18[28]),
    .c(cout_19[27]),
    .cout(cout_19[28]),
    .sum(sum_19[28]));
  AL_FADD comp19_29 (
    .a(i19[29]),
    .b(sum_18[29]),
    .c(cout_19[28]),
    .cout(cout_19[29]),
    .sum(sum_19[29]));
  AL_FADD comp19_3 (
    .a(i19[3]),
    .b(sum_18[3]),
    .c(cout_19[2]),
    .cout(cout_19[3]),
    .sum(sum_19[3]));
  AL_FADD comp19_30 (
    .a(i19[30]),
    .b(sum_18[30]),
    .c(cout_19[29]),
    .cout(cout_19[30]),
    .sum(sum_19[30]));
  AL_FADD comp19_31 (
    .a(i19[31]),
    .b(sum_18[31]),
    .c(cout_19[30]),
    .cout(cout_19[31]),
    .sum(sum_19[31]));
  AL_FADD comp19_32 (
    .a(i19[32]),
    .b(sum_18[32]),
    .c(cout_19[31]),
    .cout(cout_19[32]),
    .sum(sum_19[32]));
  AL_FADD comp19_33 (
    .a(i19[33]),
    .b(sum_18[33]),
    .c(cout_19[32]),
    .cout(cout_19[33]),
    .sum(sum_19[33]));
  AL_FADD comp19_34 (
    .a(i19[34]),
    .b(sum_18[34]),
    .c(cout_19[33]),
    .cout(cout_19[34]),
    .sum(sum_19[34]));
  AL_FADD comp19_35 (
    .a(i19[35]),
    .b(sum_18[35]),
    .c(cout_19[34]),
    .cout(cout_19[35]),
    .sum(sum_19[35]));
  AL_FADD comp19_36 (
    .a(i19[36]),
    .b(sum_18[36]),
    .c(cout_19[35]),
    .cout(cout_19[36]),
    .sum(sum_19[36]));
  AL_FADD comp19_37 (
    .a(i19[37]),
    .b(sum_18[37]),
    .c(cout_19[36]),
    .cout(cout_19[37]),
    .sum(sum_19[37]));
  AL_FADD comp19_38 (
    .a(i19[38]),
    .b(sum_18[38]),
    .c(cout_19[37]),
    .cout(cout_19[38]),
    .sum(sum_19[38]));
  AL_FADD comp19_39 (
    .a(i19[39]),
    .b(sum_18[39]),
    .c(cout_19[38]),
    .cout(cout_19[39]),
    .sum(sum_19[39]));
  AL_FADD comp19_4 (
    .a(i19[4]),
    .b(sum_18[4]),
    .c(cout_19[3]),
    .cout(cout_19[4]),
    .sum(sum_19[4]));
  AL_FADD comp19_40 (
    .a(i19[40]),
    .b(sum_18[40]),
    .c(cout_19[39]),
    .cout(cout_19[40]),
    .sum(sum_19[40]));
  AL_FADD comp19_41 (
    .a(i19[41]),
    .b(sum_18[41]),
    .c(cout_19[40]),
    .cout(cout_19[41]),
    .sum(sum_19[41]));
  AL_FADD comp19_42 (
    .a(i19[42]),
    .b(sum_18[42]),
    .c(cout_19[41]),
    .cout(cout_19[42]),
    .sum(sum_19[42]));
  AL_FADD comp19_43 (
    .a(1'b0),
    .b(sum_18[43]),
    .c(cout_19[42]),
    .cout(cout_19[43]),
    .sum(sum_19[43]));
  AL_FADD comp19_44 (
    .a(1'b0),
    .b(sum_18[44]),
    .c(cout_19[43]),
    .cout(cout_19[44]),
    .sum(sum_19[44]));
  AL_FADD comp19_45 (
    .a(1'b0),
    .b(sum_18[45]),
    .c(cout_19[44]),
    .cout(cout_19[45]),
    .sum(sum_19[45]));
  AL_FADD comp19_46 (
    .a(1'b0),
    .b(sum_18[46]),
    .c(cout_19[45]),
    .cout(cout_19[46]),
    .sum(sum_19[46]));
  AL_FADD comp19_47 (
    .a(1'b0),
    .b(sum_18[47]),
    .c(cout_19[46]),
    .cout(cout_19[47]),
    .sum(sum_19[47]));
  AL_FADD comp19_48 (
    .a(1'b0),
    .b(sum_18[48]),
    .c(cout_19[47]),
    .cout(cout_19[48]),
    .sum(sum_19[48]));
  AL_FADD comp19_49 (
    .a(1'b0),
    .b(sum_18[49]),
    .c(cout_19[48]),
    .cout(cout_19[49]),
    .sum(sum_19[49]));
  AL_FADD comp19_5 (
    .a(i19[5]),
    .b(sum_18[5]),
    .c(cout_19[4]),
    .cout(cout_19[5]),
    .sum(sum_19[5]));
  AL_FADD comp19_50 (
    .a(1'b0),
    .b(sum_18[50]),
    .c(cout_19[49]),
    .cout(cout_19[50]),
    .sum(sum_19[50]));
  AL_FADD comp19_51 (
    .a(1'b0),
    .b(sum_18[51]),
    .c(cout_19[50]),
    .cout(cout_19[51]),
    .sum(sum_19[51]));
  AL_FADD comp19_52 (
    .a(1'b0),
    .b(sum_18[52]),
    .c(cout_19[51]),
    .cout(cout_19[52]),
    .sum(sum_19[52]));
  AL_FADD comp19_53 (
    .a(1'b0),
    .b(sum_18[53]),
    .c(cout_19[52]),
    .cout(cout_19[53]),
    .sum(sum_19[53]));
  AL_FADD comp19_54 (
    .a(1'b0),
    .b(sum_18[54]),
    .c(cout_19[53]),
    .cout(cout_19[54]),
    .sum(sum_19[54]));
  AL_FADD comp19_55 (
    .a(1'b0),
    .b(sum_18[55]),
    .c(cout_19[54]),
    .cout(cout_19[55]),
    .sum(sum_19[55]));
  AL_FADD comp19_56 (
    .a(1'b0),
    .b(sum_18[56]),
    .c(cout_19[55]),
    .cout(cout_19[56]),
    .sum(sum_19[56]));
  AL_FADD comp19_57 (
    .a(1'b0),
    .b(sum_18[57]),
    .c(cout_19[56]),
    .cout(cout_19[57]),
    .sum(sum_19[57]));
  AL_FADD comp19_58 (
    .a(1'b0),
    .b(sum_18[58]),
    .c(cout_19[57]),
    .cout(cout_19[58]),
    .sum(sum_19[58]));
  AL_FADD comp19_59 (
    .a(1'b0),
    .b(sum_18[59]),
    .c(cout_19[58]),
    .cout(cout_19[59]),
    .sum(sum_19[59]));
  AL_FADD comp19_6 (
    .a(i19[6]),
    .b(sum_18[6]),
    .c(cout_19[5]),
    .cout(cout_19[6]),
    .sum(sum_19[6]));
  AL_FADD comp19_60 (
    .a(1'b0),
    .b(sum_18[60]),
    .c(cout_19[59]),
    .cout(cout_19[60]),
    .sum(sum_19[60]));
  AL_FADD comp19_61 (
    .a(1'b0),
    .b(sum_18[61]),
    .c(cout_19[60]),
    .cout(cout_19[61]),
    .sum(sum_19[61]));
  AL_FADD comp19_62 (
    .a(1'b0),
    .b(sum_18[62]),
    .c(cout_19[61]),
    .cout(cout_19[62]),
    .sum(sum_19[62]));
  AL_FADD comp19_63 (
    .a(1'b0),
    .b(sum_18[63]),
    .c(cout_19[62]),
    .cout(cout_19[63]),
    .sum(sum_19[63]));
  AL_FADD comp19_7 (
    .a(i19[7]),
    .b(sum_18[7]),
    .c(cout_19[6]),
    .cout(cout_19[7]),
    .sum(sum_19[7]));
  AL_FADD comp19_8 (
    .a(i19[8]),
    .b(sum_18[8]),
    .c(cout_19[7]),
    .cout(cout_19[8]),
    .sum(sum_19[8]));
  AL_FADD comp19_9 (
    .a(i19[9]),
    .b(sum_18[9]),
    .c(cout_19[8]),
    .cout(cout_19[9]),
    .sum(sum_19[9]));
  AL_FADD comp1_0 (
    .a(i1[0]),
    .b(i0[0]),
    .c(1'b0),
    .cout(cout_1[0]),
    .sum(sum_1[0]));
  AL_FADD comp1_1 (
    .a(i1[1]),
    .b(i0[1]),
    .c(cout_1[0]),
    .cout(cout_1[1]),
    .sum(sum_1[1]));
  AL_FADD comp1_10 (
    .a(i1[10]),
    .b(i0[10]),
    .c(cout_1[9]),
    .cout(cout_1[10]),
    .sum(sum_1[10]));
  AL_FADD comp1_11 (
    .a(i1[11]),
    .b(i0[11]),
    .c(cout_1[10]),
    .cout(cout_1[11]),
    .sum(sum_1[11]));
  AL_FADD comp1_12 (
    .a(i1[12]),
    .b(i0[12]),
    .c(cout_1[11]),
    .cout(cout_1[12]),
    .sum(sum_1[12]));
  AL_FADD comp1_13 (
    .a(i1[13]),
    .b(i0[13]),
    .c(cout_1[12]),
    .cout(cout_1[13]),
    .sum(sum_1[13]));
  AL_FADD comp1_14 (
    .a(i1[14]),
    .b(i0[14]),
    .c(cout_1[13]),
    .cout(cout_1[14]),
    .sum(sum_1[14]));
  AL_FADD comp1_15 (
    .a(i1[15]),
    .b(i0[15]),
    .c(cout_1[14]),
    .cout(cout_1[15]),
    .sum(sum_1[15]));
  AL_FADD comp1_16 (
    .a(i1[16]),
    .b(i0[16]),
    .c(cout_1[15]),
    .cout(cout_1[16]),
    .sum(sum_1[16]));
  AL_FADD comp1_17 (
    .a(i1[17]),
    .b(i0[17]),
    .c(cout_1[16]),
    .cout(cout_1[17]),
    .sum(sum_1[17]));
  AL_FADD comp1_18 (
    .a(i1[18]),
    .b(i0[18]),
    .c(cout_1[17]),
    .cout(cout_1[18]),
    .sum(sum_1[18]));
  AL_FADD comp1_19 (
    .a(i1[19]),
    .b(i0[19]),
    .c(cout_1[18]),
    .cout(cout_1[19]),
    .sum(sum_1[19]));
  AL_FADD comp1_2 (
    .a(i1[2]),
    .b(i0[2]),
    .c(cout_1[1]),
    .cout(cout_1[2]),
    .sum(sum_1[2]));
  AL_FADD comp1_20 (
    .a(i1[20]),
    .b(i0[20]),
    .c(cout_1[19]),
    .cout(cout_1[20]),
    .sum(sum_1[20]));
  AL_FADD comp1_21 (
    .a(i1[21]),
    .b(i0[21]),
    .c(cout_1[20]),
    .cout(cout_1[21]),
    .sum(sum_1[21]));
  AL_FADD comp1_22 (
    .a(i1[22]),
    .b(i0[22]),
    .c(cout_1[21]),
    .cout(cout_1[22]),
    .sum(sum_1[22]));
  AL_FADD comp1_23 (
    .a(i1[23]),
    .b(i0[23]),
    .c(cout_1[22]),
    .cout(cout_1[23]),
    .sum(sum_1[23]));
  AL_FADD comp1_24 (
    .a(i1[24]),
    .b(i0[24]),
    .c(cout_1[23]),
    .cout(cout_1[24]),
    .sum(sum_1[24]));
  AL_FADD comp1_25 (
    .a(i1[25]),
    .b(i0[25]),
    .c(cout_1[24]),
    .cout(cout_1[25]),
    .sum(sum_1[25]));
  AL_FADD comp1_26 (
    .a(i1[26]),
    .b(i0[26]),
    .c(cout_1[25]),
    .cout(cout_1[26]),
    .sum(sum_1[26]));
  AL_FADD comp1_27 (
    .a(i1[27]),
    .b(i0[27]),
    .c(cout_1[26]),
    .cout(cout_1[27]),
    .sum(sum_1[27]));
  AL_FADD comp1_28 (
    .a(i1[28]),
    .b(i0[28]),
    .c(cout_1[27]),
    .cout(cout_1[28]),
    .sum(sum_1[28]));
  AL_FADD comp1_29 (
    .a(i1[29]),
    .b(i0[29]),
    .c(cout_1[28]),
    .cout(cout_1[29]),
    .sum(sum_1[29]));
  AL_FADD comp1_3 (
    .a(i1[3]),
    .b(i0[3]),
    .c(cout_1[2]),
    .cout(cout_1[3]),
    .sum(sum_1[3]));
  AL_FADD comp1_30 (
    .a(i1[30]),
    .b(i0[30]),
    .c(cout_1[29]),
    .cout(cout_1[30]),
    .sum(sum_1[30]));
  AL_FADD comp1_31 (
    .a(i1[31]),
    .b(i0[31]),
    .c(cout_1[30]),
    .cout(cout_1[31]),
    .sum(sum_1[31]));
  AL_FADD comp1_32 (
    .a(i1[32]),
    .b(i0[32]),
    .c(cout_1[31]),
    .cout(cout_1[32]),
    .sum(sum_1[32]));
  AL_FADD comp1_33 (
    .a(i1[33]),
    .b(i0[33]),
    .c(cout_1[32]),
    .cout(cout_1[33]),
    .sum(sum_1[33]));
  AL_FADD comp1_34 (
    .a(i1[34]),
    .b(i0[34]),
    .c(cout_1[33]),
    .cout(cout_1[34]),
    .sum(sum_1[34]));
  AL_FADD comp1_35 (
    .a(i1[35]),
    .b(i0[35]),
    .c(cout_1[34]),
    .cout(cout_1[35]),
    .sum(sum_1[35]));
  AL_FADD comp1_36 (
    .a(i1[36]),
    .b(i0[36]),
    .c(cout_1[35]),
    .cout(cout_1[36]),
    .sum(sum_1[36]));
  AL_FADD comp1_37 (
    .a(i1[37]),
    .b(i0[37]),
    .c(cout_1[36]),
    .cout(cout_1[37]),
    .sum(sum_1[37]));
  AL_FADD comp1_38 (
    .a(i1[38]),
    .b(i0[38]),
    .c(cout_1[37]),
    .cout(cout_1[38]),
    .sum(sum_1[38]));
  AL_FADD comp1_39 (
    .a(i1[39]),
    .b(i0[39]),
    .c(cout_1[38]),
    .cout(cout_1[39]),
    .sum(sum_1[39]));
  AL_FADD comp1_4 (
    .a(i1[4]),
    .b(i0[4]),
    .c(cout_1[3]),
    .cout(cout_1[4]),
    .sum(sum_1[4]));
  AL_FADD comp1_40 (
    .a(i1[40]),
    .b(i0[40]),
    .c(cout_1[39]),
    .cout(cout_1[40]),
    .sum(sum_1[40]));
  AL_FADD comp1_41 (
    .a(i1[41]),
    .b(i0[41]),
    .c(cout_1[40]),
    .cout(cout_1[41]),
    .sum(sum_1[41]));
  AL_FADD comp1_42 (
    .a(i1[42]),
    .b(i0[42]),
    .c(cout_1[41]),
    .cout(cout_1[42]),
    .sum(sum_1[42]));
  AL_FADD comp1_43 (
    .a(i1[43]),
    .b(i0[43]),
    .c(cout_1[42]),
    .cout(cout_1[43]),
    .sum(sum_1[43]));
  AL_FADD comp1_44 (
    .a(i1[44]),
    .b(i0[44]),
    .c(cout_1[43]),
    .cout(cout_1[44]),
    .sum(sum_1[44]));
  AL_FADD comp1_45 (
    .a(i1[45]),
    .b(i0[45]),
    .c(cout_1[44]),
    .cout(cout_1[45]),
    .sum(sum_1[45]));
  AL_FADD comp1_46 (
    .a(i1[46]),
    .b(i0[46]),
    .c(cout_1[45]),
    .cout(cout_1[46]),
    .sum(sum_1[46]));
  AL_FADD comp1_47 (
    .a(i1[47]),
    .b(i0[47]),
    .c(cout_1[46]),
    .cout(cout_1[47]),
    .sum(sum_1[47]));
  AL_FADD comp1_48 (
    .a(i1[48]),
    .b(i0[48]),
    .c(cout_1[47]),
    .cout(cout_1[48]),
    .sum(sum_1[48]));
  AL_FADD comp1_49 (
    .a(i1[49]),
    .b(i0[49]),
    .c(cout_1[48]),
    .cout(cout_1[49]),
    .sum(sum_1[49]));
  AL_FADD comp1_5 (
    .a(i1[5]),
    .b(i0[5]),
    .c(cout_1[4]),
    .cout(cout_1[5]),
    .sum(sum_1[5]));
  AL_FADD comp1_50 (
    .a(i1[50]),
    .b(i0[50]),
    .c(cout_1[49]),
    .cout(cout_1[50]),
    .sum(sum_1[50]));
  AL_FADD comp1_51 (
    .a(i1[51]),
    .b(i0[51]),
    .c(cout_1[50]),
    .cout(cout_1[51]),
    .sum(sum_1[51]));
  AL_FADD comp1_52 (
    .a(i1[52]),
    .b(i0[52]),
    .c(cout_1[51]),
    .cout(cout_1[52]),
    .sum(sum_1[52]));
  AL_FADD comp1_53 (
    .a(i1[53]),
    .b(i0[53]),
    .c(cout_1[52]),
    .cout(cout_1[53]),
    .sum(sum_1[53]));
  AL_FADD comp1_54 (
    .a(i1[54]),
    .b(i0[54]),
    .c(cout_1[53]),
    .cout(cout_1[54]),
    .sum(sum_1[54]));
  AL_FADD comp1_55 (
    .a(i1[55]),
    .b(i0[55]),
    .c(cout_1[54]),
    .cout(cout_1[55]),
    .sum(sum_1[55]));
  AL_FADD comp1_56 (
    .a(i1[56]),
    .b(i0[56]),
    .c(cout_1[55]),
    .cout(cout_1[56]),
    .sum(sum_1[56]));
  AL_FADD comp1_57 (
    .a(i1[57]),
    .b(i0[57]),
    .c(cout_1[56]),
    .cout(cout_1[57]),
    .sum(sum_1[57]));
  AL_FADD comp1_58 (
    .a(i1[58]),
    .b(i0[58]),
    .c(cout_1[57]),
    .cout(cout_1[58]),
    .sum(sum_1[58]));
  AL_FADD comp1_59 (
    .a(i1[59]),
    .b(i0[59]),
    .c(cout_1[58]),
    .cout(cout_1[59]),
    .sum(sum_1[59]));
  AL_FADD comp1_6 (
    .a(i1[6]),
    .b(i0[6]),
    .c(cout_1[5]),
    .cout(cout_1[6]),
    .sum(sum_1[6]));
  AL_FADD comp1_60 (
    .a(i1[60]),
    .b(i0[60]),
    .c(cout_1[59]),
    .cout(cout_1[60]),
    .sum(sum_1[60]));
  AL_FADD comp1_61 (
    .a(1'b0),
    .b(i0[61]),
    .c(cout_1[60]),
    .cout(cout_1[61]),
    .sum(sum_1[61]));
  AL_FADD comp1_62 (
    .a(1'b0),
    .b(i0[62]),
    .c(cout_1[61]),
    .cout(cout_1[62]),
    .sum(sum_1[62]));
  AL_FADD comp1_63 (
    .a(1'b0),
    .b(i0[63]),
    .c(cout_1[62]),
    .cout(cout_1[63]),
    .sum(sum_1[63]));
  AL_FADD comp1_7 (
    .a(i1[7]),
    .b(i0[7]),
    .c(cout_1[6]),
    .cout(cout_1[7]),
    .sum(sum_1[7]));
  AL_FADD comp1_8 (
    .a(i1[8]),
    .b(i0[8]),
    .c(cout_1[7]),
    .cout(cout_1[8]),
    .sum(sum_1[8]));
  AL_FADD comp1_9 (
    .a(i1[9]),
    .b(i0[9]),
    .c(cout_1[8]),
    .cout(cout_1[9]),
    .sum(sum_1[9]));
  AL_FADD comp20_0 (
    .a(i20[0]),
    .b(sum_19[0]),
    .c(1'b0),
    .cout(cout_20[0]),
    .sum(sum_20[0]));
  AL_FADD comp20_1 (
    .a(i20[1]),
    .b(sum_19[1]),
    .c(cout_20[0]),
    .cout(cout_20[1]),
    .sum(sum_20[1]));
  AL_FADD comp20_10 (
    .a(i20[10]),
    .b(sum_19[10]),
    .c(cout_20[9]),
    .cout(cout_20[10]),
    .sum(sum_20[10]));
  AL_FADD comp20_11 (
    .a(i20[11]),
    .b(sum_19[11]),
    .c(cout_20[10]),
    .cout(cout_20[11]),
    .sum(sum_20[11]));
  AL_FADD comp20_12 (
    .a(i20[12]),
    .b(sum_19[12]),
    .c(cout_20[11]),
    .cout(cout_20[12]),
    .sum(sum_20[12]));
  AL_FADD comp20_13 (
    .a(i20[13]),
    .b(sum_19[13]),
    .c(cout_20[12]),
    .cout(cout_20[13]),
    .sum(sum_20[13]));
  AL_FADD comp20_14 (
    .a(i20[14]),
    .b(sum_19[14]),
    .c(cout_20[13]),
    .cout(cout_20[14]),
    .sum(sum_20[14]));
  AL_FADD comp20_15 (
    .a(i20[15]),
    .b(sum_19[15]),
    .c(cout_20[14]),
    .cout(cout_20[15]),
    .sum(sum_20[15]));
  AL_FADD comp20_16 (
    .a(i20[16]),
    .b(sum_19[16]),
    .c(cout_20[15]),
    .cout(cout_20[16]),
    .sum(sum_20[16]));
  AL_FADD comp20_17 (
    .a(i20[17]),
    .b(sum_19[17]),
    .c(cout_20[16]),
    .cout(cout_20[17]),
    .sum(sum_20[17]));
  AL_FADD comp20_18 (
    .a(i20[18]),
    .b(sum_19[18]),
    .c(cout_20[17]),
    .cout(cout_20[18]),
    .sum(sum_20[18]));
  AL_FADD comp20_19 (
    .a(i20[19]),
    .b(sum_19[19]),
    .c(cout_20[18]),
    .cout(cout_20[19]),
    .sum(sum_20[19]));
  AL_FADD comp20_2 (
    .a(i20[2]),
    .b(sum_19[2]),
    .c(cout_20[1]),
    .cout(cout_20[2]),
    .sum(sum_20[2]));
  AL_FADD comp20_20 (
    .a(i20[20]),
    .b(sum_19[20]),
    .c(cout_20[19]),
    .cout(cout_20[20]),
    .sum(sum_20[20]));
  AL_FADD comp20_21 (
    .a(i20[21]),
    .b(sum_19[21]),
    .c(cout_20[20]),
    .cout(cout_20[21]),
    .sum(sum_20[21]));
  AL_FADD comp20_22 (
    .a(i20[22]),
    .b(sum_19[22]),
    .c(cout_20[21]),
    .cout(cout_20[22]),
    .sum(sum_20[22]));
  AL_FADD comp20_23 (
    .a(i20[23]),
    .b(sum_19[23]),
    .c(cout_20[22]),
    .cout(cout_20[23]),
    .sum(sum_20[23]));
  AL_FADD comp20_24 (
    .a(i20[24]),
    .b(sum_19[24]),
    .c(cout_20[23]),
    .cout(cout_20[24]),
    .sum(sum_20[24]));
  AL_FADD comp20_25 (
    .a(i20[25]),
    .b(sum_19[25]),
    .c(cout_20[24]),
    .cout(cout_20[25]),
    .sum(sum_20[25]));
  AL_FADD comp20_26 (
    .a(i20[26]),
    .b(sum_19[26]),
    .c(cout_20[25]),
    .cout(cout_20[26]),
    .sum(sum_20[26]));
  AL_FADD comp20_27 (
    .a(i20[27]),
    .b(sum_19[27]),
    .c(cout_20[26]),
    .cout(cout_20[27]),
    .sum(sum_20[27]));
  AL_FADD comp20_28 (
    .a(i20[28]),
    .b(sum_19[28]),
    .c(cout_20[27]),
    .cout(cout_20[28]),
    .sum(sum_20[28]));
  AL_FADD comp20_29 (
    .a(i20[29]),
    .b(sum_19[29]),
    .c(cout_20[28]),
    .cout(cout_20[29]),
    .sum(sum_20[29]));
  AL_FADD comp20_3 (
    .a(i20[3]),
    .b(sum_19[3]),
    .c(cout_20[2]),
    .cout(cout_20[3]),
    .sum(sum_20[3]));
  AL_FADD comp20_30 (
    .a(i20[30]),
    .b(sum_19[30]),
    .c(cout_20[29]),
    .cout(cout_20[30]),
    .sum(sum_20[30]));
  AL_FADD comp20_31 (
    .a(i20[31]),
    .b(sum_19[31]),
    .c(cout_20[30]),
    .cout(cout_20[31]),
    .sum(sum_20[31]));
  AL_FADD comp20_32 (
    .a(i20[32]),
    .b(sum_19[32]),
    .c(cout_20[31]),
    .cout(cout_20[32]),
    .sum(sum_20[32]));
  AL_FADD comp20_33 (
    .a(i20[33]),
    .b(sum_19[33]),
    .c(cout_20[32]),
    .cout(cout_20[33]),
    .sum(sum_20[33]));
  AL_FADD comp20_34 (
    .a(i20[34]),
    .b(sum_19[34]),
    .c(cout_20[33]),
    .cout(cout_20[34]),
    .sum(sum_20[34]));
  AL_FADD comp20_35 (
    .a(i20[35]),
    .b(sum_19[35]),
    .c(cout_20[34]),
    .cout(cout_20[35]),
    .sum(sum_20[35]));
  AL_FADD comp20_36 (
    .a(i20[36]),
    .b(sum_19[36]),
    .c(cout_20[35]),
    .cout(cout_20[36]),
    .sum(sum_20[36]));
  AL_FADD comp20_37 (
    .a(i20[37]),
    .b(sum_19[37]),
    .c(cout_20[36]),
    .cout(cout_20[37]),
    .sum(sum_20[37]));
  AL_FADD comp20_38 (
    .a(i20[38]),
    .b(sum_19[38]),
    .c(cout_20[37]),
    .cout(cout_20[38]),
    .sum(sum_20[38]));
  AL_FADD comp20_39 (
    .a(i20[39]),
    .b(sum_19[39]),
    .c(cout_20[38]),
    .cout(cout_20[39]),
    .sum(sum_20[39]));
  AL_FADD comp20_4 (
    .a(i20[4]),
    .b(sum_19[4]),
    .c(cout_20[3]),
    .cout(cout_20[4]),
    .sum(sum_20[4]));
  AL_FADD comp20_40 (
    .a(i20[40]),
    .b(sum_19[40]),
    .c(cout_20[39]),
    .cout(cout_20[40]),
    .sum(sum_20[40]));
  AL_FADD comp20_41 (
    .a(i20[41]),
    .b(sum_19[41]),
    .c(cout_20[40]),
    .cout(cout_20[41]),
    .sum(sum_20[41]));
  AL_FADD comp20_42 (
    .a(1'b0),
    .b(sum_19[42]),
    .c(cout_20[41]),
    .cout(cout_20[42]),
    .sum(sum_20[42]));
  AL_FADD comp20_43 (
    .a(1'b0),
    .b(sum_19[43]),
    .c(cout_20[42]),
    .cout(cout_20[43]),
    .sum(sum_20[43]));
  AL_FADD comp20_44 (
    .a(1'b0),
    .b(sum_19[44]),
    .c(cout_20[43]),
    .cout(cout_20[44]),
    .sum(sum_20[44]));
  AL_FADD comp20_45 (
    .a(1'b0),
    .b(sum_19[45]),
    .c(cout_20[44]),
    .cout(cout_20[45]),
    .sum(sum_20[45]));
  AL_FADD comp20_46 (
    .a(1'b0),
    .b(sum_19[46]),
    .c(cout_20[45]),
    .cout(cout_20[46]),
    .sum(sum_20[46]));
  AL_FADD comp20_47 (
    .a(1'b0),
    .b(sum_19[47]),
    .c(cout_20[46]),
    .cout(cout_20[47]),
    .sum(sum_20[47]));
  AL_FADD comp20_48 (
    .a(1'b0),
    .b(sum_19[48]),
    .c(cout_20[47]),
    .cout(cout_20[48]),
    .sum(sum_20[48]));
  AL_FADD comp20_49 (
    .a(1'b0),
    .b(sum_19[49]),
    .c(cout_20[48]),
    .cout(cout_20[49]),
    .sum(sum_20[49]));
  AL_FADD comp20_5 (
    .a(i20[5]),
    .b(sum_19[5]),
    .c(cout_20[4]),
    .cout(cout_20[5]),
    .sum(sum_20[5]));
  AL_FADD comp20_50 (
    .a(1'b0),
    .b(sum_19[50]),
    .c(cout_20[49]),
    .cout(cout_20[50]),
    .sum(sum_20[50]));
  AL_FADD comp20_51 (
    .a(1'b0),
    .b(sum_19[51]),
    .c(cout_20[50]),
    .cout(cout_20[51]),
    .sum(sum_20[51]));
  AL_FADD comp20_52 (
    .a(1'b0),
    .b(sum_19[52]),
    .c(cout_20[51]),
    .cout(cout_20[52]),
    .sum(sum_20[52]));
  AL_FADD comp20_53 (
    .a(1'b0),
    .b(sum_19[53]),
    .c(cout_20[52]),
    .cout(cout_20[53]),
    .sum(sum_20[53]));
  AL_FADD comp20_54 (
    .a(1'b0),
    .b(sum_19[54]),
    .c(cout_20[53]),
    .cout(cout_20[54]),
    .sum(sum_20[54]));
  AL_FADD comp20_55 (
    .a(1'b0),
    .b(sum_19[55]),
    .c(cout_20[54]),
    .cout(cout_20[55]),
    .sum(sum_20[55]));
  AL_FADD comp20_56 (
    .a(1'b0),
    .b(sum_19[56]),
    .c(cout_20[55]),
    .cout(cout_20[56]),
    .sum(sum_20[56]));
  AL_FADD comp20_57 (
    .a(1'b0),
    .b(sum_19[57]),
    .c(cout_20[56]),
    .cout(cout_20[57]),
    .sum(sum_20[57]));
  AL_FADD comp20_58 (
    .a(1'b0),
    .b(sum_19[58]),
    .c(cout_20[57]),
    .cout(cout_20[58]),
    .sum(sum_20[58]));
  AL_FADD comp20_59 (
    .a(1'b0),
    .b(sum_19[59]),
    .c(cout_20[58]),
    .cout(cout_20[59]),
    .sum(sum_20[59]));
  AL_FADD comp20_6 (
    .a(i20[6]),
    .b(sum_19[6]),
    .c(cout_20[5]),
    .cout(cout_20[6]),
    .sum(sum_20[6]));
  AL_FADD comp20_60 (
    .a(1'b0),
    .b(sum_19[60]),
    .c(cout_20[59]),
    .cout(cout_20[60]),
    .sum(sum_20[60]));
  AL_FADD comp20_61 (
    .a(1'b0),
    .b(sum_19[61]),
    .c(cout_20[60]),
    .cout(cout_20[61]),
    .sum(sum_20[61]));
  AL_FADD comp20_62 (
    .a(1'b0),
    .b(sum_19[62]),
    .c(cout_20[61]),
    .cout(cout_20[62]),
    .sum(sum_20[62]));
  AL_FADD comp20_63 (
    .a(1'b0),
    .b(sum_19[63]),
    .c(cout_20[62]),
    .cout(cout_20[63]),
    .sum(sum_20[63]));
  AL_FADD comp20_7 (
    .a(i20[7]),
    .b(sum_19[7]),
    .c(cout_20[6]),
    .cout(cout_20[7]),
    .sum(sum_20[7]));
  AL_FADD comp20_8 (
    .a(i20[8]),
    .b(sum_19[8]),
    .c(cout_20[7]),
    .cout(cout_20[8]),
    .sum(sum_20[8]));
  AL_FADD comp20_9 (
    .a(i20[9]),
    .b(sum_19[9]),
    .c(cout_20[8]),
    .cout(cout_20[9]),
    .sum(sum_20[9]));
  AL_FADD comp21_0 (
    .a(i21[0]),
    .b(sum_20[0]),
    .c(1'b0),
    .cout(cout_21[0]),
    .sum(sum_21[0]));
  AL_FADD comp21_1 (
    .a(i21[1]),
    .b(sum_20[1]),
    .c(cout_21[0]),
    .cout(cout_21[1]),
    .sum(sum_21[1]));
  AL_FADD comp21_10 (
    .a(i21[10]),
    .b(sum_20[10]),
    .c(cout_21[9]),
    .cout(cout_21[10]),
    .sum(sum_21[10]));
  AL_FADD comp21_11 (
    .a(i21[11]),
    .b(sum_20[11]),
    .c(cout_21[10]),
    .cout(cout_21[11]),
    .sum(sum_21[11]));
  AL_FADD comp21_12 (
    .a(i21[12]),
    .b(sum_20[12]),
    .c(cout_21[11]),
    .cout(cout_21[12]),
    .sum(sum_21[12]));
  AL_FADD comp21_13 (
    .a(i21[13]),
    .b(sum_20[13]),
    .c(cout_21[12]),
    .cout(cout_21[13]),
    .sum(sum_21[13]));
  AL_FADD comp21_14 (
    .a(i21[14]),
    .b(sum_20[14]),
    .c(cout_21[13]),
    .cout(cout_21[14]),
    .sum(sum_21[14]));
  AL_FADD comp21_15 (
    .a(i21[15]),
    .b(sum_20[15]),
    .c(cout_21[14]),
    .cout(cout_21[15]),
    .sum(sum_21[15]));
  AL_FADD comp21_16 (
    .a(i21[16]),
    .b(sum_20[16]),
    .c(cout_21[15]),
    .cout(cout_21[16]),
    .sum(sum_21[16]));
  AL_FADD comp21_17 (
    .a(i21[17]),
    .b(sum_20[17]),
    .c(cout_21[16]),
    .cout(cout_21[17]),
    .sum(sum_21[17]));
  AL_FADD comp21_18 (
    .a(i21[18]),
    .b(sum_20[18]),
    .c(cout_21[17]),
    .cout(cout_21[18]),
    .sum(sum_21[18]));
  AL_FADD comp21_19 (
    .a(i21[19]),
    .b(sum_20[19]),
    .c(cout_21[18]),
    .cout(cout_21[19]),
    .sum(sum_21[19]));
  AL_FADD comp21_2 (
    .a(i21[2]),
    .b(sum_20[2]),
    .c(cout_21[1]),
    .cout(cout_21[2]),
    .sum(sum_21[2]));
  AL_FADD comp21_20 (
    .a(i21[20]),
    .b(sum_20[20]),
    .c(cout_21[19]),
    .cout(cout_21[20]),
    .sum(sum_21[20]));
  AL_FADD comp21_21 (
    .a(i21[21]),
    .b(sum_20[21]),
    .c(cout_21[20]),
    .cout(cout_21[21]),
    .sum(sum_21[21]));
  AL_FADD comp21_22 (
    .a(i21[22]),
    .b(sum_20[22]),
    .c(cout_21[21]),
    .cout(cout_21[22]),
    .sum(sum_21[22]));
  AL_FADD comp21_23 (
    .a(i21[23]),
    .b(sum_20[23]),
    .c(cout_21[22]),
    .cout(cout_21[23]),
    .sum(sum_21[23]));
  AL_FADD comp21_24 (
    .a(i21[24]),
    .b(sum_20[24]),
    .c(cout_21[23]),
    .cout(cout_21[24]),
    .sum(sum_21[24]));
  AL_FADD comp21_25 (
    .a(i21[25]),
    .b(sum_20[25]),
    .c(cout_21[24]),
    .cout(cout_21[25]),
    .sum(sum_21[25]));
  AL_FADD comp21_26 (
    .a(i21[26]),
    .b(sum_20[26]),
    .c(cout_21[25]),
    .cout(cout_21[26]),
    .sum(sum_21[26]));
  AL_FADD comp21_27 (
    .a(i21[27]),
    .b(sum_20[27]),
    .c(cout_21[26]),
    .cout(cout_21[27]),
    .sum(sum_21[27]));
  AL_FADD comp21_28 (
    .a(i21[28]),
    .b(sum_20[28]),
    .c(cout_21[27]),
    .cout(cout_21[28]),
    .sum(sum_21[28]));
  AL_FADD comp21_29 (
    .a(i21[29]),
    .b(sum_20[29]),
    .c(cout_21[28]),
    .cout(cout_21[29]),
    .sum(sum_21[29]));
  AL_FADD comp21_3 (
    .a(i21[3]),
    .b(sum_20[3]),
    .c(cout_21[2]),
    .cout(cout_21[3]),
    .sum(sum_21[3]));
  AL_FADD comp21_30 (
    .a(i21[30]),
    .b(sum_20[30]),
    .c(cout_21[29]),
    .cout(cout_21[30]),
    .sum(sum_21[30]));
  AL_FADD comp21_31 (
    .a(i21[31]),
    .b(sum_20[31]),
    .c(cout_21[30]),
    .cout(cout_21[31]),
    .sum(sum_21[31]));
  AL_FADD comp21_32 (
    .a(i21[32]),
    .b(sum_20[32]),
    .c(cout_21[31]),
    .cout(cout_21[32]),
    .sum(sum_21[32]));
  AL_FADD comp21_33 (
    .a(i21[33]),
    .b(sum_20[33]),
    .c(cout_21[32]),
    .cout(cout_21[33]),
    .sum(sum_21[33]));
  AL_FADD comp21_34 (
    .a(i21[34]),
    .b(sum_20[34]),
    .c(cout_21[33]),
    .cout(cout_21[34]),
    .sum(sum_21[34]));
  AL_FADD comp21_35 (
    .a(i21[35]),
    .b(sum_20[35]),
    .c(cout_21[34]),
    .cout(cout_21[35]),
    .sum(sum_21[35]));
  AL_FADD comp21_36 (
    .a(i21[36]),
    .b(sum_20[36]),
    .c(cout_21[35]),
    .cout(cout_21[36]),
    .sum(sum_21[36]));
  AL_FADD comp21_37 (
    .a(i21[37]),
    .b(sum_20[37]),
    .c(cout_21[36]),
    .cout(cout_21[37]),
    .sum(sum_21[37]));
  AL_FADD comp21_38 (
    .a(i21[38]),
    .b(sum_20[38]),
    .c(cout_21[37]),
    .cout(cout_21[38]),
    .sum(sum_21[38]));
  AL_FADD comp21_39 (
    .a(i21[39]),
    .b(sum_20[39]),
    .c(cout_21[38]),
    .cout(cout_21[39]),
    .sum(sum_21[39]));
  AL_FADD comp21_4 (
    .a(i21[4]),
    .b(sum_20[4]),
    .c(cout_21[3]),
    .cout(cout_21[4]),
    .sum(sum_21[4]));
  AL_FADD comp21_40 (
    .a(i21[40]),
    .b(sum_20[40]),
    .c(cout_21[39]),
    .cout(cout_21[40]),
    .sum(sum_21[40]));
  AL_FADD comp21_41 (
    .a(1'b0),
    .b(sum_20[41]),
    .c(cout_21[40]),
    .cout(cout_21[41]),
    .sum(sum_21[41]));
  AL_FADD comp21_42 (
    .a(1'b0),
    .b(sum_20[42]),
    .c(cout_21[41]),
    .cout(cout_21[42]),
    .sum(sum_21[42]));
  AL_FADD comp21_43 (
    .a(1'b0),
    .b(sum_20[43]),
    .c(cout_21[42]),
    .cout(cout_21[43]),
    .sum(sum_21[43]));
  AL_FADD comp21_44 (
    .a(1'b0),
    .b(sum_20[44]),
    .c(cout_21[43]),
    .cout(cout_21[44]),
    .sum(sum_21[44]));
  AL_FADD comp21_45 (
    .a(1'b0),
    .b(sum_20[45]),
    .c(cout_21[44]),
    .cout(cout_21[45]),
    .sum(sum_21[45]));
  AL_FADD comp21_46 (
    .a(1'b0),
    .b(sum_20[46]),
    .c(cout_21[45]),
    .cout(cout_21[46]),
    .sum(sum_21[46]));
  AL_FADD comp21_47 (
    .a(1'b0),
    .b(sum_20[47]),
    .c(cout_21[46]),
    .cout(cout_21[47]),
    .sum(sum_21[47]));
  AL_FADD comp21_48 (
    .a(1'b0),
    .b(sum_20[48]),
    .c(cout_21[47]),
    .cout(cout_21[48]),
    .sum(sum_21[48]));
  AL_FADD comp21_49 (
    .a(1'b0),
    .b(sum_20[49]),
    .c(cout_21[48]),
    .cout(cout_21[49]),
    .sum(sum_21[49]));
  AL_FADD comp21_5 (
    .a(i21[5]),
    .b(sum_20[5]),
    .c(cout_21[4]),
    .cout(cout_21[5]),
    .sum(sum_21[5]));
  AL_FADD comp21_50 (
    .a(1'b0),
    .b(sum_20[50]),
    .c(cout_21[49]),
    .cout(cout_21[50]),
    .sum(sum_21[50]));
  AL_FADD comp21_51 (
    .a(1'b0),
    .b(sum_20[51]),
    .c(cout_21[50]),
    .cout(cout_21[51]),
    .sum(sum_21[51]));
  AL_FADD comp21_52 (
    .a(1'b0),
    .b(sum_20[52]),
    .c(cout_21[51]),
    .cout(cout_21[52]),
    .sum(sum_21[52]));
  AL_FADD comp21_53 (
    .a(1'b0),
    .b(sum_20[53]),
    .c(cout_21[52]),
    .cout(cout_21[53]),
    .sum(sum_21[53]));
  AL_FADD comp21_54 (
    .a(1'b0),
    .b(sum_20[54]),
    .c(cout_21[53]),
    .cout(cout_21[54]),
    .sum(sum_21[54]));
  AL_FADD comp21_55 (
    .a(1'b0),
    .b(sum_20[55]),
    .c(cout_21[54]),
    .cout(cout_21[55]),
    .sum(sum_21[55]));
  AL_FADD comp21_56 (
    .a(1'b0),
    .b(sum_20[56]),
    .c(cout_21[55]),
    .cout(cout_21[56]),
    .sum(sum_21[56]));
  AL_FADD comp21_57 (
    .a(1'b0),
    .b(sum_20[57]),
    .c(cout_21[56]),
    .cout(cout_21[57]),
    .sum(sum_21[57]));
  AL_FADD comp21_58 (
    .a(1'b0),
    .b(sum_20[58]),
    .c(cout_21[57]),
    .cout(cout_21[58]),
    .sum(sum_21[58]));
  AL_FADD comp21_59 (
    .a(1'b0),
    .b(sum_20[59]),
    .c(cout_21[58]),
    .cout(cout_21[59]),
    .sum(sum_21[59]));
  AL_FADD comp21_6 (
    .a(i21[6]),
    .b(sum_20[6]),
    .c(cout_21[5]),
    .cout(cout_21[6]),
    .sum(sum_21[6]));
  AL_FADD comp21_60 (
    .a(1'b0),
    .b(sum_20[60]),
    .c(cout_21[59]),
    .cout(cout_21[60]),
    .sum(sum_21[60]));
  AL_FADD comp21_61 (
    .a(1'b0),
    .b(sum_20[61]),
    .c(cout_21[60]),
    .cout(cout_21[61]),
    .sum(sum_21[61]));
  AL_FADD comp21_62 (
    .a(1'b0),
    .b(sum_20[62]),
    .c(cout_21[61]),
    .cout(cout_21[62]),
    .sum(sum_21[62]));
  AL_FADD comp21_63 (
    .a(1'b0),
    .b(sum_20[63]),
    .c(cout_21[62]),
    .cout(cout_21[63]),
    .sum(sum_21[63]));
  AL_FADD comp21_7 (
    .a(i21[7]),
    .b(sum_20[7]),
    .c(cout_21[6]),
    .cout(cout_21[7]),
    .sum(sum_21[7]));
  AL_FADD comp21_8 (
    .a(i21[8]),
    .b(sum_20[8]),
    .c(cout_21[7]),
    .cout(cout_21[8]),
    .sum(sum_21[8]));
  AL_FADD comp21_9 (
    .a(i21[9]),
    .b(sum_20[9]),
    .c(cout_21[8]),
    .cout(cout_21[9]),
    .sum(sum_21[9]));
  AL_FADD comp22_0 (
    .a(i22[0]),
    .b(sum_21[0]),
    .c(1'b0),
    .cout(cout_22[0]),
    .sum(sum_22[0]));
  AL_FADD comp22_1 (
    .a(i22[1]),
    .b(sum_21[1]),
    .c(cout_22[0]),
    .cout(cout_22[1]),
    .sum(sum_22[1]));
  AL_FADD comp22_10 (
    .a(i22[10]),
    .b(sum_21[10]),
    .c(cout_22[9]),
    .cout(cout_22[10]),
    .sum(sum_22[10]));
  AL_FADD comp22_11 (
    .a(i22[11]),
    .b(sum_21[11]),
    .c(cout_22[10]),
    .cout(cout_22[11]),
    .sum(sum_22[11]));
  AL_FADD comp22_12 (
    .a(i22[12]),
    .b(sum_21[12]),
    .c(cout_22[11]),
    .cout(cout_22[12]),
    .sum(sum_22[12]));
  AL_FADD comp22_13 (
    .a(i22[13]),
    .b(sum_21[13]),
    .c(cout_22[12]),
    .cout(cout_22[13]),
    .sum(sum_22[13]));
  AL_FADD comp22_14 (
    .a(i22[14]),
    .b(sum_21[14]),
    .c(cout_22[13]),
    .cout(cout_22[14]),
    .sum(sum_22[14]));
  AL_FADD comp22_15 (
    .a(i22[15]),
    .b(sum_21[15]),
    .c(cout_22[14]),
    .cout(cout_22[15]),
    .sum(sum_22[15]));
  AL_FADD comp22_16 (
    .a(i22[16]),
    .b(sum_21[16]),
    .c(cout_22[15]),
    .cout(cout_22[16]),
    .sum(sum_22[16]));
  AL_FADD comp22_17 (
    .a(i22[17]),
    .b(sum_21[17]),
    .c(cout_22[16]),
    .cout(cout_22[17]),
    .sum(sum_22[17]));
  AL_FADD comp22_18 (
    .a(i22[18]),
    .b(sum_21[18]),
    .c(cout_22[17]),
    .cout(cout_22[18]),
    .sum(sum_22[18]));
  AL_FADD comp22_19 (
    .a(i22[19]),
    .b(sum_21[19]),
    .c(cout_22[18]),
    .cout(cout_22[19]),
    .sum(sum_22[19]));
  AL_FADD comp22_2 (
    .a(i22[2]),
    .b(sum_21[2]),
    .c(cout_22[1]),
    .cout(cout_22[2]),
    .sum(sum_22[2]));
  AL_FADD comp22_20 (
    .a(i22[20]),
    .b(sum_21[20]),
    .c(cout_22[19]),
    .cout(cout_22[20]),
    .sum(sum_22[20]));
  AL_FADD comp22_21 (
    .a(i22[21]),
    .b(sum_21[21]),
    .c(cout_22[20]),
    .cout(cout_22[21]),
    .sum(sum_22[21]));
  AL_FADD comp22_22 (
    .a(i22[22]),
    .b(sum_21[22]),
    .c(cout_22[21]),
    .cout(cout_22[22]),
    .sum(sum_22[22]));
  AL_FADD comp22_23 (
    .a(i22[23]),
    .b(sum_21[23]),
    .c(cout_22[22]),
    .cout(cout_22[23]),
    .sum(sum_22[23]));
  AL_FADD comp22_24 (
    .a(i22[24]),
    .b(sum_21[24]),
    .c(cout_22[23]),
    .cout(cout_22[24]),
    .sum(sum_22[24]));
  AL_FADD comp22_25 (
    .a(i22[25]),
    .b(sum_21[25]),
    .c(cout_22[24]),
    .cout(cout_22[25]),
    .sum(sum_22[25]));
  AL_FADD comp22_26 (
    .a(i22[26]),
    .b(sum_21[26]),
    .c(cout_22[25]),
    .cout(cout_22[26]),
    .sum(sum_22[26]));
  AL_FADD comp22_27 (
    .a(i22[27]),
    .b(sum_21[27]),
    .c(cout_22[26]),
    .cout(cout_22[27]),
    .sum(sum_22[27]));
  AL_FADD comp22_28 (
    .a(i22[28]),
    .b(sum_21[28]),
    .c(cout_22[27]),
    .cout(cout_22[28]),
    .sum(sum_22[28]));
  AL_FADD comp22_29 (
    .a(i22[29]),
    .b(sum_21[29]),
    .c(cout_22[28]),
    .cout(cout_22[29]),
    .sum(sum_22[29]));
  AL_FADD comp22_3 (
    .a(i22[3]),
    .b(sum_21[3]),
    .c(cout_22[2]),
    .cout(cout_22[3]),
    .sum(sum_22[3]));
  AL_FADD comp22_30 (
    .a(i22[30]),
    .b(sum_21[30]),
    .c(cout_22[29]),
    .cout(cout_22[30]),
    .sum(sum_22[30]));
  AL_FADD comp22_31 (
    .a(i22[31]),
    .b(sum_21[31]),
    .c(cout_22[30]),
    .cout(cout_22[31]),
    .sum(sum_22[31]));
  AL_FADD comp22_32 (
    .a(i22[32]),
    .b(sum_21[32]),
    .c(cout_22[31]),
    .cout(cout_22[32]),
    .sum(sum_22[32]));
  AL_FADD comp22_33 (
    .a(i22[33]),
    .b(sum_21[33]),
    .c(cout_22[32]),
    .cout(cout_22[33]),
    .sum(sum_22[33]));
  AL_FADD comp22_34 (
    .a(i22[34]),
    .b(sum_21[34]),
    .c(cout_22[33]),
    .cout(cout_22[34]),
    .sum(sum_22[34]));
  AL_FADD comp22_35 (
    .a(i22[35]),
    .b(sum_21[35]),
    .c(cout_22[34]),
    .cout(cout_22[35]),
    .sum(sum_22[35]));
  AL_FADD comp22_36 (
    .a(i22[36]),
    .b(sum_21[36]),
    .c(cout_22[35]),
    .cout(cout_22[36]),
    .sum(sum_22[36]));
  AL_FADD comp22_37 (
    .a(i22[37]),
    .b(sum_21[37]),
    .c(cout_22[36]),
    .cout(cout_22[37]),
    .sum(sum_22[37]));
  AL_FADD comp22_38 (
    .a(i22[38]),
    .b(sum_21[38]),
    .c(cout_22[37]),
    .cout(cout_22[38]),
    .sum(sum_22[38]));
  AL_FADD comp22_39 (
    .a(i22[39]),
    .b(sum_21[39]),
    .c(cout_22[38]),
    .cout(cout_22[39]),
    .sum(sum_22[39]));
  AL_FADD comp22_4 (
    .a(i22[4]),
    .b(sum_21[4]),
    .c(cout_22[3]),
    .cout(cout_22[4]),
    .sum(sum_22[4]));
  AL_FADD comp22_40 (
    .a(1'b0),
    .b(sum_21[40]),
    .c(cout_22[39]),
    .cout(cout_22[40]),
    .sum(sum_22[40]));
  AL_FADD comp22_41 (
    .a(1'b0),
    .b(sum_21[41]),
    .c(cout_22[40]),
    .cout(cout_22[41]),
    .sum(sum_22[41]));
  AL_FADD comp22_42 (
    .a(1'b0),
    .b(sum_21[42]),
    .c(cout_22[41]),
    .cout(cout_22[42]),
    .sum(sum_22[42]));
  AL_FADD comp22_43 (
    .a(1'b0),
    .b(sum_21[43]),
    .c(cout_22[42]),
    .cout(cout_22[43]),
    .sum(sum_22[43]));
  AL_FADD comp22_44 (
    .a(1'b0),
    .b(sum_21[44]),
    .c(cout_22[43]),
    .cout(cout_22[44]),
    .sum(sum_22[44]));
  AL_FADD comp22_45 (
    .a(1'b0),
    .b(sum_21[45]),
    .c(cout_22[44]),
    .cout(cout_22[45]),
    .sum(sum_22[45]));
  AL_FADD comp22_46 (
    .a(1'b0),
    .b(sum_21[46]),
    .c(cout_22[45]),
    .cout(cout_22[46]),
    .sum(sum_22[46]));
  AL_FADD comp22_47 (
    .a(1'b0),
    .b(sum_21[47]),
    .c(cout_22[46]),
    .cout(cout_22[47]),
    .sum(sum_22[47]));
  AL_FADD comp22_48 (
    .a(1'b0),
    .b(sum_21[48]),
    .c(cout_22[47]),
    .cout(cout_22[48]),
    .sum(sum_22[48]));
  AL_FADD comp22_49 (
    .a(1'b0),
    .b(sum_21[49]),
    .c(cout_22[48]),
    .cout(cout_22[49]),
    .sum(sum_22[49]));
  AL_FADD comp22_5 (
    .a(i22[5]),
    .b(sum_21[5]),
    .c(cout_22[4]),
    .cout(cout_22[5]),
    .sum(sum_22[5]));
  AL_FADD comp22_50 (
    .a(1'b0),
    .b(sum_21[50]),
    .c(cout_22[49]),
    .cout(cout_22[50]),
    .sum(sum_22[50]));
  AL_FADD comp22_51 (
    .a(1'b0),
    .b(sum_21[51]),
    .c(cout_22[50]),
    .cout(cout_22[51]),
    .sum(sum_22[51]));
  AL_FADD comp22_52 (
    .a(1'b0),
    .b(sum_21[52]),
    .c(cout_22[51]),
    .cout(cout_22[52]),
    .sum(sum_22[52]));
  AL_FADD comp22_53 (
    .a(1'b0),
    .b(sum_21[53]),
    .c(cout_22[52]),
    .cout(cout_22[53]),
    .sum(sum_22[53]));
  AL_FADD comp22_54 (
    .a(1'b0),
    .b(sum_21[54]),
    .c(cout_22[53]),
    .cout(cout_22[54]),
    .sum(sum_22[54]));
  AL_FADD comp22_55 (
    .a(1'b0),
    .b(sum_21[55]),
    .c(cout_22[54]),
    .cout(cout_22[55]),
    .sum(sum_22[55]));
  AL_FADD comp22_56 (
    .a(1'b0),
    .b(sum_21[56]),
    .c(cout_22[55]),
    .cout(cout_22[56]),
    .sum(sum_22[56]));
  AL_FADD comp22_57 (
    .a(1'b0),
    .b(sum_21[57]),
    .c(cout_22[56]),
    .cout(cout_22[57]),
    .sum(sum_22[57]));
  AL_FADD comp22_58 (
    .a(1'b0),
    .b(sum_21[58]),
    .c(cout_22[57]),
    .cout(cout_22[58]),
    .sum(sum_22[58]));
  AL_FADD comp22_59 (
    .a(1'b0),
    .b(sum_21[59]),
    .c(cout_22[58]),
    .cout(cout_22[59]),
    .sum(sum_22[59]));
  AL_FADD comp22_6 (
    .a(i22[6]),
    .b(sum_21[6]),
    .c(cout_22[5]),
    .cout(cout_22[6]),
    .sum(sum_22[6]));
  AL_FADD comp22_60 (
    .a(1'b0),
    .b(sum_21[60]),
    .c(cout_22[59]),
    .cout(cout_22[60]),
    .sum(sum_22[60]));
  AL_FADD comp22_61 (
    .a(1'b0),
    .b(sum_21[61]),
    .c(cout_22[60]),
    .cout(cout_22[61]),
    .sum(sum_22[61]));
  AL_FADD comp22_62 (
    .a(1'b0),
    .b(sum_21[62]),
    .c(cout_22[61]),
    .cout(cout_22[62]),
    .sum(sum_22[62]));
  AL_FADD comp22_63 (
    .a(1'b0),
    .b(sum_21[63]),
    .c(cout_22[62]),
    .cout(cout_22[63]),
    .sum(sum_22[63]));
  AL_FADD comp22_7 (
    .a(i22[7]),
    .b(sum_21[7]),
    .c(cout_22[6]),
    .cout(cout_22[7]),
    .sum(sum_22[7]));
  AL_FADD comp22_8 (
    .a(i22[8]),
    .b(sum_21[8]),
    .c(cout_22[7]),
    .cout(cout_22[8]),
    .sum(sum_22[8]));
  AL_FADD comp22_9 (
    .a(i22[9]),
    .b(sum_21[9]),
    .c(cout_22[8]),
    .cout(cout_22[9]),
    .sum(sum_22[9]));
  AL_FADD comp23_0 (
    .a(i23[0]),
    .b(sum_22[0]),
    .c(1'b0),
    .cout(cout_23[0]),
    .sum(sum_23[0]));
  AL_FADD comp23_1 (
    .a(i23[1]),
    .b(sum_22[1]),
    .c(cout_23[0]),
    .cout(cout_23[1]),
    .sum(sum_23[1]));
  AL_FADD comp23_10 (
    .a(i23[10]),
    .b(sum_22[10]),
    .c(cout_23[9]),
    .cout(cout_23[10]),
    .sum(sum_23[10]));
  AL_FADD comp23_11 (
    .a(i23[11]),
    .b(sum_22[11]),
    .c(cout_23[10]),
    .cout(cout_23[11]),
    .sum(sum_23[11]));
  AL_FADD comp23_12 (
    .a(i23[12]),
    .b(sum_22[12]),
    .c(cout_23[11]),
    .cout(cout_23[12]),
    .sum(sum_23[12]));
  AL_FADD comp23_13 (
    .a(i23[13]),
    .b(sum_22[13]),
    .c(cout_23[12]),
    .cout(cout_23[13]),
    .sum(sum_23[13]));
  AL_FADD comp23_14 (
    .a(i23[14]),
    .b(sum_22[14]),
    .c(cout_23[13]),
    .cout(cout_23[14]),
    .sum(sum_23[14]));
  AL_FADD comp23_15 (
    .a(i23[15]),
    .b(sum_22[15]),
    .c(cout_23[14]),
    .cout(cout_23[15]),
    .sum(sum_23[15]));
  AL_FADD comp23_16 (
    .a(i23[16]),
    .b(sum_22[16]),
    .c(cout_23[15]),
    .cout(cout_23[16]),
    .sum(sum_23[16]));
  AL_FADD comp23_17 (
    .a(i23[17]),
    .b(sum_22[17]),
    .c(cout_23[16]),
    .cout(cout_23[17]),
    .sum(sum_23[17]));
  AL_FADD comp23_18 (
    .a(i23[18]),
    .b(sum_22[18]),
    .c(cout_23[17]),
    .cout(cout_23[18]),
    .sum(sum_23[18]));
  AL_FADD comp23_19 (
    .a(i23[19]),
    .b(sum_22[19]),
    .c(cout_23[18]),
    .cout(cout_23[19]),
    .sum(sum_23[19]));
  AL_FADD comp23_2 (
    .a(i23[2]),
    .b(sum_22[2]),
    .c(cout_23[1]),
    .cout(cout_23[2]),
    .sum(sum_23[2]));
  AL_FADD comp23_20 (
    .a(i23[20]),
    .b(sum_22[20]),
    .c(cout_23[19]),
    .cout(cout_23[20]),
    .sum(sum_23[20]));
  AL_FADD comp23_21 (
    .a(i23[21]),
    .b(sum_22[21]),
    .c(cout_23[20]),
    .cout(cout_23[21]),
    .sum(sum_23[21]));
  AL_FADD comp23_22 (
    .a(i23[22]),
    .b(sum_22[22]),
    .c(cout_23[21]),
    .cout(cout_23[22]),
    .sum(sum_23[22]));
  AL_FADD comp23_23 (
    .a(i23[23]),
    .b(sum_22[23]),
    .c(cout_23[22]),
    .cout(cout_23[23]),
    .sum(sum_23[23]));
  AL_FADD comp23_24 (
    .a(i23[24]),
    .b(sum_22[24]),
    .c(cout_23[23]),
    .cout(cout_23[24]),
    .sum(sum_23[24]));
  AL_FADD comp23_25 (
    .a(i23[25]),
    .b(sum_22[25]),
    .c(cout_23[24]),
    .cout(cout_23[25]),
    .sum(sum_23[25]));
  AL_FADD comp23_26 (
    .a(i23[26]),
    .b(sum_22[26]),
    .c(cout_23[25]),
    .cout(cout_23[26]),
    .sum(sum_23[26]));
  AL_FADD comp23_27 (
    .a(i23[27]),
    .b(sum_22[27]),
    .c(cout_23[26]),
    .cout(cout_23[27]),
    .sum(sum_23[27]));
  AL_FADD comp23_28 (
    .a(i23[28]),
    .b(sum_22[28]),
    .c(cout_23[27]),
    .cout(cout_23[28]),
    .sum(sum_23[28]));
  AL_FADD comp23_29 (
    .a(i23[29]),
    .b(sum_22[29]),
    .c(cout_23[28]),
    .cout(cout_23[29]),
    .sum(sum_23[29]));
  AL_FADD comp23_3 (
    .a(i23[3]),
    .b(sum_22[3]),
    .c(cout_23[2]),
    .cout(cout_23[3]),
    .sum(sum_23[3]));
  AL_FADD comp23_30 (
    .a(i23[30]),
    .b(sum_22[30]),
    .c(cout_23[29]),
    .cout(cout_23[30]),
    .sum(sum_23[30]));
  AL_FADD comp23_31 (
    .a(i23[31]),
    .b(sum_22[31]),
    .c(cout_23[30]),
    .cout(cout_23[31]),
    .sum(sum_23[31]));
  AL_FADD comp23_32 (
    .a(i23[32]),
    .b(sum_22[32]),
    .c(cout_23[31]),
    .cout(cout_23[32]),
    .sum(sum_23[32]));
  AL_FADD comp23_33 (
    .a(i23[33]),
    .b(sum_22[33]),
    .c(cout_23[32]),
    .cout(cout_23[33]),
    .sum(sum_23[33]));
  AL_FADD comp23_34 (
    .a(i23[34]),
    .b(sum_22[34]),
    .c(cout_23[33]),
    .cout(cout_23[34]),
    .sum(sum_23[34]));
  AL_FADD comp23_35 (
    .a(i23[35]),
    .b(sum_22[35]),
    .c(cout_23[34]),
    .cout(cout_23[35]),
    .sum(sum_23[35]));
  AL_FADD comp23_36 (
    .a(i23[36]),
    .b(sum_22[36]),
    .c(cout_23[35]),
    .cout(cout_23[36]),
    .sum(sum_23[36]));
  AL_FADD comp23_37 (
    .a(i23[37]),
    .b(sum_22[37]),
    .c(cout_23[36]),
    .cout(cout_23[37]),
    .sum(sum_23[37]));
  AL_FADD comp23_38 (
    .a(i23[38]),
    .b(sum_22[38]),
    .c(cout_23[37]),
    .cout(cout_23[38]),
    .sum(sum_23[38]));
  AL_FADD comp23_39 (
    .a(1'b0),
    .b(sum_22[39]),
    .c(cout_23[38]),
    .cout(cout_23[39]),
    .sum(sum_23[39]));
  AL_FADD comp23_4 (
    .a(i23[4]),
    .b(sum_22[4]),
    .c(cout_23[3]),
    .cout(cout_23[4]),
    .sum(sum_23[4]));
  AL_FADD comp23_40 (
    .a(1'b0),
    .b(sum_22[40]),
    .c(cout_23[39]),
    .cout(cout_23[40]),
    .sum(sum_23[40]));
  AL_FADD comp23_41 (
    .a(1'b0),
    .b(sum_22[41]),
    .c(cout_23[40]),
    .cout(cout_23[41]),
    .sum(sum_23[41]));
  AL_FADD comp23_42 (
    .a(1'b0),
    .b(sum_22[42]),
    .c(cout_23[41]),
    .cout(cout_23[42]),
    .sum(sum_23[42]));
  AL_FADD comp23_43 (
    .a(1'b0),
    .b(sum_22[43]),
    .c(cout_23[42]),
    .cout(cout_23[43]),
    .sum(sum_23[43]));
  AL_FADD comp23_44 (
    .a(1'b0),
    .b(sum_22[44]),
    .c(cout_23[43]),
    .cout(cout_23[44]),
    .sum(sum_23[44]));
  AL_FADD comp23_45 (
    .a(1'b0),
    .b(sum_22[45]),
    .c(cout_23[44]),
    .cout(cout_23[45]),
    .sum(sum_23[45]));
  AL_FADD comp23_46 (
    .a(1'b0),
    .b(sum_22[46]),
    .c(cout_23[45]),
    .cout(cout_23[46]),
    .sum(sum_23[46]));
  AL_FADD comp23_47 (
    .a(1'b0),
    .b(sum_22[47]),
    .c(cout_23[46]),
    .cout(cout_23[47]),
    .sum(sum_23[47]));
  AL_FADD comp23_48 (
    .a(1'b0),
    .b(sum_22[48]),
    .c(cout_23[47]),
    .cout(cout_23[48]),
    .sum(sum_23[48]));
  AL_FADD comp23_49 (
    .a(1'b0),
    .b(sum_22[49]),
    .c(cout_23[48]),
    .cout(cout_23[49]),
    .sum(sum_23[49]));
  AL_FADD comp23_5 (
    .a(i23[5]),
    .b(sum_22[5]),
    .c(cout_23[4]),
    .cout(cout_23[5]),
    .sum(sum_23[5]));
  AL_FADD comp23_50 (
    .a(1'b0),
    .b(sum_22[50]),
    .c(cout_23[49]),
    .cout(cout_23[50]),
    .sum(sum_23[50]));
  AL_FADD comp23_51 (
    .a(1'b0),
    .b(sum_22[51]),
    .c(cout_23[50]),
    .cout(cout_23[51]),
    .sum(sum_23[51]));
  AL_FADD comp23_52 (
    .a(1'b0),
    .b(sum_22[52]),
    .c(cout_23[51]),
    .cout(cout_23[52]),
    .sum(sum_23[52]));
  AL_FADD comp23_53 (
    .a(1'b0),
    .b(sum_22[53]),
    .c(cout_23[52]),
    .cout(cout_23[53]),
    .sum(sum_23[53]));
  AL_FADD comp23_54 (
    .a(1'b0),
    .b(sum_22[54]),
    .c(cout_23[53]),
    .cout(cout_23[54]),
    .sum(sum_23[54]));
  AL_FADD comp23_55 (
    .a(1'b0),
    .b(sum_22[55]),
    .c(cout_23[54]),
    .cout(cout_23[55]),
    .sum(sum_23[55]));
  AL_FADD comp23_56 (
    .a(1'b0),
    .b(sum_22[56]),
    .c(cout_23[55]),
    .cout(cout_23[56]),
    .sum(sum_23[56]));
  AL_FADD comp23_57 (
    .a(1'b0),
    .b(sum_22[57]),
    .c(cout_23[56]),
    .cout(cout_23[57]),
    .sum(sum_23[57]));
  AL_FADD comp23_58 (
    .a(1'b0),
    .b(sum_22[58]),
    .c(cout_23[57]),
    .cout(cout_23[58]),
    .sum(sum_23[58]));
  AL_FADD comp23_59 (
    .a(1'b0),
    .b(sum_22[59]),
    .c(cout_23[58]),
    .cout(cout_23[59]),
    .sum(sum_23[59]));
  AL_FADD comp23_6 (
    .a(i23[6]),
    .b(sum_22[6]),
    .c(cout_23[5]),
    .cout(cout_23[6]),
    .sum(sum_23[6]));
  AL_FADD comp23_60 (
    .a(1'b0),
    .b(sum_22[60]),
    .c(cout_23[59]),
    .cout(cout_23[60]),
    .sum(sum_23[60]));
  AL_FADD comp23_61 (
    .a(1'b0),
    .b(sum_22[61]),
    .c(cout_23[60]),
    .cout(cout_23[61]),
    .sum(sum_23[61]));
  AL_FADD comp23_62 (
    .a(1'b0),
    .b(sum_22[62]),
    .c(cout_23[61]),
    .cout(cout_23[62]),
    .sum(sum_23[62]));
  AL_FADD comp23_63 (
    .a(1'b0),
    .b(sum_22[63]),
    .c(cout_23[62]),
    .cout(cout_23[63]),
    .sum(sum_23[63]));
  AL_FADD comp23_7 (
    .a(i23[7]),
    .b(sum_22[7]),
    .c(cout_23[6]),
    .cout(cout_23[7]),
    .sum(sum_23[7]));
  AL_FADD comp23_8 (
    .a(i23[8]),
    .b(sum_22[8]),
    .c(cout_23[7]),
    .cout(cout_23[8]),
    .sum(sum_23[8]));
  AL_FADD comp23_9 (
    .a(i23[9]),
    .b(sum_22[9]),
    .c(cout_23[8]),
    .cout(cout_23[9]),
    .sum(sum_23[9]));
  AL_FADD comp24_0 (
    .a(i24[0]),
    .b(sum_23[0]),
    .c(1'b0),
    .cout(cout_24[0]),
    .sum(sum_24[0]));
  AL_FADD comp24_1 (
    .a(i24[1]),
    .b(sum_23[1]),
    .c(cout_24[0]),
    .cout(cout_24[1]),
    .sum(sum_24[1]));
  AL_FADD comp24_10 (
    .a(i24[10]),
    .b(sum_23[10]),
    .c(cout_24[9]),
    .cout(cout_24[10]),
    .sum(sum_24[10]));
  AL_FADD comp24_11 (
    .a(i24[11]),
    .b(sum_23[11]),
    .c(cout_24[10]),
    .cout(cout_24[11]),
    .sum(sum_24[11]));
  AL_FADD comp24_12 (
    .a(i24[12]),
    .b(sum_23[12]),
    .c(cout_24[11]),
    .cout(cout_24[12]),
    .sum(sum_24[12]));
  AL_FADD comp24_13 (
    .a(i24[13]),
    .b(sum_23[13]),
    .c(cout_24[12]),
    .cout(cout_24[13]),
    .sum(sum_24[13]));
  AL_FADD comp24_14 (
    .a(i24[14]),
    .b(sum_23[14]),
    .c(cout_24[13]),
    .cout(cout_24[14]),
    .sum(sum_24[14]));
  AL_FADD comp24_15 (
    .a(i24[15]),
    .b(sum_23[15]),
    .c(cout_24[14]),
    .cout(cout_24[15]),
    .sum(sum_24[15]));
  AL_FADD comp24_16 (
    .a(i24[16]),
    .b(sum_23[16]),
    .c(cout_24[15]),
    .cout(cout_24[16]),
    .sum(sum_24[16]));
  AL_FADD comp24_17 (
    .a(i24[17]),
    .b(sum_23[17]),
    .c(cout_24[16]),
    .cout(cout_24[17]),
    .sum(sum_24[17]));
  AL_FADD comp24_18 (
    .a(i24[18]),
    .b(sum_23[18]),
    .c(cout_24[17]),
    .cout(cout_24[18]),
    .sum(sum_24[18]));
  AL_FADD comp24_19 (
    .a(i24[19]),
    .b(sum_23[19]),
    .c(cout_24[18]),
    .cout(cout_24[19]),
    .sum(sum_24[19]));
  AL_FADD comp24_2 (
    .a(i24[2]),
    .b(sum_23[2]),
    .c(cout_24[1]),
    .cout(cout_24[2]),
    .sum(sum_24[2]));
  AL_FADD comp24_20 (
    .a(i24[20]),
    .b(sum_23[20]),
    .c(cout_24[19]),
    .cout(cout_24[20]),
    .sum(sum_24[20]));
  AL_FADD comp24_21 (
    .a(i24[21]),
    .b(sum_23[21]),
    .c(cout_24[20]),
    .cout(cout_24[21]),
    .sum(sum_24[21]));
  AL_FADD comp24_22 (
    .a(i24[22]),
    .b(sum_23[22]),
    .c(cout_24[21]),
    .cout(cout_24[22]),
    .sum(sum_24[22]));
  AL_FADD comp24_23 (
    .a(i24[23]),
    .b(sum_23[23]),
    .c(cout_24[22]),
    .cout(cout_24[23]),
    .sum(sum_24[23]));
  AL_FADD comp24_24 (
    .a(i24[24]),
    .b(sum_23[24]),
    .c(cout_24[23]),
    .cout(cout_24[24]),
    .sum(sum_24[24]));
  AL_FADD comp24_25 (
    .a(i24[25]),
    .b(sum_23[25]),
    .c(cout_24[24]),
    .cout(cout_24[25]),
    .sum(sum_24[25]));
  AL_FADD comp24_26 (
    .a(i24[26]),
    .b(sum_23[26]),
    .c(cout_24[25]),
    .cout(cout_24[26]),
    .sum(sum_24[26]));
  AL_FADD comp24_27 (
    .a(i24[27]),
    .b(sum_23[27]),
    .c(cout_24[26]),
    .cout(cout_24[27]),
    .sum(sum_24[27]));
  AL_FADD comp24_28 (
    .a(i24[28]),
    .b(sum_23[28]),
    .c(cout_24[27]),
    .cout(cout_24[28]),
    .sum(sum_24[28]));
  AL_FADD comp24_29 (
    .a(i24[29]),
    .b(sum_23[29]),
    .c(cout_24[28]),
    .cout(cout_24[29]),
    .sum(sum_24[29]));
  AL_FADD comp24_3 (
    .a(i24[3]),
    .b(sum_23[3]),
    .c(cout_24[2]),
    .cout(cout_24[3]),
    .sum(sum_24[3]));
  AL_FADD comp24_30 (
    .a(i24[30]),
    .b(sum_23[30]),
    .c(cout_24[29]),
    .cout(cout_24[30]),
    .sum(sum_24[30]));
  AL_FADD comp24_31 (
    .a(i24[31]),
    .b(sum_23[31]),
    .c(cout_24[30]),
    .cout(cout_24[31]),
    .sum(sum_24[31]));
  AL_FADD comp24_32 (
    .a(i24[32]),
    .b(sum_23[32]),
    .c(cout_24[31]),
    .cout(cout_24[32]),
    .sum(sum_24[32]));
  AL_FADD comp24_33 (
    .a(i24[33]),
    .b(sum_23[33]),
    .c(cout_24[32]),
    .cout(cout_24[33]),
    .sum(sum_24[33]));
  AL_FADD comp24_34 (
    .a(i24[34]),
    .b(sum_23[34]),
    .c(cout_24[33]),
    .cout(cout_24[34]),
    .sum(sum_24[34]));
  AL_FADD comp24_35 (
    .a(i24[35]),
    .b(sum_23[35]),
    .c(cout_24[34]),
    .cout(cout_24[35]),
    .sum(sum_24[35]));
  AL_FADD comp24_36 (
    .a(i24[36]),
    .b(sum_23[36]),
    .c(cout_24[35]),
    .cout(cout_24[36]),
    .sum(sum_24[36]));
  AL_FADD comp24_37 (
    .a(i24[37]),
    .b(sum_23[37]),
    .c(cout_24[36]),
    .cout(cout_24[37]),
    .sum(sum_24[37]));
  AL_FADD comp24_38 (
    .a(1'b0),
    .b(sum_23[38]),
    .c(cout_24[37]),
    .cout(cout_24[38]),
    .sum(sum_24[38]));
  AL_FADD comp24_39 (
    .a(1'b0),
    .b(sum_23[39]),
    .c(cout_24[38]),
    .cout(cout_24[39]),
    .sum(sum_24[39]));
  AL_FADD comp24_4 (
    .a(i24[4]),
    .b(sum_23[4]),
    .c(cout_24[3]),
    .cout(cout_24[4]),
    .sum(sum_24[4]));
  AL_FADD comp24_40 (
    .a(1'b0),
    .b(sum_23[40]),
    .c(cout_24[39]),
    .cout(cout_24[40]),
    .sum(sum_24[40]));
  AL_FADD comp24_41 (
    .a(1'b0),
    .b(sum_23[41]),
    .c(cout_24[40]),
    .cout(cout_24[41]),
    .sum(sum_24[41]));
  AL_FADD comp24_42 (
    .a(1'b0),
    .b(sum_23[42]),
    .c(cout_24[41]),
    .cout(cout_24[42]),
    .sum(sum_24[42]));
  AL_FADD comp24_43 (
    .a(1'b0),
    .b(sum_23[43]),
    .c(cout_24[42]),
    .cout(cout_24[43]),
    .sum(sum_24[43]));
  AL_FADD comp24_44 (
    .a(1'b0),
    .b(sum_23[44]),
    .c(cout_24[43]),
    .cout(cout_24[44]),
    .sum(sum_24[44]));
  AL_FADD comp24_45 (
    .a(1'b0),
    .b(sum_23[45]),
    .c(cout_24[44]),
    .cout(cout_24[45]),
    .sum(sum_24[45]));
  AL_FADD comp24_46 (
    .a(1'b0),
    .b(sum_23[46]),
    .c(cout_24[45]),
    .cout(cout_24[46]),
    .sum(sum_24[46]));
  AL_FADD comp24_47 (
    .a(1'b0),
    .b(sum_23[47]),
    .c(cout_24[46]),
    .cout(cout_24[47]),
    .sum(sum_24[47]));
  AL_FADD comp24_48 (
    .a(1'b0),
    .b(sum_23[48]),
    .c(cout_24[47]),
    .cout(cout_24[48]),
    .sum(sum_24[48]));
  AL_FADD comp24_49 (
    .a(1'b0),
    .b(sum_23[49]),
    .c(cout_24[48]),
    .cout(cout_24[49]),
    .sum(sum_24[49]));
  AL_FADD comp24_5 (
    .a(i24[5]),
    .b(sum_23[5]),
    .c(cout_24[4]),
    .cout(cout_24[5]),
    .sum(sum_24[5]));
  AL_FADD comp24_50 (
    .a(1'b0),
    .b(sum_23[50]),
    .c(cout_24[49]),
    .cout(cout_24[50]),
    .sum(sum_24[50]));
  AL_FADD comp24_51 (
    .a(1'b0),
    .b(sum_23[51]),
    .c(cout_24[50]),
    .cout(cout_24[51]),
    .sum(sum_24[51]));
  AL_FADD comp24_52 (
    .a(1'b0),
    .b(sum_23[52]),
    .c(cout_24[51]),
    .cout(cout_24[52]),
    .sum(sum_24[52]));
  AL_FADD comp24_53 (
    .a(1'b0),
    .b(sum_23[53]),
    .c(cout_24[52]),
    .cout(cout_24[53]),
    .sum(sum_24[53]));
  AL_FADD comp24_54 (
    .a(1'b0),
    .b(sum_23[54]),
    .c(cout_24[53]),
    .cout(cout_24[54]),
    .sum(sum_24[54]));
  AL_FADD comp24_55 (
    .a(1'b0),
    .b(sum_23[55]),
    .c(cout_24[54]),
    .cout(cout_24[55]),
    .sum(sum_24[55]));
  AL_FADD comp24_56 (
    .a(1'b0),
    .b(sum_23[56]),
    .c(cout_24[55]),
    .cout(cout_24[56]),
    .sum(sum_24[56]));
  AL_FADD comp24_57 (
    .a(1'b0),
    .b(sum_23[57]),
    .c(cout_24[56]),
    .cout(cout_24[57]),
    .sum(sum_24[57]));
  AL_FADD comp24_58 (
    .a(1'b0),
    .b(sum_23[58]),
    .c(cout_24[57]),
    .cout(cout_24[58]),
    .sum(sum_24[58]));
  AL_FADD comp24_59 (
    .a(1'b0),
    .b(sum_23[59]),
    .c(cout_24[58]),
    .cout(cout_24[59]),
    .sum(sum_24[59]));
  AL_FADD comp24_6 (
    .a(i24[6]),
    .b(sum_23[6]),
    .c(cout_24[5]),
    .cout(cout_24[6]),
    .sum(sum_24[6]));
  AL_FADD comp24_60 (
    .a(1'b0),
    .b(sum_23[60]),
    .c(cout_24[59]),
    .cout(cout_24[60]),
    .sum(sum_24[60]));
  AL_FADD comp24_61 (
    .a(1'b0),
    .b(sum_23[61]),
    .c(cout_24[60]),
    .cout(cout_24[61]),
    .sum(sum_24[61]));
  AL_FADD comp24_62 (
    .a(1'b0),
    .b(sum_23[62]),
    .c(cout_24[61]),
    .cout(cout_24[62]),
    .sum(sum_24[62]));
  AL_FADD comp24_63 (
    .a(1'b0),
    .b(sum_23[63]),
    .c(cout_24[62]),
    .cout(cout_24[63]),
    .sum(sum_24[63]));
  AL_FADD comp24_7 (
    .a(i24[7]),
    .b(sum_23[7]),
    .c(cout_24[6]),
    .cout(cout_24[7]),
    .sum(sum_24[7]));
  AL_FADD comp24_8 (
    .a(i24[8]),
    .b(sum_23[8]),
    .c(cout_24[7]),
    .cout(cout_24[8]),
    .sum(sum_24[8]));
  AL_FADD comp24_9 (
    .a(i24[9]),
    .b(sum_23[9]),
    .c(cout_24[8]),
    .cout(cout_24[9]),
    .sum(sum_24[9]));
  AL_FADD comp25_0 (
    .a(i25[0]),
    .b(sum_24[0]),
    .c(1'b0),
    .cout(cout_25[0]),
    .sum(sum_25[0]));
  AL_FADD comp25_1 (
    .a(i25[1]),
    .b(sum_24[1]),
    .c(cout_25[0]),
    .cout(cout_25[1]),
    .sum(sum_25[1]));
  AL_FADD comp25_10 (
    .a(i25[10]),
    .b(sum_24[10]),
    .c(cout_25[9]),
    .cout(cout_25[10]),
    .sum(sum_25[10]));
  AL_FADD comp25_11 (
    .a(i25[11]),
    .b(sum_24[11]),
    .c(cout_25[10]),
    .cout(cout_25[11]),
    .sum(sum_25[11]));
  AL_FADD comp25_12 (
    .a(i25[12]),
    .b(sum_24[12]),
    .c(cout_25[11]),
    .cout(cout_25[12]),
    .sum(sum_25[12]));
  AL_FADD comp25_13 (
    .a(i25[13]),
    .b(sum_24[13]),
    .c(cout_25[12]),
    .cout(cout_25[13]),
    .sum(sum_25[13]));
  AL_FADD comp25_14 (
    .a(i25[14]),
    .b(sum_24[14]),
    .c(cout_25[13]),
    .cout(cout_25[14]),
    .sum(sum_25[14]));
  AL_FADD comp25_15 (
    .a(i25[15]),
    .b(sum_24[15]),
    .c(cout_25[14]),
    .cout(cout_25[15]),
    .sum(sum_25[15]));
  AL_FADD comp25_16 (
    .a(i25[16]),
    .b(sum_24[16]),
    .c(cout_25[15]),
    .cout(cout_25[16]),
    .sum(sum_25[16]));
  AL_FADD comp25_17 (
    .a(i25[17]),
    .b(sum_24[17]),
    .c(cout_25[16]),
    .cout(cout_25[17]),
    .sum(sum_25[17]));
  AL_FADD comp25_18 (
    .a(i25[18]),
    .b(sum_24[18]),
    .c(cout_25[17]),
    .cout(cout_25[18]),
    .sum(sum_25[18]));
  AL_FADD comp25_19 (
    .a(i25[19]),
    .b(sum_24[19]),
    .c(cout_25[18]),
    .cout(cout_25[19]),
    .sum(sum_25[19]));
  AL_FADD comp25_2 (
    .a(i25[2]),
    .b(sum_24[2]),
    .c(cout_25[1]),
    .cout(cout_25[2]),
    .sum(sum_25[2]));
  AL_FADD comp25_20 (
    .a(i25[20]),
    .b(sum_24[20]),
    .c(cout_25[19]),
    .cout(cout_25[20]),
    .sum(sum_25[20]));
  AL_FADD comp25_21 (
    .a(i25[21]),
    .b(sum_24[21]),
    .c(cout_25[20]),
    .cout(cout_25[21]),
    .sum(sum_25[21]));
  AL_FADD comp25_22 (
    .a(i25[22]),
    .b(sum_24[22]),
    .c(cout_25[21]),
    .cout(cout_25[22]),
    .sum(sum_25[22]));
  AL_FADD comp25_23 (
    .a(i25[23]),
    .b(sum_24[23]),
    .c(cout_25[22]),
    .cout(cout_25[23]),
    .sum(sum_25[23]));
  AL_FADD comp25_24 (
    .a(i25[24]),
    .b(sum_24[24]),
    .c(cout_25[23]),
    .cout(cout_25[24]),
    .sum(sum_25[24]));
  AL_FADD comp25_25 (
    .a(i25[25]),
    .b(sum_24[25]),
    .c(cout_25[24]),
    .cout(cout_25[25]),
    .sum(sum_25[25]));
  AL_FADD comp25_26 (
    .a(i25[26]),
    .b(sum_24[26]),
    .c(cout_25[25]),
    .cout(cout_25[26]),
    .sum(sum_25[26]));
  AL_FADD comp25_27 (
    .a(i25[27]),
    .b(sum_24[27]),
    .c(cout_25[26]),
    .cout(cout_25[27]),
    .sum(sum_25[27]));
  AL_FADD comp25_28 (
    .a(i25[28]),
    .b(sum_24[28]),
    .c(cout_25[27]),
    .cout(cout_25[28]),
    .sum(sum_25[28]));
  AL_FADD comp25_29 (
    .a(i25[29]),
    .b(sum_24[29]),
    .c(cout_25[28]),
    .cout(cout_25[29]),
    .sum(sum_25[29]));
  AL_FADD comp25_3 (
    .a(i25[3]),
    .b(sum_24[3]),
    .c(cout_25[2]),
    .cout(cout_25[3]),
    .sum(sum_25[3]));
  AL_FADD comp25_30 (
    .a(i25[30]),
    .b(sum_24[30]),
    .c(cout_25[29]),
    .cout(cout_25[30]),
    .sum(sum_25[30]));
  AL_FADD comp25_31 (
    .a(i25[31]),
    .b(sum_24[31]),
    .c(cout_25[30]),
    .cout(cout_25[31]),
    .sum(sum_25[31]));
  AL_FADD comp25_32 (
    .a(i25[32]),
    .b(sum_24[32]),
    .c(cout_25[31]),
    .cout(cout_25[32]),
    .sum(sum_25[32]));
  AL_FADD comp25_33 (
    .a(i25[33]),
    .b(sum_24[33]),
    .c(cout_25[32]),
    .cout(cout_25[33]),
    .sum(sum_25[33]));
  AL_FADD comp25_34 (
    .a(i25[34]),
    .b(sum_24[34]),
    .c(cout_25[33]),
    .cout(cout_25[34]),
    .sum(sum_25[34]));
  AL_FADD comp25_35 (
    .a(i25[35]),
    .b(sum_24[35]),
    .c(cout_25[34]),
    .cout(cout_25[35]),
    .sum(sum_25[35]));
  AL_FADD comp25_36 (
    .a(i25[36]),
    .b(sum_24[36]),
    .c(cout_25[35]),
    .cout(cout_25[36]),
    .sum(sum_25[36]));
  AL_FADD comp25_37 (
    .a(1'b0),
    .b(sum_24[37]),
    .c(cout_25[36]),
    .cout(cout_25[37]),
    .sum(sum_25[37]));
  AL_FADD comp25_38 (
    .a(1'b0),
    .b(sum_24[38]),
    .c(cout_25[37]),
    .cout(cout_25[38]),
    .sum(sum_25[38]));
  AL_FADD comp25_39 (
    .a(1'b0),
    .b(sum_24[39]),
    .c(cout_25[38]),
    .cout(cout_25[39]),
    .sum(sum_25[39]));
  AL_FADD comp25_4 (
    .a(i25[4]),
    .b(sum_24[4]),
    .c(cout_25[3]),
    .cout(cout_25[4]),
    .sum(sum_25[4]));
  AL_FADD comp25_40 (
    .a(1'b0),
    .b(sum_24[40]),
    .c(cout_25[39]),
    .cout(cout_25[40]),
    .sum(sum_25[40]));
  AL_FADD comp25_41 (
    .a(1'b0),
    .b(sum_24[41]),
    .c(cout_25[40]),
    .cout(cout_25[41]),
    .sum(sum_25[41]));
  AL_FADD comp25_42 (
    .a(1'b0),
    .b(sum_24[42]),
    .c(cout_25[41]),
    .cout(cout_25[42]),
    .sum(sum_25[42]));
  AL_FADD comp25_43 (
    .a(1'b0),
    .b(sum_24[43]),
    .c(cout_25[42]),
    .cout(cout_25[43]),
    .sum(sum_25[43]));
  AL_FADD comp25_44 (
    .a(1'b0),
    .b(sum_24[44]),
    .c(cout_25[43]),
    .cout(cout_25[44]),
    .sum(sum_25[44]));
  AL_FADD comp25_45 (
    .a(1'b0),
    .b(sum_24[45]),
    .c(cout_25[44]),
    .cout(cout_25[45]),
    .sum(sum_25[45]));
  AL_FADD comp25_46 (
    .a(1'b0),
    .b(sum_24[46]),
    .c(cout_25[45]),
    .cout(cout_25[46]),
    .sum(sum_25[46]));
  AL_FADD comp25_47 (
    .a(1'b0),
    .b(sum_24[47]),
    .c(cout_25[46]),
    .cout(cout_25[47]),
    .sum(sum_25[47]));
  AL_FADD comp25_48 (
    .a(1'b0),
    .b(sum_24[48]),
    .c(cout_25[47]),
    .cout(cout_25[48]),
    .sum(sum_25[48]));
  AL_FADD comp25_49 (
    .a(1'b0),
    .b(sum_24[49]),
    .c(cout_25[48]),
    .cout(cout_25[49]),
    .sum(sum_25[49]));
  AL_FADD comp25_5 (
    .a(i25[5]),
    .b(sum_24[5]),
    .c(cout_25[4]),
    .cout(cout_25[5]),
    .sum(sum_25[5]));
  AL_FADD comp25_50 (
    .a(1'b0),
    .b(sum_24[50]),
    .c(cout_25[49]),
    .cout(cout_25[50]),
    .sum(sum_25[50]));
  AL_FADD comp25_51 (
    .a(1'b0),
    .b(sum_24[51]),
    .c(cout_25[50]),
    .cout(cout_25[51]),
    .sum(sum_25[51]));
  AL_FADD comp25_52 (
    .a(1'b0),
    .b(sum_24[52]),
    .c(cout_25[51]),
    .cout(cout_25[52]),
    .sum(sum_25[52]));
  AL_FADD comp25_53 (
    .a(1'b0),
    .b(sum_24[53]),
    .c(cout_25[52]),
    .cout(cout_25[53]),
    .sum(sum_25[53]));
  AL_FADD comp25_54 (
    .a(1'b0),
    .b(sum_24[54]),
    .c(cout_25[53]),
    .cout(cout_25[54]),
    .sum(sum_25[54]));
  AL_FADD comp25_55 (
    .a(1'b0),
    .b(sum_24[55]),
    .c(cout_25[54]),
    .cout(cout_25[55]),
    .sum(sum_25[55]));
  AL_FADD comp25_56 (
    .a(1'b0),
    .b(sum_24[56]),
    .c(cout_25[55]),
    .cout(cout_25[56]),
    .sum(sum_25[56]));
  AL_FADD comp25_57 (
    .a(1'b0),
    .b(sum_24[57]),
    .c(cout_25[56]),
    .cout(cout_25[57]),
    .sum(sum_25[57]));
  AL_FADD comp25_58 (
    .a(1'b0),
    .b(sum_24[58]),
    .c(cout_25[57]),
    .cout(cout_25[58]),
    .sum(sum_25[58]));
  AL_FADD comp25_59 (
    .a(1'b0),
    .b(sum_24[59]),
    .c(cout_25[58]),
    .cout(cout_25[59]),
    .sum(sum_25[59]));
  AL_FADD comp25_6 (
    .a(i25[6]),
    .b(sum_24[6]),
    .c(cout_25[5]),
    .cout(cout_25[6]),
    .sum(sum_25[6]));
  AL_FADD comp25_60 (
    .a(1'b0),
    .b(sum_24[60]),
    .c(cout_25[59]),
    .cout(cout_25[60]),
    .sum(sum_25[60]));
  AL_FADD comp25_61 (
    .a(1'b0),
    .b(sum_24[61]),
    .c(cout_25[60]),
    .cout(cout_25[61]),
    .sum(sum_25[61]));
  AL_FADD comp25_62 (
    .a(1'b0),
    .b(sum_24[62]),
    .c(cout_25[61]),
    .cout(cout_25[62]),
    .sum(sum_25[62]));
  AL_FADD comp25_63 (
    .a(1'b0),
    .b(sum_24[63]),
    .c(cout_25[62]),
    .cout(cout_25[63]),
    .sum(sum_25[63]));
  AL_FADD comp25_7 (
    .a(i25[7]),
    .b(sum_24[7]),
    .c(cout_25[6]),
    .cout(cout_25[7]),
    .sum(sum_25[7]));
  AL_FADD comp25_8 (
    .a(i25[8]),
    .b(sum_24[8]),
    .c(cout_25[7]),
    .cout(cout_25[8]),
    .sum(sum_25[8]));
  AL_FADD comp25_9 (
    .a(i25[9]),
    .b(sum_24[9]),
    .c(cout_25[8]),
    .cout(cout_25[9]),
    .sum(sum_25[9]));
  AL_FADD comp26_0 (
    .a(i26[0]),
    .b(sum_25[0]),
    .c(1'b0),
    .cout(cout_26[0]),
    .sum(sum_26[0]));
  AL_FADD comp26_1 (
    .a(i26[1]),
    .b(sum_25[1]),
    .c(cout_26[0]),
    .cout(cout_26[1]),
    .sum(sum_26[1]));
  AL_FADD comp26_10 (
    .a(i26[10]),
    .b(sum_25[10]),
    .c(cout_26[9]),
    .cout(cout_26[10]),
    .sum(sum_26[10]));
  AL_FADD comp26_11 (
    .a(i26[11]),
    .b(sum_25[11]),
    .c(cout_26[10]),
    .cout(cout_26[11]),
    .sum(sum_26[11]));
  AL_FADD comp26_12 (
    .a(i26[12]),
    .b(sum_25[12]),
    .c(cout_26[11]),
    .cout(cout_26[12]),
    .sum(sum_26[12]));
  AL_FADD comp26_13 (
    .a(i26[13]),
    .b(sum_25[13]),
    .c(cout_26[12]),
    .cout(cout_26[13]),
    .sum(sum_26[13]));
  AL_FADD comp26_14 (
    .a(i26[14]),
    .b(sum_25[14]),
    .c(cout_26[13]),
    .cout(cout_26[14]),
    .sum(sum_26[14]));
  AL_FADD comp26_15 (
    .a(i26[15]),
    .b(sum_25[15]),
    .c(cout_26[14]),
    .cout(cout_26[15]),
    .sum(sum_26[15]));
  AL_FADD comp26_16 (
    .a(i26[16]),
    .b(sum_25[16]),
    .c(cout_26[15]),
    .cout(cout_26[16]),
    .sum(sum_26[16]));
  AL_FADD comp26_17 (
    .a(i26[17]),
    .b(sum_25[17]),
    .c(cout_26[16]),
    .cout(cout_26[17]),
    .sum(sum_26[17]));
  AL_FADD comp26_18 (
    .a(i26[18]),
    .b(sum_25[18]),
    .c(cout_26[17]),
    .cout(cout_26[18]),
    .sum(sum_26[18]));
  AL_FADD comp26_19 (
    .a(i26[19]),
    .b(sum_25[19]),
    .c(cout_26[18]),
    .cout(cout_26[19]),
    .sum(sum_26[19]));
  AL_FADD comp26_2 (
    .a(i26[2]),
    .b(sum_25[2]),
    .c(cout_26[1]),
    .cout(cout_26[2]),
    .sum(sum_26[2]));
  AL_FADD comp26_20 (
    .a(i26[20]),
    .b(sum_25[20]),
    .c(cout_26[19]),
    .cout(cout_26[20]),
    .sum(sum_26[20]));
  AL_FADD comp26_21 (
    .a(i26[21]),
    .b(sum_25[21]),
    .c(cout_26[20]),
    .cout(cout_26[21]),
    .sum(sum_26[21]));
  AL_FADD comp26_22 (
    .a(i26[22]),
    .b(sum_25[22]),
    .c(cout_26[21]),
    .cout(cout_26[22]),
    .sum(sum_26[22]));
  AL_FADD comp26_23 (
    .a(i26[23]),
    .b(sum_25[23]),
    .c(cout_26[22]),
    .cout(cout_26[23]),
    .sum(sum_26[23]));
  AL_FADD comp26_24 (
    .a(i26[24]),
    .b(sum_25[24]),
    .c(cout_26[23]),
    .cout(cout_26[24]),
    .sum(sum_26[24]));
  AL_FADD comp26_25 (
    .a(i26[25]),
    .b(sum_25[25]),
    .c(cout_26[24]),
    .cout(cout_26[25]),
    .sum(sum_26[25]));
  AL_FADD comp26_26 (
    .a(i26[26]),
    .b(sum_25[26]),
    .c(cout_26[25]),
    .cout(cout_26[26]),
    .sum(sum_26[26]));
  AL_FADD comp26_27 (
    .a(i26[27]),
    .b(sum_25[27]),
    .c(cout_26[26]),
    .cout(cout_26[27]),
    .sum(sum_26[27]));
  AL_FADD comp26_28 (
    .a(i26[28]),
    .b(sum_25[28]),
    .c(cout_26[27]),
    .cout(cout_26[28]),
    .sum(sum_26[28]));
  AL_FADD comp26_29 (
    .a(i26[29]),
    .b(sum_25[29]),
    .c(cout_26[28]),
    .cout(cout_26[29]),
    .sum(sum_26[29]));
  AL_FADD comp26_3 (
    .a(i26[3]),
    .b(sum_25[3]),
    .c(cout_26[2]),
    .cout(cout_26[3]),
    .sum(sum_26[3]));
  AL_FADD comp26_30 (
    .a(i26[30]),
    .b(sum_25[30]),
    .c(cout_26[29]),
    .cout(cout_26[30]),
    .sum(sum_26[30]));
  AL_FADD comp26_31 (
    .a(i26[31]),
    .b(sum_25[31]),
    .c(cout_26[30]),
    .cout(cout_26[31]),
    .sum(sum_26[31]));
  AL_FADD comp26_32 (
    .a(i26[32]),
    .b(sum_25[32]),
    .c(cout_26[31]),
    .cout(cout_26[32]),
    .sum(sum_26[32]));
  AL_FADD comp26_33 (
    .a(i26[33]),
    .b(sum_25[33]),
    .c(cout_26[32]),
    .cout(cout_26[33]),
    .sum(sum_26[33]));
  AL_FADD comp26_34 (
    .a(i26[34]),
    .b(sum_25[34]),
    .c(cout_26[33]),
    .cout(cout_26[34]),
    .sum(sum_26[34]));
  AL_FADD comp26_35 (
    .a(i26[35]),
    .b(sum_25[35]),
    .c(cout_26[34]),
    .cout(cout_26[35]),
    .sum(sum_26[35]));
  AL_FADD comp26_36 (
    .a(1'b0),
    .b(sum_25[36]),
    .c(cout_26[35]),
    .cout(cout_26[36]),
    .sum(sum_26[36]));
  AL_FADD comp26_37 (
    .a(1'b0),
    .b(sum_25[37]),
    .c(cout_26[36]),
    .cout(cout_26[37]),
    .sum(sum_26[37]));
  AL_FADD comp26_38 (
    .a(1'b0),
    .b(sum_25[38]),
    .c(cout_26[37]),
    .cout(cout_26[38]),
    .sum(sum_26[38]));
  AL_FADD comp26_39 (
    .a(1'b0),
    .b(sum_25[39]),
    .c(cout_26[38]),
    .cout(cout_26[39]),
    .sum(sum_26[39]));
  AL_FADD comp26_4 (
    .a(i26[4]),
    .b(sum_25[4]),
    .c(cout_26[3]),
    .cout(cout_26[4]),
    .sum(sum_26[4]));
  AL_FADD comp26_40 (
    .a(1'b0),
    .b(sum_25[40]),
    .c(cout_26[39]),
    .cout(cout_26[40]),
    .sum(sum_26[40]));
  AL_FADD comp26_41 (
    .a(1'b0),
    .b(sum_25[41]),
    .c(cout_26[40]),
    .cout(cout_26[41]),
    .sum(sum_26[41]));
  AL_FADD comp26_42 (
    .a(1'b0),
    .b(sum_25[42]),
    .c(cout_26[41]),
    .cout(cout_26[42]),
    .sum(sum_26[42]));
  AL_FADD comp26_43 (
    .a(1'b0),
    .b(sum_25[43]),
    .c(cout_26[42]),
    .cout(cout_26[43]),
    .sum(sum_26[43]));
  AL_FADD comp26_44 (
    .a(1'b0),
    .b(sum_25[44]),
    .c(cout_26[43]),
    .cout(cout_26[44]),
    .sum(sum_26[44]));
  AL_FADD comp26_45 (
    .a(1'b0),
    .b(sum_25[45]),
    .c(cout_26[44]),
    .cout(cout_26[45]),
    .sum(sum_26[45]));
  AL_FADD comp26_46 (
    .a(1'b0),
    .b(sum_25[46]),
    .c(cout_26[45]),
    .cout(cout_26[46]),
    .sum(sum_26[46]));
  AL_FADD comp26_47 (
    .a(1'b0),
    .b(sum_25[47]),
    .c(cout_26[46]),
    .cout(cout_26[47]),
    .sum(sum_26[47]));
  AL_FADD comp26_48 (
    .a(1'b0),
    .b(sum_25[48]),
    .c(cout_26[47]),
    .cout(cout_26[48]),
    .sum(sum_26[48]));
  AL_FADD comp26_49 (
    .a(1'b0),
    .b(sum_25[49]),
    .c(cout_26[48]),
    .cout(cout_26[49]),
    .sum(sum_26[49]));
  AL_FADD comp26_5 (
    .a(i26[5]),
    .b(sum_25[5]),
    .c(cout_26[4]),
    .cout(cout_26[5]),
    .sum(sum_26[5]));
  AL_FADD comp26_50 (
    .a(1'b0),
    .b(sum_25[50]),
    .c(cout_26[49]),
    .cout(cout_26[50]),
    .sum(sum_26[50]));
  AL_FADD comp26_51 (
    .a(1'b0),
    .b(sum_25[51]),
    .c(cout_26[50]),
    .cout(cout_26[51]),
    .sum(sum_26[51]));
  AL_FADD comp26_52 (
    .a(1'b0),
    .b(sum_25[52]),
    .c(cout_26[51]),
    .cout(cout_26[52]),
    .sum(sum_26[52]));
  AL_FADD comp26_53 (
    .a(1'b0),
    .b(sum_25[53]),
    .c(cout_26[52]),
    .cout(cout_26[53]),
    .sum(sum_26[53]));
  AL_FADD comp26_54 (
    .a(1'b0),
    .b(sum_25[54]),
    .c(cout_26[53]),
    .cout(cout_26[54]),
    .sum(sum_26[54]));
  AL_FADD comp26_55 (
    .a(1'b0),
    .b(sum_25[55]),
    .c(cout_26[54]),
    .cout(cout_26[55]),
    .sum(sum_26[55]));
  AL_FADD comp26_56 (
    .a(1'b0),
    .b(sum_25[56]),
    .c(cout_26[55]),
    .cout(cout_26[56]),
    .sum(sum_26[56]));
  AL_FADD comp26_57 (
    .a(1'b0),
    .b(sum_25[57]),
    .c(cout_26[56]),
    .cout(cout_26[57]),
    .sum(sum_26[57]));
  AL_FADD comp26_58 (
    .a(1'b0),
    .b(sum_25[58]),
    .c(cout_26[57]),
    .cout(cout_26[58]),
    .sum(sum_26[58]));
  AL_FADD comp26_59 (
    .a(1'b0),
    .b(sum_25[59]),
    .c(cout_26[58]),
    .cout(cout_26[59]),
    .sum(sum_26[59]));
  AL_FADD comp26_6 (
    .a(i26[6]),
    .b(sum_25[6]),
    .c(cout_26[5]),
    .cout(cout_26[6]),
    .sum(sum_26[6]));
  AL_FADD comp26_60 (
    .a(1'b0),
    .b(sum_25[60]),
    .c(cout_26[59]),
    .cout(cout_26[60]),
    .sum(sum_26[60]));
  AL_FADD comp26_61 (
    .a(1'b0),
    .b(sum_25[61]),
    .c(cout_26[60]),
    .cout(cout_26[61]),
    .sum(sum_26[61]));
  AL_FADD comp26_62 (
    .a(1'b0),
    .b(sum_25[62]),
    .c(cout_26[61]),
    .cout(cout_26[62]),
    .sum(sum_26[62]));
  AL_FADD comp26_63 (
    .a(1'b0),
    .b(sum_25[63]),
    .c(cout_26[62]),
    .cout(cout_26[63]),
    .sum(sum_26[63]));
  AL_FADD comp26_7 (
    .a(i26[7]),
    .b(sum_25[7]),
    .c(cout_26[6]),
    .cout(cout_26[7]),
    .sum(sum_26[7]));
  AL_FADD comp26_8 (
    .a(i26[8]),
    .b(sum_25[8]),
    .c(cout_26[7]),
    .cout(cout_26[8]),
    .sum(sum_26[8]));
  AL_FADD comp26_9 (
    .a(i26[9]),
    .b(sum_25[9]),
    .c(cout_26[8]),
    .cout(cout_26[9]),
    .sum(sum_26[9]));
  AL_FADD comp27_0 (
    .a(i27[0]),
    .b(sum_26[0]),
    .c(1'b0),
    .cout(cout_27[0]),
    .sum(sum_27[0]));
  AL_FADD comp27_1 (
    .a(i27[1]),
    .b(sum_26[1]),
    .c(cout_27[0]),
    .cout(cout_27[1]),
    .sum(sum_27[1]));
  AL_FADD comp27_10 (
    .a(i27[10]),
    .b(sum_26[10]),
    .c(cout_27[9]),
    .cout(cout_27[10]),
    .sum(sum_27[10]));
  AL_FADD comp27_11 (
    .a(i27[11]),
    .b(sum_26[11]),
    .c(cout_27[10]),
    .cout(cout_27[11]),
    .sum(sum_27[11]));
  AL_FADD comp27_12 (
    .a(i27[12]),
    .b(sum_26[12]),
    .c(cout_27[11]),
    .cout(cout_27[12]),
    .sum(sum_27[12]));
  AL_FADD comp27_13 (
    .a(i27[13]),
    .b(sum_26[13]),
    .c(cout_27[12]),
    .cout(cout_27[13]),
    .sum(sum_27[13]));
  AL_FADD comp27_14 (
    .a(i27[14]),
    .b(sum_26[14]),
    .c(cout_27[13]),
    .cout(cout_27[14]),
    .sum(sum_27[14]));
  AL_FADD comp27_15 (
    .a(i27[15]),
    .b(sum_26[15]),
    .c(cout_27[14]),
    .cout(cout_27[15]),
    .sum(sum_27[15]));
  AL_FADD comp27_16 (
    .a(i27[16]),
    .b(sum_26[16]),
    .c(cout_27[15]),
    .cout(cout_27[16]),
    .sum(sum_27[16]));
  AL_FADD comp27_17 (
    .a(i27[17]),
    .b(sum_26[17]),
    .c(cout_27[16]),
    .cout(cout_27[17]),
    .sum(sum_27[17]));
  AL_FADD comp27_18 (
    .a(i27[18]),
    .b(sum_26[18]),
    .c(cout_27[17]),
    .cout(cout_27[18]),
    .sum(sum_27[18]));
  AL_FADD comp27_19 (
    .a(i27[19]),
    .b(sum_26[19]),
    .c(cout_27[18]),
    .cout(cout_27[19]),
    .sum(sum_27[19]));
  AL_FADD comp27_2 (
    .a(i27[2]),
    .b(sum_26[2]),
    .c(cout_27[1]),
    .cout(cout_27[2]),
    .sum(sum_27[2]));
  AL_FADD comp27_20 (
    .a(i27[20]),
    .b(sum_26[20]),
    .c(cout_27[19]),
    .cout(cout_27[20]),
    .sum(sum_27[20]));
  AL_FADD comp27_21 (
    .a(i27[21]),
    .b(sum_26[21]),
    .c(cout_27[20]),
    .cout(cout_27[21]),
    .sum(sum_27[21]));
  AL_FADD comp27_22 (
    .a(i27[22]),
    .b(sum_26[22]),
    .c(cout_27[21]),
    .cout(cout_27[22]),
    .sum(sum_27[22]));
  AL_FADD comp27_23 (
    .a(i27[23]),
    .b(sum_26[23]),
    .c(cout_27[22]),
    .cout(cout_27[23]),
    .sum(sum_27[23]));
  AL_FADD comp27_24 (
    .a(i27[24]),
    .b(sum_26[24]),
    .c(cout_27[23]),
    .cout(cout_27[24]),
    .sum(sum_27[24]));
  AL_FADD comp27_25 (
    .a(i27[25]),
    .b(sum_26[25]),
    .c(cout_27[24]),
    .cout(cout_27[25]),
    .sum(sum_27[25]));
  AL_FADD comp27_26 (
    .a(i27[26]),
    .b(sum_26[26]),
    .c(cout_27[25]),
    .cout(cout_27[26]),
    .sum(sum_27[26]));
  AL_FADD comp27_27 (
    .a(i27[27]),
    .b(sum_26[27]),
    .c(cout_27[26]),
    .cout(cout_27[27]),
    .sum(sum_27[27]));
  AL_FADD comp27_28 (
    .a(i27[28]),
    .b(sum_26[28]),
    .c(cout_27[27]),
    .cout(cout_27[28]),
    .sum(sum_27[28]));
  AL_FADD comp27_29 (
    .a(i27[29]),
    .b(sum_26[29]),
    .c(cout_27[28]),
    .cout(cout_27[29]),
    .sum(sum_27[29]));
  AL_FADD comp27_3 (
    .a(i27[3]),
    .b(sum_26[3]),
    .c(cout_27[2]),
    .cout(cout_27[3]),
    .sum(sum_27[3]));
  AL_FADD comp27_30 (
    .a(i27[30]),
    .b(sum_26[30]),
    .c(cout_27[29]),
    .cout(cout_27[30]),
    .sum(sum_27[30]));
  AL_FADD comp27_31 (
    .a(i27[31]),
    .b(sum_26[31]),
    .c(cout_27[30]),
    .cout(cout_27[31]),
    .sum(sum_27[31]));
  AL_FADD comp27_32 (
    .a(i27[32]),
    .b(sum_26[32]),
    .c(cout_27[31]),
    .cout(cout_27[32]),
    .sum(sum_27[32]));
  AL_FADD comp27_33 (
    .a(i27[33]),
    .b(sum_26[33]),
    .c(cout_27[32]),
    .cout(cout_27[33]),
    .sum(sum_27[33]));
  AL_FADD comp27_34 (
    .a(i27[34]),
    .b(sum_26[34]),
    .c(cout_27[33]),
    .cout(cout_27[34]),
    .sum(sum_27[34]));
  AL_FADD comp27_35 (
    .a(1'b0),
    .b(sum_26[35]),
    .c(cout_27[34]),
    .cout(cout_27[35]),
    .sum(sum_27[35]));
  AL_FADD comp27_36 (
    .a(1'b0),
    .b(sum_26[36]),
    .c(cout_27[35]),
    .cout(cout_27[36]),
    .sum(sum_27[36]));
  AL_FADD comp27_37 (
    .a(1'b0),
    .b(sum_26[37]),
    .c(cout_27[36]),
    .cout(cout_27[37]),
    .sum(sum_27[37]));
  AL_FADD comp27_38 (
    .a(1'b0),
    .b(sum_26[38]),
    .c(cout_27[37]),
    .cout(cout_27[38]),
    .sum(sum_27[38]));
  AL_FADD comp27_39 (
    .a(1'b0),
    .b(sum_26[39]),
    .c(cout_27[38]),
    .cout(cout_27[39]),
    .sum(sum_27[39]));
  AL_FADD comp27_4 (
    .a(i27[4]),
    .b(sum_26[4]),
    .c(cout_27[3]),
    .cout(cout_27[4]),
    .sum(sum_27[4]));
  AL_FADD comp27_40 (
    .a(1'b0),
    .b(sum_26[40]),
    .c(cout_27[39]),
    .cout(cout_27[40]),
    .sum(sum_27[40]));
  AL_FADD comp27_41 (
    .a(1'b0),
    .b(sum_26[41]),
    .c(cout_27[40]),
    .cout(cout_27[41]),
    .sum(sum_27[41]));
  AL_FADD comp27_42 (
    .a(1'b0),
    .b(sum_26[42]),
    .c(cout_27[41]),
    .cout(cout_27[42]),
    .sum(sum_27[42]));
  AL_FADD comp27_43 (
    .a(1'b0),
    .b(sum_26[43]),
    .c(cout_27[42]),
    .cout(cout_27[43]),
    .sum(sum_27[43]));
  AL_FADD comp27_44 (
    .a(1'b0),
    .b(sum_26[44]),
    .c(cout_27[43]),
    .cout(cout_27[44]),
    .sum(sum_27[44]));
  AL_FADD comp27_45 (
    .a(1'b0),
    .b(sum_26[45]),
    .c(cout_27[44]),
    .cout(cout_27[45]),
    .sum(sum_27[45]));
  AL_FADD comp27_46 (
    .a(1'b0),
    .b(sum_26[46]),
    .c(cout_27[45]),
    .cout(cout_27[46]),
    .sum(sum_27[46]));
  AL_FADD comp27_47 (
    .a(1'b0),
    .b(sum_26[47]),
    .c(cout_27[46]),
    .cout(cout_27[47]),
    .sum(sum_27[47]));
  AL_FADD comp27_48 (
    .a(1'b0),
    .b(sum_26[48]),
    .c(cout_27[47]),
    .cout(cout_27[48]),
    .sum(sum_27[48]));
  AL_FADD comp27_49 (
    .a(1'b0),
    .b(sum_26[49]),
    .c(cout_27[48]),
    .cout(cout_27[49]),
    .sum(sum_27[49]));
  AL_FADD comp27_5 (
    .a(i27[5]),
    .b(sum_26[5]),
    .c(cout_27[4]),
    .cout(cout_27[5]),
    .sum(sum_27[5]));
  AL_FADD comp27_50 (
    .a(1'b0),
    .b(sum_26[50]),
    .c(cout_27[49]),
    .cout(cout_27[50]),
    .sum(sum_27[50]));
  AL_FADD comp27_51 (
    .a(1'b0),
    .b(sum_26[51]),
    .c(cout_27[50]),
    .cout(cout_27[51]),
    .sum(sum_27[51]));
  AL_FADD comp27_52 (
    .a(1'b0),
    .b(sum_26[52]),
    .c(cout_27[51]),
    .cout(cout_27[52]),
    .sum(sum_27[52]));
  AL_FADD comp27_53 (
    .a(1'b0),
    .b(sum_26[53]),
    .c(cout_27[52]),
    .cout(cout_27[53]),
    .sum(sum_27[53]));
  AL_FADD comp27_54 (
    .a(1'b0),
    .b(sum_26[54]),
    .c(cout_27[53]),
    .cout(cout_27[54]),
    .sum(sum_27[54]));
  AL_FADD comp27_55 (
    .a(1'b0),
    .b(sum_26[55]),
    .c(cout_27[54]),
    .cout(cout_27[55]),
    .sum(sum_27[55]));
  AL_FADD comp27_56 (
    .a(1'b0),
    .b(sum_26[56]),
    .c(cout_27[55]),
    .cout(cout_27[56]),
    .sum(sum_27[56]));
  AL_FADD comp27_57 (
    .a(1'b0),
    .b(sum_26[57]),
    .c(cout_27[56]),
    .cout(cout_27[57]),
    .sum(sum_27[57]));
  AL_FADD comp27_58 (
    .a(1'b0),
    .b(sum_26[58]),
    .c(cout_27[57]),
    .cout(cout_27[58]),
    .sum(sum_27[58]));
  AL_FADD comp27_59 (
    .a(1'b0),
    .b(sum_26[59]),
    .c(cout_27[58]),
    .cout(cout_27[59]),
    .sum(sum_27[59]));
  AL_FADD comp27_6 (
    .a(i27[6]),
    .b(sum_26[6]),
    .c(cout_27[5]),
    .cout(cout_27[6]),
    .sum(sum_27[6]));
  AL_FADD comp27_60 (
    .a(1'b0),
    .b(sum_26[60]),
    .c(cout_27[59]),
    .cout(cout_27[60]),
    .sum(sum_27[60]));
  AL_FADD comp27_61 (
    .a(1'b0),
    .b(sum_26[61]),
    .c(cout_27[60]),
    .cout(cout_27[61]),
    .sum(sum_27[61]));
  AL_FADD comp27_62 (
    .a(1'b0),
    .b(sum_26[62]),
    .c(cout_27[61]),
    .cout(cout_27[62]),
    .sum(sum_27[62]));
  AL_FADD comp27_63 (
    .a(1'b0),
    .b(sum_26[63]),
    .c(cout_27[62]),
    .cout(cout_27[63]),
    .sum(sum_27[63]));
  AL_FADD comp27_7 (
    .a(i27[7]),
    .b(sum_26[7]),
    .c(cout_27[6]),
    .cout(cout_27[7]),
    .sum(sum_27[7]));
  AL_FADD comp27_8 (
    .a(i27[8]),
    .b(sum_26[8]),
    .c(cout_27[7]),
    .cout(cout_27[8]),
    .sum(sum_27[8]));
  AL_FADD comp27_9 (
    .a(i27[9]),
    .b(sum_26[9]),
    .c(cout_27[8]),
    .cout(cout_27[9]),
    .sum(sum_27[9]));
  AL_FADD comp28_0 (
    .a(i28[0]),
    .b(sum_27[0]),
    .c(1'b0),
    .cout(cout_28[0]),
    .sum(sum_28[0]));
  AL_FADD comp28_1 (
    .a(i28[1]),
    .b(sum_27[1]),
    .c(cout_28[0]),
    .cout(cout_28[1]),
    .sum(sum_28[1]));
  AL_FADD comp28_10 (
    .a(i28[10]),
    .b(sum_27[10]),
    .c(cout_28[9]),
    .cout(cout_28[10]),
    .sum(sum_28[10]));
  AL_FADD comp28_11 (
    .a(i28[11]),
    .b(sum_27[11]),
    .c(cout_28[10]),
    .cout(cout_28[11]),
    .sum(sum_28[11]));
  AL_FADD comp28_12 (
    .a(i28[12]),
    .b(sum_27[12]),
    .c(cout_28[11]),
    .cout(cout_28[12]),
    .sum(sum_28[12]));
  AL_FADD comp28_13 (
    .a(i28[13]),
    .b(sum_27[13]),
    .c(cout_28[12]),
    .cout(cout_28[13]),
    .sum(sum_28[13]));
  AL_FADD comp28_14 (
    .a(i28[14]),
    .b(sum_27[14]),
    .c(cout_28[13]),
    .cout(cout_28[14]),
    .sum(sum_28[14]));
  AL_FADD comp28_15 (
    .a(i28[15]),
    .b(sum_27[15]),
    .c(cout_28[14]),
    .cout(cout_28[15]),
    .sum(sum_28[15]));
  AL_FADD comp28_16 (
    .a(i28[16]),
    .b(sum_27[16]),
    .c(cout_28[15]),
    .cout(cout_28[16]),
    .sum(sum_28[16]));
  AL_FADD comp28_17 (
    .a(i28[17]),
    .b(sum_27[17]),
    .c(cout_28[16]),
    .cout(cout_28[17]),
    .sum(sum_28[17]));
  AL_FADD comp28_18 (
    .a(i28[18]),
    .b(sum_27[18]),
    .c(cout_28[17]),
    .cout(cout_28[18]),
    .sum(sum_28[18]));
  AL_FADD comp28_19 (
    .a(i28[19]),
    .b(sum_27[19]),
    .c(cout_28[18]),
    .cout(cout_28[19]),
    .sum(sum_28[19]));
  AL_FADD comp28_2 (
    .a(i28[2]),
    .b(sum_27[2]),
    .c(cout_28[1]),
    .cout(cout_28[2]),
    .sum(sum_28[2]));
  AL_FADD comp28_20 (
    .a(i28[20]),
    .b(sum_27[20]),
    .c(cout_28[19]),
    .cout(cout_28[20]),
    .sum(sum_28[20]));
  AL_FADD comp28_21 (
    .a(i28[21]),
    .b(sum_27[21]),
    .c(cout_28[20]),
    .cout(cout_28[21]),
    .sum(sum_28[21]));
  AL_FADD comp28_22 (
    .a(i28[22]),
    .b(sum_27[22]),
    .c(cout_28[21]),
    .cout(cout_28[22]),
    .sum(sum_28[22]));
  AL_FADD comp28_23 (
    .a(i28[23]),
    .b(sum_27[23]),
    .c(cout_28[22]),
    .cout(cout_28[23]),
    .sum(sum_28[23]));
  AL_FADD comp28_24 (
    .a(i28[24]),
    .b(sum_27[24]),
    .c(cout_28[23]),
    .cout(cout_28[24]),
    .sum(sum_28[24]));
  AL_FADD comp28_25 (
    .a(i28[25]),
    .b(sum_27[25]),
    .c(cout_28[24]),
    .cout(cout_28[25]),
    .sum(sum_28[25]));
  AL_FADD comp28_26 (
    .a(i28[26]),
    .b(sum_27[26]),
    .c(cout_28[25]),
    .cout(cout_28[26]),
    .sum(sum_28[26]));
  AL_FADD comp28_27 (
    .a(i28[27]),
    .b(sum_27[27]),
    .c(cout_28[26]),
    .cout(cout_28[27]),
    .sum(sum_28[27]));
  AL_FADD comp28_28 (
    .a(i28[28]),
    .b(sum_27[28]),
    .c(cout_28[27]),
    .cout(cout_28[28]),
    .sum(sum_28[28]));
  AL_FADD comp28_29 (
    .a(i28[29]),
    .b(sum_27[29]),
    .c(cout_28[28]),
    .cout(cout_28[29]),
    .sum(sum_28[29]));
  AL_FADD comp28_3 (
    .a(i28[3]),
    .b(sum_27[3]),
    .c(cout_28[2]),
    .cout(cout_28[3]),
    .sum(sum_28[3]));
  AL_FADD comp28_30 (
    .a(i28[30]),
    .b(sum_27[30]),
    .c(cout_28[29]),
    .cout(cout_28[30]),
    .sum(sum_28[30]));
  AL_FADD comp28_31 (
    .a(i28[31]),
    .b(sum_27[31]),
    .c(cout_28[30]),
    .cout(cout_28[31]),
    .sum(sum_28[31]));
  AL_FADD comp28_32 (
    .a(i28[32]),
    .b(sum_27[32]),
    .c(cout_28[31]),
    .cout(cout_28[32]),
    .sum(sum_28[32]));
  AL_FADD comp28_33 (
    .a(i28[33]),
    .b(sum_27[33]),
    .c(cout_28[32]),
    .cout(cout_28[33]),
    .sum(sum_28[33]));
  AL_FADD comp28_34 (
    .a(1'b0),
    .b(sum_27[34]),
    .c(cout_28[33]),
    .cout(cout_28[34]),
    .sum(sum_28[34]));
  AL_FADD comp28_35 (
    .a(1'b0),
    .b(sum_27[35]),
    .c(cout_28[34]),
    .cout(cout_28[35]),
    .sum(sum_28[35]));
  AL_FADD comp28_36 (
    .a(1'b0),
    .b(sum_27[36]),
    .c(cout_28[35]),
    .cout(cout_28[36]),
    .sum(sum_28[36]));
  AL_FADD comp28_37 (
    .a(1'b0),
    .b(sum_27[37]),
    .c(cout_28[36]),
    .cout(cout_28[37]),
    .sum(sum_28[37]));
  AL_FADD comp28_38 (
    .a(1'b0),
    .b(sum_27[38]),
    .c(cout_28[37]),
    .cout(cout_28[38]),
    .sum(sum_28[38]));
  AL_FADD comp28_39 (
    .a(1'b0),
    .b(sum_27[39]),
    .c(cout_28[38]),
    .cout(cout_28[39]),
    .sum(sum_28[39]));
  AL_FADD comp28_4 (
    .a(i28[4]),
    .b(sum_27[4]),
    .c(cout_28[3]),
    .cout(cout_28[4]),
    .sum(sum_28[4]));
  AL_FADD comp28_40 (
    .a(1'b0),
    .b(sum_27[40]),
    .c(cout_28[39]),
    .cout(cout_28[40]),
    .sum(sum_28[40]));
  AL_FADD comp28_41 (
    .a(1'b0),
    .b(sum_27[41]),
    .c(cout_28[40]),
    .cout(cout_28[41]),
    .sum(sum_28[41]));
  AL_FADD comp28_42 (
    .a(1'b0),
    .b(sum_27[42]),
    .c(cout_28[41]),
    .cout(cout_28[42]),
    .sum(sum_28[42]));
  AL_FADD comp28_43 (
    .a(1'b0),
    .b(sum_27[43]),
    .c(cout_28[42]),
    .cout(cout_28[43]),
    .sum(sum_28[43]));
  AL_FADD comp28_44 (
    .a(1'b0),
    .b(sum_27[44]),
    .c(cout_28[43]),
    .cout(cout_28[44]),
    .sum(sum_28[44]));
  AL_FADD comp28_45 (
    .a(1'b0),
    .b(sum_27[45]),
    .c(cout_28[44]),
    .cout(cout_28[45]),
    .sum(sum_28[45]));
  AL_FADD comp28_46 (
    .a(1'b0),
    .b(sum_27[46]),
    .c(cout_28[45]),
    .cout(cout_28[46]),
    .sum(sum_28[46]));
  AL_FADD comp28_47 (
    .a(1'b0),
    .b(sum_27[47]),
    .c(cout_28[46]),
    .cout(cout_28[47]),
    .sum(sum_28[47]));
  AL_FADD comp28_48 (
    .a(1'b0),
    .b(sum_27[48]),
    .c(cout_28[47]),
    .cout(cout_28[48]),
    .sum(sum_28[48]));
  AL_FADD comp28_49 (
    .a(1'b0),
    .b(sum_27[49]),
    .c(cout_28[48]),
    .cout(cout_28[49]),
    .sum(sum_28[49]));
  AL_FADD comp28_5 (
    .a(i28[5]),
    .b(sum_27[5]),
    .c(cout_28[4]),
    .cout(cout_28[5]),
    .sum(sum_28[5]));
  AL_FADD comp28_50 (
    .a(1'b0),
    .b(sum_27[50]),
    .c(cout_28[49]),
    .cout(cout_28[50]),
    .sum(sum_28[50]));
  AL_FADD comp28_51 (
    .a(1'b0),
    .b(sum_27[51]),
    .c(cout_28[50]),
    .cout(cout_28[51]),
    .sum(sum_28[51]));
  AL_FADD comp28_52 (
    .a(1'b0),
    .b(sum_27[52]),
    .c(cout_28[51]),
    .cout(cout_28[52]),
    .sum(sum_28[52]));
  AL_FADD comp28_53 (
    .a(1'b0),
    .b(sum_27[53]),
    .c(cout_28[52]),
    .cout(cout_28[53]),
    .sum(sum_28[53]));
  AL_FADD comp28_54 (
    .a(1'b0),
    .b(sum_27[54]),
    .c(cout_28[53]),
    .cout(cout_28[54]),
    .sum(sum_28[54]));
  AL_FADD comp28_55 (
    .a(1'b0),
    .b(sum_27[55]),
    .c(cout_28[54]),
    .cout(cout_28[55]),
    .sum(sum_28[55]));
  AL_FADD comp28_56 (
    .a(1'b0),
    .b(sum_27[56]),
    .c(cout_28[55]),
    .cout(cout_28[56]),
    .sum(sum_28[56]));
  AL_FADD comp28_57 (
    .a(1'b0),
    .b(sum_27[57]),
    .c(cout_28[56]),
    .cout(cout_28[57]),
    .sum(sum_28[57]));
  AL_FADD comp28_58 (
    .a(1'b0),
    .b(sum_27[58]),
    .c(cout_28[57]),
    .cout(cout_28[58]),
    .sum(sum_28[58]));
  AL_FADD comp28_59 (
    .a(1'b0),
    .b(sum_27[59]),
    .c(cout_28[58]),
    .cout(cout_28[59]),
    .sum(sum_28[59]));
  AL_FADD comp28_6 (
    .a(i28[6]),
    .b(sum_27[6]),
    .c(cout_28[5]),
    .cout(cout_28[6]),
    .sum(sum_28[6]));
  AL_FADD comp28_60 (
    .a(1'b0),
    .b(sum_27[60]),
    .c(cout_28[59]),
    .cout(cout_28[60]),
    .sum(sum_28[60]));
  AL_FADD comp28_61 (
    .a(1'b0),
    .b(sum_27[61]),
    .c(cout_28[60]),
    .cout(cout_28[61]),
    .sum(sum_28[61]));
  AL_FADD comp28_62 (
    .a(1'b0),
    .b(sum_27[62]),
    .c(cout_28[61]),
    .cout(cout_28[62]),
    .sum(sum_28[62]));
  AL_FADD comp28_63 (
    .a(1'b0),
    .b(sum_27[63]),
    .c(cout_28[62]),
    .cout(cout_28[63]),
    .sum(sum_28[63]));
  AL_FADD comp28_7 (
    .a(i28[7]),
    .b(sum_27[7]),
    .c(cout_28[6]),
    .cout(cout_28[7]),
    .sum(sum_28[7]));
  AL_FADD comp28_8 (
    .a(i28[8]),
    .b(sum_27[8]),
    .c(cout_28[7]),
    .cout(cout_28[8]),
    .sum(sum_28[8]));
  AL_FADD comp28_9 (
    .a(i28[9]),
    .b(sum_27[9]),
    .c(cout_28[8]),
    .cout(cout_28[9]),
    .sum(sum_28[9]));
  AL_FADD comp29_0 (
    .a(i29[0]),
    .b(sum_28[0]),
    .c(1'b0),
    .cout(cout_29[0]),
    .sum(sum_29[0]));
  AL_FADD comp29_1 (
    .a(i29[1]),
    .b(sum_28[1]),
    .c(cout_29[0]),
    .cout(cout_29[1]),
    .sum(sum_29[1]));
  AL_FADD comp29_10 (
    .a(i29[10]),
    .b(sum_28[10]),
    .c(cout_29[9]),
    .cout(cout_29[10]),
    .sum(sum_29[10]));
  AL_FADD comp29_11 (
    .a(i29[11]),
    .b(sum_28[11]),
    .c(cout_29[10]),
    .cout(cout_29[11]),
    .sum(sum_29[11]));
  AL_FADD comp29_12 (
    .a(i29[12]),
    .b(sum_28[12]),
    .c(cout_29[11]),
    .cout(cout_29[12]),
    .sum(sum_29[12]));
  AL_FADD comp29_13 (
    .a(i29[13]),
    .b(sum_28[13]),
    .c(cout_29[12]),
    .cout(cout_29[13]),
    .sum(sum_29[13]));
  AL_FADD comp29_14 (
    .a(i29[14]),
    .b(sum_28[14]),
    .c(cout_29[13]),
    .cout(cout_29[14]),
    .sum(sum_29[14]));
  AL_FADD comp29_15 (
    .a(i29[15]),
    .b(sum_28[15]),
    .c(cout_29[14]),
    .cout(cout_29[15]),
    .sum(sum_29[15]));
  AL_FADD comp29_16 (
    .a(i29[16]),
    .b(sum_28[16]),
    .c(cout_29[15]),
    .cout(cout_29[16]),
    .sum(sum_29[16]));
  AL_FADD comp29_17 (
    .a(i29[17]),
    .b(sum_28[17]),
    .c(cout_29[16]),
    .cout(cout_29[17]),
    .sum(sum_29[17]));
  AL_FADD comp29_18 (
    .a(i29[18]),
    .b(sum_28[18]),
    .c(cout_29[17]),
    .cout(cout_29[18]),
    .sum(sum_29[18]));
  AL_FADD comp29_19 (
    .a(i29[19]),
    .b(sum_28[19]),
    .c(cout_29[18]),
    .cout(cout_29[19]),
    .sum(sum_29[19]));
  AL_FADD comp29_2 (
    .a(i29[2]),
    .b(sum_28[2]),
    .c(cout_29[1]),
    .cout(cout_29[2]),
    .sum(sum_29[2]));
  AL_FADD comp29_20 (
    .a(i29[20]),
    .b(sum_28[20]),
    .c(cout_29[19]),
    .cout(cout_29[20]),
    .sum(sum_29[20]));
  AL_FADD comp29_21 (
    .a(i29[21]),
    .b(sum_28[21]),
    .c(cout_29[20]),
    .cout(cout_29[21]),
    .sum(sum_29[21]));
  AL_FADD comp29_22 (
    .a(i29[22]),
    .b(sum_28[22]),
    .c(cout_29[21]),
    .cout(cout_29[22]),
    .sum(sum_29[22]));
  AL_FADD comp29_23 (
    .a(i29[23]),
    .b(sum_28[23]),
    .c(cout_29[22]),
    .cout(cout_29[23]),
    .sum(sum_29[23]));
  AL_FADD comp29_24 (
    .a(i29[24]),
    .b(sum_28[24]),
    .c(cout_29[23]),
    .cout(cout_29[24]),
    .sum(sum_29[24]));
  AL_FADD comp29_25 (
    .a(i29[25]),
    .b(sum_28[25]),
    .c(cout_29[24]),
    .cout(cout_29[25]),
    .sum(sum_29[25]));
  AL_FADD comp29_26 (
    .a(i29[26]),
    .b(sum_28[26]),
    .c(cout_29[25]),
    .cout(cout_29[26]),
    .sum(sum_29[26]));
  AL_FADD comp29_27 (
    .a(i29[27]),
    .b(sum_28[27]),
    .c(cout_29[26]),
    .cout(cout_29[27]),
    .sum(sum_29[27]));
  AL_FADD comp29_28 (
    .a(i29[28]),
    .b(sum_28[28]),
    .c(cout_29[27]),
    .cout(cout_29[28]),
    .sum(sum_29[28]));
  AL_FADD comp29_29 (
    .a(i29[29]),
    .b(sum_28[29]),
    .c(cout_29[28]),
    .cout(cout_29[29]),
    .sum(sum_29[29]));
  AL_FADD comp29_3 (
    .a(i29[3]),
    .b(sum_28[3]),
    .c(cout_29[2]),
    .cout(cout_29[3]),
    .sum(sum_29[3]));
  AL_FADD comp29_30 (
    .a(i29[30]),
    .b(sum_28[30]),
    .c(cout_29[29]),
    .cout(cout_29[30]),
    .sum(sum_29[30]));
  AL_FADD comp29_31 (
    .a(i29[31]),
    .b(sum_28[31]),
    .c(cout_29[30]),
    .cout(cout_29[31]),
    .sum(sum_29[31]));
  AL_FADD comp29_32 (
    .a(i29[32]),
    .b(sum_28[32]),
    .c(cout_29[31]),
    .cout(cout_29[32]),
    .sum(sum_29[32]));
  AL_FADD comp29_33 (
    .a(1'b0),
    .b(sum_28[33]),
    .c(cout_29[32]),
    .cout(cout_29[33]),
    .sum(sum_29[33]));
  AL_FADD comp29_34 (
    .a(1'b0),
    .b(sum_28[34]),
    .c(cout_29[33]),
    .cout(cout_29[34]),
    .sum(sum_29[34]));
  AL_FADD comp29_35 (
    .a(1'b0),
    .b(sum_28[35]),
    .c(cout_29[34]),
    .cout(cout_29[35]),
    .sum(sum_29[35]));
  AL_FADD comp29_36 (
    .a(1'b0),
    .b(sum_28[36]),
    .c(cout_29[35]),
    .cout(cout_29[36]),
    .sum(sum_29[36]));
  AL_FADD comp29_37 (
    .a(1'b0),
    .b(sum_28[37]),
    .c(cout_29[36]),
    .cout(cout_29[37]),
    .sum(sum_29[37]));
  AL_FADD comp29_38 (
    .a(1'b0),
    .b(sum_28[38]),
    .c(cout_29[37]),
    .cout(cout_29[38]),
    .sum(sum_29[38]));
  AL_FADD comp29_39 (
    .a(1'b0),
    .b(sum_28[39]),
    .c(cout_29[38]),
    .cout(cout_29[39]),
    .sum(sum_29[39]));
  AL_FADD comp29_4 (
    .a(i29[4]),
    .b(sum_28[4]),
    .c(cout_29[3]),
    .cout(cout_29[4]),
    .sum(sum_29[4]));
  AL_FADD comp29_40 (
    .a(1'b0),
    .b(sum_28[40]),
    .c(cout_29[39]),
    .cout(cout_29[40]),
    .sum(sum_29[40]));
  AL_FADD comp29_41 (
    .a(1'b0),
    .b(sum_28[41]),
    .c(cout_29[40]),
    .cout(cout_29[41]),
    .sum(sum_29[41]));
  AL_FADD comp29_42 (
    .a(1'b0),
    .b(sum_28[42]),
    .c(cout_29[41]),
    .cout(cout_29[42]),
    .sum(sum_29[42]));
  AL_FADD comp29_43 (
    .a(1'b0),
    .b(sum_28[43]),
    .c(cout_29[42]),
    .cout(cout_29[43]),
    .sum(sum_29[43]));
  AL_FADD comp29_44 (
    .a(1'b0),
    .b(sum_28[44]),
    .c(cout_29[43]),
    .cout(cout_29[44]),
    .sum(sum_29[44]));
  AL_FADD comp29_45 (
    .a(1'b0),
    .b(sum_28[45]),
    .c(cout_29[44]),
    .cout(cout_29[45]),
    .sum(sum_29[45]));
  AL_FADD comp29_46 (
    .a(1'b0),
    .b(sum_28[46]),
    .c(cout_29[45]),
    .cout(cout_29[46]),
    .sum(sum_29[46]));
  AL_FADD comp29_47 (
    .a(1'b0),
    .b(sum_28[47]),
    .c(cout_29[46]),
    .cout(cout_29[47]),
    .sum(sum_29[47]));
  AL_FADD comp29_48 (
    .a(1'b0),
    .b(sum_28[48]),
    .c(cout_29[47]),
    .cout(cout_29[48]),
    .sum(sum_29[48]));
  AL_FADD comp29_49 (
    .a(1'b0),
    .b(sum_28[49]),
    .c(cout_29[48]),
    .cout(cout_29[49]),
    .sum(sum_29[49]));
  AL_FADD comp29_5 (
    .a(i29[5]),
    .b(sum_28[5]),
    .c(cout_29[4]),
    .cout(cout_29[5]),
    .sum(sum_29[5]));
  AL_FADD comp29_50 (
    .a(1'b0),
    .b(sum_28[50]),
    .c(cout_29[49]),
    .cout(cout_29[50]),
    .sum(sum_29[50]));
  AL_FADD comp29_51 (
    .a(1'b0),
    .b(sum_28[51]),
    .c(cout_29[50]),
    .cout(cout_29[51]),
    .sum(sum_29[51]));
  AL_FADD comp29_52 (
    .a(1'b0),
    .b(sum_28[52]),
    .c(cout_29[51]),
    .cout(cout_29[52]),
    .sum(sum_29[52]));
  AL_FADD comp29_53 (
    .a(1'b0),
    .b(sum_28[53]),
    .c(cout_29[52]),
    .cout(cout_29[53]),
    .sum(sum_29[53]));
  AL_FADD comp29_54 (
    .a(1'b0),
    .b(sum_28[54]),
    .c(cout_29[53]),
    .cout(cout_29[54]),
    .sum(sum_29[54]));
  AL_FADD comp29_55 (
    .a(1'b0),
    .b(sum_28[55]),
    .c(cout_29[54]),
    .cout(cout_29[55]),
    .sum(sum_29[55]));
  AL_FADD comp29_56 (
    .a(1'b0),
    .b(sum_28[56]),
    .c(cout_29[55]),
    .cout(cout_29[56]),
    .sum(sum_29[56]));
  AL_FADD comp29_57 (
    .a(1'b0),
    .b(sum_28[57]),
    .c(cout_29[56]),
    .cout(cout_29[57]),
    .sum(sum_29[57]));
  AL_FADD comp29_58 (
    .a(1'b0),
    .b(sum_28[58]),
    .c(cout_29[57]),
    .cout(cout_29[58]),
    .sum(sum_29[58]));
  AL_FADD comp29_59 (
    .a(1'b0),
    .b(sum_28[59]),
    .c(cout_29[58]),
    .cout(cout_29[59]),
    .sum(sum_29[59]));
  AL_FADD comp29_6 (
    .a(i29[6]),
    .b(sum_28[6]),
    .c(cout_29[5]),
    .cout(cout_29[6]),
    .sum(sum_29[6]));
  AL_FADD comp29_60 (
    .a(1'b0),
    .b(sum_28[60]),
    .c(cout_29[59]),
    .cout(cout_29[60]),
    .sum(sum_29[60]));
  AL_FADD comp29_61 (
    .a(1'b0),
    .b(sum_28[61]),
    .c(cout_29[60]),
    .cout(cout_29[61]),
    .sum(sum_29[61]));
  AL_FADD comp29_62 (
    .a(1'b0),
    .b(sum_28[62]),
    .c(cout_29[61]),
    .cout(cout_29[62]),
    .sum(sum_29[62]));
  AL_FADD comp29_63 (
    .a(1'b0),
    .b(sum_28[63]),
    .c(cout_29[62]),
    .cout(cout_29[63]),
    .sum(sum_29[63]));
  AL_FADD comp29_7 (
    .a(i29[7]),
    .b(sum_28[7]),
    .c(cout_29[6]),
    .cout(cout_29[7]),
    .sum(sum_29[7]));
  AL_FADD comp29_8 (
    .a(i29[8]),
    .b(sum_28[8]),
    .c(cout_29[7]),
    .cout(cout_29[8]),
    .sum(sum_29[8]));
  AL_FADD comp29_9 (
    .a(i29[9]),
    .b(sum_28[9]),
    .c(cout_29[8]),
    .cout(cout_29[9]),
    .sum(sum_29[9]));
  AL_FADD comp2_0 (
    .a(i2[0]),
    .b(sum_1[0]),
    .c(1'b0),
    .cout(cout_2[0]),
    .sum(sum_2[0]));
  AL_FADD comp2_1 (
    .a(i2[1]),
    .b(sum_1[1]),
    .c(cout_2[0]),
    .cout(cout_2[1]),
    .sum(sum_2[1]));
  AL_FADD comp2_10 (
    .a(i2[10]),
    .b(sum_1[10]),
    .c(cout_2[9]),
    .cout(cout_2[10]),
    .sum(sum_2[10]));
  AL_FADD comp2_11 (
    .a(i2[11]),
    .b(sum_1[11]),
    .c(cout_2[10]),
    .cout(cout_2[11]),
    .sum(sum_2[11]));
  AL_FADD comp2_12 (
    .a(i2[12]),
    .b(sum_1[12]),
    .c(cout_2[11]),
    .cout(cout_2[12]),
    .sum(sum_2[12]));
  AL_FADD comp2_13 (
    .a(i2[13]),
    .b(sum_1[13]),
    .c(cout_2[12]),
    .cout(cout_2[13]),
    .sum(sum_2[13]));
  AL_FADD comp2_14 (
    .a(i2[14]),
    .b(sum_1[14]),
    .c(cout_2[13]),
    .cout(cout_2[14]),
    .sum(sum_2[14]));
  AL_FADD comp2_15 (
    .a(i2[15]),
    .b(sum_1[15]),
    .c(cout_2[14]),
    .cout(cout_2[15]),
    .sum(sum_2[15]));
  AL_FADD comp2_16 (
    .a(i2[16]),
    .b(sum_1[16]),
    .c(cout_2[15]),
    .cout(cout_2[16]),
    .sum(sum_2[16]));
  AL_FADD comp2_17 (
    .a(i2[17]),
    .b(sum_1[17]),
    .c(cout_2[16]),
    .cout(cout_2[17]),
    .sum(sum_2[17]));
  AL_FADD comp2_18 (
    .a(i2[18]),
    .b(sum_1[18]),
    .c(cout_2[17]),
    .cout(cout_2[18]),
    .sum(sum_2[18]));
  AL_FADD comp2_19 (
    .a(i2[19]),
    .b(sum_1[19]),
    .c(cout_2[18]),
    .cout(cout_2[19]),
    .sum(sum_2[19]));
  AL_FADD comp2_2 (
    .a(i2[2]),
    .b(sum_1[2]),
    .c(cout_2[1]),
    .cout(cout_2[2]),
    .sum(sum_2[2]));
  AL_FADD comp2_20 (
    .a(i2[20]),
    .b(sum_1[20]),
    .c(cout_2[19]),
    .cout(cout_2[20]),
    .sum(sum_2[20]));
  AL_FADD comp2_21 (
    .a(i2[21]),
    .b(sum_1[21]),
    .c(cout_2[20]),
    .cout(cout_2[21]),
    .sum(sum_2[21]));
  AL_FADD comp2_22 (
    .a(i2[22]),
    .b(sum_1[22]),
    .c(cout_2[21]),
    .cout(cout_2[22]),
    .sum(sum_2[22]));
  AL_FADD comp2_23 (
    .a(i2[23]),
    .b(sum_1[23]),
    .c(cout_2[22]),
    .cout(cout_2[23]),
    .sum(sum_2[23]));
  AL_FADD comp2_24 (
    .a(i2[24]),
    .b(sum_1[24]),
    .c(cout_2[23]),
    .cout(cout_2[24]),
    .sum(sum_2[24]));
  AL_FADD comp2_25 (
    .a(i2[25]),
    .b(sum_1[25]),
    .c(cout_2[24]),
    .cout(cout_2[25]),
    .sum(sum_2[25]));
  AL_FADD comp2_26 (
    .a(i2[26]),
    .b(sum_1[26]),
    .c(cout_2[25]),
    .cout(cout_2[26]),
    .sum(sum_2[26]));
  AL_FADD comp2_27 (
    .a(i2[27]),
    .b(sum_1[27]),
    .c(cout_2[26]),
    .cout(cout_2[27]),
    .sum(sum_2[27]));
  AL_FADD comp2_28 (
    .a(i2[28]),
    .b(sum_1[28]),
    .c(cout_2[27]),
    .cout(cout_2[28]),
    .sum(sum_2[28]));
  AL_FADD comp2_29 (
    .a(i2[29]),
    .b(sum_1[29]),
    .c(cout_2[28]),
    .cout(cout_2[29]),
    .sum(sum_2[29]));
  AL_FADD comp2_3 (
    .a(i2[3]),
    .b(sum_1[3]),
    .c(cout_2[2]),
    .cout(cout_2[3]),
    .sum(sum_2[3]));
  AL_FADD comp2_30 (
    .a(i2[30]),
    .b(sum_1[30]),
    .c(cout_2[29]),
    .cout(cout_2[30]),
    .sum(sum_2[30]));
  AL_FADD comp2_31 (
    .a(i2[31]),
    .b(sum_1[31]),
    .c(cout_2[30]),
    .cout(cout_2[31]),
    .sum(sum_2[31]));
  AL_FADD comp2_32 (
    .a(i2[32]),
    .b(sum_1[32]),
    .c(cout_2[31]),
    .cout(cout_2[32]),
    .sum(sum_2[32]));
  AL_FADD comp2_33 (
    .a(i2[33]),
    .b(sum_1[33]),
    .c(cout_2[32]),
    .cout(cout_2[33]),
    .sum(sum_2[33]));
  AL_FADD comp2_34 (
    .a(i2[34]),
    .b(sum_1[34]),
    .c(cout_2[33]),
    .cout(cout_2[34]),
    .sum(sum_2[34]));
  AL_FADD comp2_35 (
    .a(i2[35]),
    .b(sum_1[35]),
    .c(cout_2[34]),
    .cout(cout_2[35]),
    .sum(sum_2[35]));
  AL_FADD comp2_36 (
    .a(i2[36]),
    .b(sum_1[36]),
    .c(cout_2[35]),
    .cout(cout_2[36]),
    .sum(sum_2[36]));
  AL_FADD comp2_37 (
    .a(i2[37]),
    .b(sum_1[37]),
    .c(cout_2[36]),
    .cout(cout_2[37]),
    .sum(sum_2[37]));
  AL_FADD comp2_38 (
    .a(i2[38]),
    .b(sum_1[38]),
    .c(cout_2[37]),
    .cout(cout_2[38]),
    .sum(sum_2[38]));
  AL_FADD comp2_39 (
    .a(i2[39]),
    .b(sum_1[39]),
    .c(cout_2[38]),
    .cout(cout_2[39]),
    .sum(sum_2[39]));
  AL_FADD comp2_4 (
    .a(i2[4]),
    .b(sum_1[4]),
    .c(cout_2[3]),
    .cout(cout_2[4]),
    .sum(sum_2[4]));
  AL_FADD comp2_40 (
    .a(i2[40]),
    .b(sum_1[40]),
    .c(cout_2[39]),
    .cout(cout_2[40]),
    .sum(sum_2[40]));
  AL_FADD comp2_41 (
    .a(i2[41]),
    .b(sum_1[41]),
    .c(cout_2[40]),
    .cout(cout_2[41]),
    .sum(sum_2[41]));
  AL_FADD comp2_42 (
    .a(i2[42]),
    .b(sum_1[42]),
    .c(cout_2[41]),
    .cout(cout_2[42]),
    .sum(sum_2[42]));
  AL_FADD comp2_43 (
    .a(i2[43]),
    .b(sum_1[43]),
    .c(cout_2[42]),
    .cout(cout_2[43]),
    .sum(sum_2[43]));
  AL_FADD comp2_44 (
    .a(i2[44]),
    .b(sum_1[44]),
    .c(cout_2[43]),
    .cout(cout_2[44]),
    .sum(sum_2[44]));
  AL_FADD comp2_45 (
    .a(i2[45]),
    .b(sum_1[45]),
    .c(cout_2[44]),
    .cout(cout_2[45]),
    .sum(sum_2[45]));
  AL_FADD comp2_46 (
    .a(i2[46]),
    .b(sum_1[46]),
    .c(cout_2[45]),
    .cout(cout_2[46]),
    .sum(sum_2[46]));
  AL_FADD comp2_47 (
    .a(i2[47]),
    .b(sum_1[47]),
    .c(cout_2[46]),
    .cout(cout_2[47]),
    .sum(sum_2[47]));
  AL_FADD comp2_48 (
    .a(i2[48]),
    .b(sum_1[48]),
    .c(cout_2[47]),
    .cout(cout_2[48]),
    .sum(sum_2[48]));
  AL_FADD comp2_49 (
    .a(i2[49]),
    .b(sum_1[49]),
    .c(cout_2[48]),
    .cout(cout_2[49]),
    .sum(sum_2[49]));
  AL_FADD comp2_5 (
    .a(i2[5]),
    .b(sum_1[5]),
    .c(cout_2[4]),
    .cout(cout_2[5]),
    .sum(sum_2[5]));
  AL_FADD comp2_50 (
    .a(i2[50]),
    .b(sum_1[50]),
    .c(cout_2[49]),
    .cout(cout_2[50]),
    .sum(sum_2[50]));
  AL_FADD comp2_51 (
    .a(i2[51]),
    .b(sum_1[51]),
    .c(cout_2[50]),
    .cout(cout_2[51]),
    .sum(sum_2[51]));
  AL_FADD comp2_52 (
    .a(i2[52]),
    .b(sum_1[52]),
    .c(cout_2[51]),
    .cout(cout_2[52]),
    .sum(sum_2[52]));
  AL_FADD comp2_53 (
    .a(i2[53]),
    .b(sum_1[53]),
    .c(cout_2[52]),
    .cout(cout_2[53]),
    .sum(sum_2[53]));
  AL_FADD comp2_54 (
    .a(i2[54]),
    .b(sum_1[54]),
    .c(cout_2[53]),
    .cout(cout_2[54]),
    .sum(sum_2[54]));
  AL_FADD comp2_55 (
    .a(i2[55]),
    .b(sum_1[55]),
    .c(cout_2[54]),
    .cout(cout_2[55]),
    .sum(sum_2[55]));
  AL_FADD comp2_56 (
    .a(i2[56]),
    .b(sum_1[56]),
    .c(cout_2[55]),
    .cout(cout_2[56]),
    .sum(sum_2[56]));
  AL_FADD comp2_57 (
    .a(i2[57]),
    .b(sum_1[57]),
    .c(cout_2[56]),
    .cout(cout_2[57]),
    .sum(sum_2[57]));
  AL_FADD comp2_58 (
    .a(i2[58]),
    .b(sum_1[58]),
    .c(cout_2[57]),
    .cout(cout_2[58]),
    .sum(sum_2[58]));
  AL_FADD comp2_59 (
    .a(i2[59]),
    .b(sum_1[59]),
    .c(cout_2[58]),
    .cout(cout_2[59]),
    .sum(sum_2[59]));
  AL_FADD comp2_6 (
    .a(i2[6]),
    .b(sum_1[6]),
    .c(cout_2[5]),
    .cout(cout_2[6]),
    .sum(sum_2[6]));
  AL_FADD comp2_60 (
    .a(1'b0),
    .b(sum_1[60]),
    .c(cout_2[59]),
    .cout(cout_2[60]),
    .sum(sum_2[60]));
  AL_FADD comp2_61 (
    .a(1'b0),
    .b(sum_1[61]),
    .c(cout_2[60]),
    .cout(cout_2[61]),
    .sum(sum_2[61]));
  AL_FADD comp2_62 (
    .a(1'b0),
    .b(sum_1[62]),
    .c(cout_2[61]),
    .cout(cout_2[62]),
    .sum(sum_2[62]));
  AL_FADD comp2_63 (
    .a(1'b0),
    .b(sum_1[63]),
    .c(cout_2[62]),
    .cout(cout_2[63]),
    .sum(sum_2[63]));
  AL_FADD comp2_7 (
    .a(i2[7]),
    .b(sum_1[7]),
    .c(cout_2[6]),
    .cout(cout_2[7]),
    .sum(sum_2[7]));
  AL_FADD comp2_8 (
    .a(i2[8]),
    .b(sum_1[8]),
    .c(cout_2[7]),
    .cout(cout_2[8]),
    .sum(sum_2[8]));
  AL_FADD comp2_9 (
    .a(i2[9]),
    .b(sum_1[9]),
    .c(cout_2[8]),
    .cout(cout_2[9]),
    .sum(sum_2[9]));
  AL_FADD comp30_0 (
    .a(i30[0]),
    .b(sum_29[0]),
    .c(1'b0),
    .cout(cout_30[0]),
    .sum(sum_30[0]));
  AL_FADD comp30_1 (
    .a(i30[1]),
    .b(sum_29[1]),
    .c(cout_30[0]),
    .cout(cout_30[1]),
    .sum(sum_30[1]));
  AL_FADD comp30_10 (
    .a(i30[10]),
    .b(sum_29[10]),
    .c(cout_30[9]),
    .cout(cout_30[10]),
    .sum(sum_30[10]));
  AL_FADD comp30_11 (
    .a(i30[11]),
    .b(sum_29[11]),
    .c(cout_30[10]),
    .cout(cout_30[11]),
    .sum(sum_30[11]));
  AL_FADD comp30_12 (
    .a(i30[12]),
    .b(sum_29[12]),
    .c(cout_30[11]),
    .cout(cout_30[12]),
    .sum(sum_30[12]));
  AL_FADD comp30_13 (
    .a(i30[13]),
    .b(sum_29[13]),
    .c(cout_30[12]),
    .cout(cout_30[13]),
    .sum(sum_30[13]));
  AL_FADD comp30_14 (
    .a(i30[14]),
    .b(sum_29[14]),
    .c(cout_30[13]),
    .cout(cout_30[14]),
    .sum(sum_30[14]));
  AL_FADD comp30_15 (
    .a(i30[15]),
    .b(sum_29[15]),
    .c(cout_30[14]),
    .cout(cout_30[15]),
    .sum(sum_30[15]));
  AL_FADD comp30_16 (
    .a(i30[16]),
    .b(sum_29[16]),
    .c(cout_30[15]),
    .cout(cout_30[16]),
    .sum(sum_30[16]));
  AL_FADD comp30_17 (
    .a(i30[17]),
    .b(sum_29[17]),
    .c(cout_30[16]),
    .cout(cout_30[17]),
    .sum(sum_30[17]));
  AL_FADD comp30_18 (
    .a(i30[18]),
    .b(sum_29[18]),
    .c(cout_30[17]),
    .cout(cout_30[18]),
    .sum(sum_30[18]));
  AL_FADD comp30_19 (
    .a(i30[19]),
    .b(sum_29[19]),
    .c(cout_30[18]),
    .cout(cout_30[19]),
    .sum(sum_30[19]));
  AL_FADD comp30_2 (
    .a(i30[2]),
    .b(sum_29[2]),
    .c(cout_30[1]),
    .cout(cout_30[2]),
    .sum(sum_30[2]));
  AL_FADD comp30_20 (
    .a(i30[20]),
    .b(sum_29[20]),
    .c(cout_30[19]),
    .cout(cout_30[20]),
    .sum(sum_30[20]));
  AL_FADD comp30_21 (
    .a(i30[21]),
    .b(sum_29[21]),
    .c(cout_30[20]),
    .cout(cout_30[21]),
    .sum(sum_30[21]));
  AL_FADD comp30_22 (
    .a(i30[22]),
    .b(sum_29[22]),
    .c(cout_30[21]),
    .cout(cout_30[22]),
    .sum(sum_30[22]));
  AL_FADD comp30_23 (
    .a(i30[23]),
    .b(sum_29[23]),
    .c(cout_30[22]),
    .cout(cout_30[23]),
    .sum(sum_30[23]));
  AL_FADD comp30_24 (
    .a(i30[24]),
    .b(sum_29[24]),
    .c(cout_30[23]),
    .cout(cout_30[24]),
    .sum(sum_30[24]));
  AL_FADD comp30_25 (
    .a(i30[25]),
    .b(sum_29[25]),
    .c(cout_30[24]),
    .cout(cout_30[25]),
    .sum(sum_30[25]));
  AL_FADD comp30_26 (
    .a(i30[26]),
    .b(sum_29[26]),
    .c(cout_30[25]),
    .cout(cout_30[26]),
    .sum(sum_30[26]));
  AL_FADD comp30_27 (
    .a(i30[27]),
    .b(sum_29[27]),
    .c(cout_30[26]),
    .cout(cout_30[27]),
    .sum(sum_30[27]));
  AL_FADD comp30_28 (
    .a(i30[28]),
    .b(sum_29[28]),
    .c(cout_30[27]),
    .cout(cout_30[28]),
    .sum(sum_30[28]));
  AL_FADD comp30_29 (
    .a(i30[29]),
    .b(sum_29[29]),
    .c(cout_30[28]),
    .cout(cout_30[29]),
    .sum(sum_30[29]));
  AL_FADD comp30_3 (
    .a(i30[3]),
    .b(sum_29[3]),
    .c(cout_30[2]),
    .cout(cout_30[3]),
    .sum(sum_30[3]));
  AL_FADD comp30_30 (
    .a(i30[30]),
    .b(sum_29[30]),
    .c(cout_30[29]),
    .cout(cout_30[30]),
    .sum(sum_30[30]));
  AL_FADD comp30_31 (
    .a(i30[31]),
    .b(sum_29[31]),
    .c(cout_30[30]),
    .cout(cout_30[31]),
    .sum(sum_30[31]));
  AL_FADD comp30_32 (
    .a(1'b0),
    .b(sum_29[32]),
    .c(cout_30[31]),
    .cout(cout_30[32]),
    .sum(sum_30[32]));
  AL_FADD comp30_33 (
    .a(1'b0),
    .b(sum_29[33]),
    .c(cout_30[32]),
    .cout(cout_30[33]),
    .sum(sum_30[33]));
  AL_FADD comp30_34 (
    .a(1'b0),
    .b(sum_29[34]),
    .c(cout_30[33]),
    .cout(cout_30[34]),
    .sum(sum_30[34]));
  AL_FADD comp30_35 (
    .a(1'b0),
    .b(sum_29[35]),
    .c(cout_30[34]),
    .cout(cout_30[35]),
    .sum(sum_30[35]));
  AL_FADD comp30_36 (
    .a(1'b0),
    .b(sum_29[36]),
    .c(cout_30[35]),
    .cout(cout_30[36]),
    .sum(sum_30[36]));
  AL_FADD comp30_37 (
    .a(1'b0),
    .b(sum_29[37]),
    .c(cout_30[36]),
    .cout(cout_30[37]),
    .sum(sum_30[37]));
  AL_FADD comp30_38 (
    .a(1'b0),
    .b(sum_29[38]),
    .c(cout_30[37]),
    .cout(cout_30[38]),
    .sum(sum_30[38]));
  AL_FADD comp30_39 (
    .a(1'b0),
    .b(sum_29[39]),
    .c(cout_30[38]),
    .cout(cout_30[39]),
    .sum(sum_30[39]));
  AL_FADD comp30_4 (
    .a(i30[4]),
    .b(sum_29[4]),
    .c(cout_30[3]),
    .cout(cout_30[4]),
    .sum(sum_30[4]));
  AL_FADD comp30_40 (
    .a(1'b0),
    .b(sum_29[40]),
    .c(cout_30[39]),
    .cout(cout_30[40]),
    .sum(sum_30[40]));
  AL_FADD comp30_41 (
    .a(1'b0),
    .b(sum_29[41]),
    .c(cout_30[40]),
    .cout(cout_30[41]),
    .sum(sum_30[41]));
  AL_FADD comp30_42 (
    .a(1'b0),
    .b(sum_29[42]),
    .c(cout_30[41]),
    .cout(cout_30[42]),
    .sum(sum_30[42]));
  AL_FADD comp30_43 (
    .a(1'b0),
    .b(sum_29[43]),
    .c(cout_30[42]),
    .cout(cout_30[43]),
    .sum(sum_30[43]));
  AL_FADD comp30_44 (
    .a(1'b0),
    .b(sum_29[44]),
    .c(cout_30[43]),
    .cout(cout_30[44]),
    .sum(sum_30[44]));
  AL_FADD comp30_45 (
    .a(1'b0),
    .b(sum_29[45]),
    .c(cout_30[44]),
    .cout(cout_30[45]),
    .sum(sum_30[45]));
  AL_FADD comp30_46 (
    .a(1'b0),
    .b(sum_29[46]),
    .c(cout_30[45]),
    .cout(cout_30[46]),
    .sum(sum_30[46]));
  AL_FADD comp30_47 (
    .a(1'b0),
    .b(sum_29[47]),
    .c(cout_30[46]),
    .cout(cout_30[47]),
    .sum(sum_30[47]));
  AL_FADD comp30_48 (
    .a(1'b0),
    .b(sum_29[48]),
    .c(cout_30[47]),
    .cout(cout_30[48]),
    .sum(sum_30[48]));
  AL_FADD comp30_49 (
    .a(1'b0),
    .b(sum_29[49]),
    .c(cout_30[48]),
    .cout(cout_30[49]),
    .sum(sum_30[49]));
  AL_FADD comp30_5 (
    .a(i30[5]),
    .b(sum_29[5]),
    .c(cout_30[4]),
    .cout(cout_30[5]),
    .sum(sum_30[5]));
  AL_FADD comp30_50 (
    .a(1'b0),
    .b(sum_29[50]),
    .c(cout_30[49]),
    .cout(cout_30[50]),
    .sum(sum_30[50]));
  AL_FADD comp30_51 (
    .a(1'b0),
    .b(sum_29[51]),
    .c(cout_30[50]),
    .cout(cout_30[51]),
    .sum(sum_30[51]));
  AL_FADD comp30_52 (
    .a(1'b0),
    .b(sum_29[52]),
    .c(cout_30[51]),
    .cout(cout_30[52]),
    .sum(sum_30[52]));
  AL_FADD comp30_53 (
    .a(1'b0),
    .b(sum_29[53]),
    .c(cout_30[52]),
    .cout(cout_30[53]),
    .sum(sum_30[53]));
  AL_FADD comp30_54 (
    .a(1'b0),
    .b(sum_29[54]),
    .c(cout_30[53]),
    .cout(cout_30[54]),
    .sum(sum_30[54]));
  AL_FADD comp30_55 (
    .a(1'b0),
    .b(sum_29[55]),
    .c(cout_30[54]),
    .cout(cout_30[55]),
    .sum(sum_30[55]));
  AL_FADD comp30_56 (
    .a(1'b0),
    .b(sum_29[56]),
    .c(cout_30[55]),
    .cout(cout_30[56]),
    .sum(sum_30[56]));
  AL_FADD comp30_57 (
    .a(1'b0),
    .b(sum_29[57]),
    .c(cout_30[56]),
    .cout(cout_30[57]),
    .sum(sum_30[57]));
  AL_FADD comp30_58 (
    .a(1'b0),
    .b(sum_29[58]),
    .c(cout_30[57]),
    .cout(cout_30[58]),
    .sum(sum_30[58]));
  AL_FADD comp30_59 (
    .a(1'b0),
    .b(sum_29[59]),
    .c(cout_30[58]),
    .cout(cout_30[59]),
    .sum(sum_30[59]));
  AL_FADD comp30_6 (
    .a(i30[6]),
    .b(sum_29[6]),
    .c(cout_30[5]),
    .cout(cout_30[6]),
    .sum(sum_30[6]));
  AL_FADD comp30_60 (
    .a(1'b0),
    .b(sum_29[60]),
    .c(cout_30[59]),
    .cout(cout_30[60]),
    .sum(sum_30[60]));
  AL_FADD comp30_61 (
    .a(1'b0),
    .b(sum_29[61]),
    .c(cout_30[60]),
    .cout(cout_30[61]),
    .sum(sum_30[61]));
  AL_FADD comp30_62 (
    .a(1'b0),
    .b(sum_29[62]),
    .c(cout_30[61]),
    .cout(cout_30[62]),
    .sum(sum_30[62]));
  AL_FADD comp30_63 (
    .a(1'b0),
    .b(sum_29[63]),
    .c(cout_30[62]),
    .cout(cout_30[63]),
    .sum(sum_30[63]));
  AL_FADD comp30_7 (
    .a(i30[7]),
    .b(sum_29[7]),
    .c(cout_30[6]),
    .cout(cout_30[7]),
    .sum(sum_30[7]));
  AL_FADD comp30_8 (
    .a(i30[8]),
    .b(sum_29[8]),
    .c(cout_30[7]),
    .cout(cout_30[8]),
    .sum(sum_30[8]));
  AL_FADD comp30_9 (
    .a(i30[9]),
    .b(sum_29[9]),
    .c(cout_30[8]),
    .cout(cout_30[9]),
    .sum(sum_30[9]));
  AL_FADD comp31_0 (
    .a(sum_30[0]),
    .b(net_nb31_0),
    .c(1'b1),
    .cout(cout_31[0]),
    .sum(sum_31[0]));
  AL_FADD comp31_1 (
    .a(sum_30[1]),
    .b(net_nb31_1),
    .c(cout_31[0]),
    .cout(cout_31[1]),
    .sum(sum_31[1]));
  AL_FADD comp31_10 (
    .a(sum_30[10]),
    .b(net_nb31_10),
    .c(cout_31[9]),
    .cout(cout_31[10]),
    .sum(sum_31[10]));
  AL_FADD comp31_11 (
    .a(sum_30[11]),
    .b(net_nb31_11),
    .c(cout_31[10]),
    .cout(cout_31[11]),
    .sum(sum_31[11]));
  AL_FADD comp31_12 (
    .a(sum_30[12]),
    .b(net_nb31_12),
    .c(cout_31[11]),
    .cout(cout_31[12]),
    .sum(sum_31[12]));
  AL_FADD comp31_13 (
    .a(sum_30[13]),
    .b(net_nb31_13),
    .c(cout_31[12]),
    .cout(cout_31[13]),
    .sum(sum_31[13]));
  AL_FADD comp31_14 (
    .a(sum_30[14]),
    .b(net_nb31_14),
    .c(cout_31[13]),
    .cout(cout_31[14]),
    .sum(sum_31[14]));
  AL_FADD comp31_15 (
    .a(sum_30[15]),
    .b(net_nb31_15),
    .c(cout_31[14]),
    .cout(cout_31[15]),
    .sum(sum_31[15]));
  AL_FADD comp31_16 (
    .a(sum_30[16]),
    .b(net_nb31_16),
    .c(cout_31[15]),
    .cout(cout_31[16]),
    .sum(sum_31[16]));
  AL_FADD comp31_17 (
    .a(sum_30[17]),
    .b(net_nb31_17),
    .c(cout_31[16]),
    .cout(cout_31[17]),
    .sum(sum_31[17]));
  AL_FADD comp31_18 (
    .a(sum_30[18]),
    .b(net_nb31_18),
    .c(cout_31[17]),
    .cout(cout_31[18]),
    .sum(sum_31[18]));
  AL_FADD comp31_19 (
    .a(sum_30[19]),
    .b(net_nb31_19),
    .c(cout_31[18]),
    .cout(cout_31[19]),
    .sum(sum_31[19]));
  AL_FADD comp31_2 (
    .a(sum_30[2]),
    .b(net_nb31_2),
    .c(cout_31[1]),
    .cout(cout_31[2]),
    .sum(sum_31[2]));
  AL_FADD comp31_20 (
    .a(sum_30[20]),
    .b(net_nb31_20),
    .c(cout_31[19]),
    .cout(cout_31[20]),
    .sum(sum_31[20]));
  AL_FADD comp31_21 (
    .a(sum_30[21]),
    .b(net_nb31_21),
    .c(cout_31[20]),
    .cout(cout_31[21]),
    .sum(sum_31[21]));
  AL_FADD comp31_22 (
    .a(sum_30[22]),
    .b(net_nb31_22),
    .c(cout_31[21]),
    .cout(cout_31[22]),
    .sum(sum_31[22]));
  AL_FADD comp31_23 (
    .a(sum_30[23]),
    .b(net_nb31_23),
    .c(cout_31[22]),
    .cout(cout_31[23]),
    .sum(sum_31[23]));
  AL_FADD comp31_24 (
    .a(sum_30[24]),
    .b(net_nb31_24),
    .c(cout_31[23]),
    .cout(cout_31[24]),
    .sum(sum_31[24]));
  AL_FADD comp31_25 (
    .a(sum_30[25]),
    .b(net_nb31_25),
    .c(cout_31[24]),
    .cout(cout_31[25]),
    .sum(sum_31[25]));
  AL_FADD comp31_26 (
    .a(sum_30[26]),
    .b(net_nb31_26),
    .c(cout_31[25]),
    .cout(cout_31[26]),
    .sum(sum_31[26]));
  AL_FADD comp31_27 (
    .a(sum_30[27]),
    .b(net_nb31_27),
    .c(cout_31[26]),
    .cout(cout_31[27]),
    .sum(sum_31[27]));
  AL_FADD comp31_28 (
    .a(sum_30[28]),
    .b(net_nb31_28),
    .c(cout_31[27]),
    .cout(cout_31[28]),
    .sum(sum_31[28]));
  AL_FADD comp31_29 (
    .a(sum_30[29]),
    .b(net_nb31_29),
    .c(cout_31[28]),
    .cout(cout_31[29]),
    .sum(sum_31[29]));
  AL_FADD comp31_3 (
    .a(sum_30[3]),
    .b(net_nb31_3),
    .c(cout_31[2]),
    .cout(cout_31[3]),
    .sum(sum_31[3]));
  AL_FADD comp31_30 (
    .a(sum_30[30]),
    .b(net_nb31_30),
    .c(cout_31[29]),
    .cout(cout_31[30]),
    .sum(sum_31[30]));
  AL_FADD comp31_31 (
    .a(sum_30[31]),
    .b(net_nb31_31),
    .c(cout_31[30]),
    .cout(cout_31[31]),
    .sum(sum_31[31]));
  AL_FADD comp31_32 (
    .a(sum_30[32]),
    .b(net_nb31_32),
    .c(cout_31[31]),
    .cout(cout_31[32]),
    .sum(sum_31[32]));
  AL_FADD comp31_33 (
    .a(sum_30[33]),
    .b(net_nb31_33),
    .c(cout_31[32]),
    .cout(cout_31[33]),
    .sum(sum_31[33]));
  AL_FADD comp31_34 (
    .a(sum_30[34]),
    .b(net_nb31_34),
    .c(cout_31[33]),
    .cout(cout_31[34]),
    .sum(sum_31[34]));
  AL_FADD comp31_35 (
    .a(sum_30[35]),
    .b(net_nb31_35),
    .c(cout_31[34]),
    .cout(cout_31[35]),
    .sum(sum_31[35]));
  AL_FADD comp31_36 (
    .a(sum_30[36]),
    .b(net_nb31_36),
    .c(cout_31[35]),
    .cout(cout_31[36]),
    .sum(sum_31[36]));
  AL_FADD comp31_37 (
    .a(sum_30[37]),
    .b(net_nb31_37),
    .c(cout_31[36]),
    .cout(cout_31[37]),
    .sum(sum_31[37]));
  AL_FADD comp31_38 (
    .a(sum_30[38]),
    .b(net_nb31_38),
    .c(cout_31[37]),
    .cout(cout_31[38]),
    .sum(sum_31[38]));
  AL_FADD comp31_39 (
    .a(sum_30[39]),
    .b(net_nb31_39),
    .c(cout_31[38]),
    .cout(cout_31[39]),
    .sum(sum_31[39]));
  AL_FADD comp31_4 (
    .a(sum_30[4]),
    .b(net_nb31_4),
    .c(cout_31[3]),
    .cout(cout_31[4]),
    .sum(sum_31[4]));
  AL_FADD comp31_40 (
    .a(sum_30[40]),
    .b(net_nb31_40),
    .c(cout_31[39]),
    .cout(cout_31[40]),
    .sum(sum_31[40]));
  AL_FADD comp31_41 (
    .a(sum_30[41]),
    .b(net_nb31_41),
    .c(cout_31[40]),
    .cout(cout_31[41]),
    .sum(sum_31[41]));
  AL_FADD comp31_42 (
    .a(sum_30[42]),
    .b(net_nb31_42),
    .c(cout_31[41]),
    .cout(cout_31[42]),
    .sum(sum_31[42]));
  AL_FADD comp31_43 (
    .a(sum_30[43]),
    .b(net_nb31_43),
    .c(cout_31[42]),
    .cout(cout_31[43]),
    .sum(sum_31[43]));
  AL_FADD comp31_44 (
    .a(sum_30[44]),
    .b(net_nb31_44),
    .c(cout_31[43]),
    .cout(cout_31[44]),
    .sum(sum_31[44]));
  AL_FADD comp31_45 (
    .a(sum_30[45]),
    .b(net_nb31_45),
    .c(cout_31[44]),
    .cout(cout_31[45]),
    .sum(sum_31[45]));
  AL_FADD comp31_46 (
    .a(sum_30[46]),
    .b(net_nb31_46),
    .c(cout_31[45]),
    .cout(cout_31[46]),
    .sum(sum_31[46]));
  AL_FADD comp31_47 (
    .a(sum_30[47]),
    .b(net_nb31_47),
    .c(cout_31[46]),
    .cout(cout_31[47]),
    .sum(sum_31[47]));
  AL_FADD comp31_48 (
    .a(sum_30[48]),
    .b(net_nb31_48),
    .c(cout_31[47]),
    .cout(cout_31[48]),
    .sum(sum_31[48]));
  AL_FADD comp31_49 (
    .a(sum_30[49]),
    .b(net_nb31_49),
    .c(cout_31[48]),
    .cout(cout_31[49]),
    .sum(sum_31[49]));
  AL_FADD comp31_5 (
    .a(sum_30[5]),
    .b(net_nb31_5),
    .c(cout_31[4]),
    .cout(cout_31[5]),
    .sum(sum_31[5]));
  AL_FADD comp31_50 (
    .a(sum_30[50]),
    .b(net_nb31_50),
    .c(cout_31[49]),
    .cout(cout_31[50]),
    .sum(sum_31[50]));
  AL_FADD comp31_51 (
    .a(sum_30[51]),
    .b(net_nb31_51),
    .c(cout_31[50]),
    .cout(cout_31[51]),
    .sum(sum_31[51]));
  AL_FADD comp31_52 (
    .a(sum_30[52]),
    .b(net_nb31_52),
    .c(cout_31[51]),
    .cout(cout_31[52]),
    .sum(sum_31[52]));
  AL_FADD comp31_53 (
    .a(sum_30[53]),
    .b(net_nb31_53),
    .c(cout_31[52]),
    .cout(cout_31[53]),
    .sum(sum_31[53]));
  AL_FADD comp31_54 (
    .a(sum_30[54]),
    .b(net_nb31_54),
    .c(cout_31[53]),
    .cout(cout_31[54]),
    .sum(sum_31[54]));
  AL_FADD comp31_55 (
    .a(sum_30[55]),
    .b(net_nb31_55),
    .c(cout_31[54]),
    .cout(cout_31[55]),
    .sum(sum_31[55]));
  AL_FADD comp31_56 (
    .a(sum_30[56]),
    .b(net_nb31_56),
    .c(cout_31[55]),
    .cout(cout_31[56]),
    .sum(sum_31[56]));
  AL_FADD comp31_57 (
    .a(sum_30[57]),
    .b(net_nb31_57),
    .c(cout_31[56]),
    .cout(cout_31[57]),
    .sum(sum_31[57]));
  AL_FADD comp31_58 (
    .a(sum_30[58]),
    .b(net_nb31_58),
    .c(cout_31[57]),
    .cout(cout_31[58]),
    .sum(sum_31[58]));
  AL_FADD comp31_59 (
    .a(sum_30[59]),
    .b(net_nb31_59),
    .c(cout_31[58]),
    .cout(cout_31[59]),
    .sum(sum_31[59]));
  AL_FADD comp31_6 (
    .a(sum_30[6]),
    .b(net_nb31_6),
    .c(cout_31[5]),
    .cout(cout_31[6]),
    .sum(sum_31[6]));
  AL_FADD comp31_60 (
    .a(sum_30[60]),
    .b(net_nb31_60),
    .c(cout_31[59]),
    .cout(cout_31[60]),
    .sum(sum_31[60]));
  AL_FADD comp31_61 (
    .a(sum_30[61]),
    .b(net_nb31_61),
    .c(cout_31[60]),
    .cout(cout_31[61]),
    .sum(sum_31[61]));
  AL_FADD comp31_62 (
    .a(sum_30[62]),
    .b(net_nb31_62),
    .c(cout_31[61]),
    .cout(cout_31[62]),
    .sum(sum_31[62]));
  AL_FADD comp31_63 (
    .a(sum_30[63]),
    .b(net_nb31_63),
    .c(cout_31[62]),
    .cout(cout_31[63]),
    .sum(sum_31[63]));
  AL_FADD comp31_7 (
    .a(sum_30[7]),
    .b(net_nb31_7),
    .c(cout_31[6]),
    .cout(cout_31[7]),
    .sum(sum_31[7]));
  AL_FADD comp31_8 (
    .a(sum_30[8]),
    .b(net_nb31_8),
    .c(cout_31[7]),
    .cout(cout_31[8]),
    .sum(sum_31[8]));
  AL_FADD comp31_9 (
    .a(sum_30[9]),
    .b(net_nb31_9),
    .c(cout_31[8]),
    .cout(cout_31[9]),
    .sum(sum_31[9]));
  AL_FADD comp32_0 (
    .a(sum_31[0]),
    .b(net_nb32_0),
    .c(1'b1),
    .cout(cout_32[0]),
    .sum(sum_32[0]));
  AL_FADD comp32_1 (
    .a(sum_31[1]),
    .b(net_nb32_1),
    .c(cout_32[0]),
    .cout(cout_32[1]),
    .sum(sum_32[1]));
  AL_FADD comp32_10 (
    .a(sum_31[10]),
    .b(net_nb32_10),
    .c(cout_32[9]),
    .cout(cout_32[10]),
    .sum(sum_32[10]));
  AL_FADD comp32_11 (
    .a(sum_31[11]),
    .b(net_nb32_11),
    .c(cout_32[10]),
    .cout(cout_32[11]),
    .sum(sum_32[11]));
  AL_FADD comp32_12 (
    .a(sum_31[12]),
    .b(net_nb32_12),
    .c(cout_32[11]),
    .cout(cout_32[12]),
    .sum(sum_32[12]));
  AL_FADD comp32_13 (
    .a(sum_31[13]),
    .b(net_nb32_13),
    .c(cout_32[12]),
    .cout(cout_32[13]),
    .sum(sum_32[13]));
  AL_FADD comp32_14 (
    .a(sum_31[14]),
    .b(net_nb32_14),
    .c(cout_32[13]),
    .cout(cout_32[14]),
    .sum(sum_32[14]));
  AL_FADD comp32_15 (
    .a(sum_31[15]),
    .b(net_nb32_15),
    .c(cout_32[14]),
    .cout(cout_32[15]),
    .sum(sum_32[15]));
  AL_FADD comp32_16 (
    .a(sum_31[16]),
    .b(net_nb32_16),
    .c(cout_32[15]),
    .cout(cout_32[16]),
    .sum(sum_32[16]));
  AL_FADD comp32_17 (
    .a(sum_31[17]),
    .b(net_nb32_17),
    .c(cout_32[16]),
    .cout(cout_32[17]),
    .sum(sum_32[17]));
  AL_FADD comp32_18 (
    .a(sum_31[18]),
    .b(net_nb32_18),
    .c(cout_32[17]),
    .cout(cout_32[18]),
    .sum(sum_32[18]));
  AL_FADD comp32_19 (
    .a(sum_31[19]),
    .b(net_nb32_19),
    .c(cout_32[18]),
    .cout(cout_32[19]),
    .sum(sum_32[19]));
  AL_FADD comp32_2 (
    .a(sum_31[2]),
    .b(net_nb32_2),
    .c(cout_32[1]),
    .cout(cout_32[2]),
    .sum(sum_32[2]));
  AL_FADD comp32_20 (
    .a(sum_31[20]),
    .b(net_nb32_20),
    .c(cout_32[19]),
    .cout(cout_32[20]),
    .sum(sum_32[20]));
  AL_FADD comp32_21 (
    .a(sum_31[21]),
    .b(net_nb32_21),
    .c(cout_32[20]),
    .cout(cout_32[21]),
    .sum(sum_32[21]));
  AL_FADD comp32_22 (
    .a(sum_31[22]),
    .b(net_nb32_22),
    .c(cout_32[21]),
    .cout(cout_32[22]),
    .sum(sum_32[22]));
  AL_FADD comp32_23 (
    .a(sum_31[23]),
    .b(net_nb32_23),
    .c(cout_32[22]),
    .cout(cout_32[23]),
    .sum(sum_32[23]));
  AL_FADD comp32_24 (
    .a(sum_31[24]),
    .b(net_nb32_24),
    .c(cout_32[23]),
    .cout(cout_32[24]),
    .sum(sum_32[24]));
  AL_FADD comp32_25 (
    .a(sum_31[25]),
    .b(net_nb32_25),
    .c(cout_32[24]),
    .cout(cout_32[25]),
    .sum(sum_32[25]));
  AL_FADD comp32_26 (
    .a(sum_31[26]),
    .b(net_nb32_26),
    .c(cout_32[25]),
    .cout(cout_32[26]),
    .sum(sum_32[26]));
  AL_FADD comp32_27 (
    .a(sum_31[27]),
    .b(net_nb32_27),
    .c(cout_32[26]),
    .cout(cout_32[27]),
    .sum(sum_32[27]));
  AL_FADD comp32_28 (
    .a(sum_31[28]),
    .b(net_nb32_28),
    .c(cout_32[27]),
    .cout(cout_32[28]),
    .sum(sum_32[28]));
  AL_FADD comp32_29 (
    .a(sum_31[29]),
    .b(net_nb32_29),
    .c(cout_32[28]),
    .cout(cout_32[29]),
    .sum(sum_32[29]));
  AL_FADD comp32_3 (
    .a(sum_31[3]),
    .b(net_nb32_3),
    .c(cout_32[2]),
    .cout(cout_32[3]),
    .sum(sum_32[3]));
  AL_FADD comp32_30 (
    .a(sum_31[30]),
    .b(net_nb32_30),
    .c(cout_32[29]),
    .cout(cout_32[30]),
    .sum(sum_32[30]));
  AL_FADD comp32_31 (
    .a(sum_31[31]),
    .b(net_nb32_31),
    .c(cout_32[30]),
    .cout(cout_32[31]),
    .sum(sum_32[31]));
  AL_FADD comp32_32 (
    .a(sum_31[32]),
    .b(net_nb32_32),
    .c(cout_32[31]),
    .cout(cout_32[32]),
    .sum(sum_32[32]));
  AL_FADD comp32_33 (
    .a(sum_31[33]),
    .b(net_nb32_33),
    .c(cout_32[32]),
    .cout(cout_32[33]),
    .sum(sum_32[33]));
  AL_FADD comp32_34 (
    .a(sum_31[34]),
    .b(net_nb32_34),
    .c(cout_32[33]),
    .cout(cout_32[34]),
    .sum(sum_32[34]));
  AL_FADD comp32_35 (
    .a(sum_31[35]),
    .b(net_nb32_35),
    .c(cout_32[34]),
    .cout(cout_32[35]),
    .sum(sum_32[35]));
  AL_FADD comp32_36 (
    .a(sum_31[36]),
    .b(net_nb32_36),
    .c(cout_32[35]),
    .cout(cout_32[36]),
    .sum(sum_32[36]));
  AL_FADD comp32_37 (
    .a(sum_31[37]),
    .b(net_nb32_37),
    .c(cout_32[36]),
    .cout(cout_32[37]),
    .sum(sum_32[37]));
  AL_FADD comp32_38 (
    .a(sum_31[38]),
    .b(net_nb32_38),
    .c(cout_32[37]),
    .cout(cout_32[38]),
    .sum(sum_32[38]));
  AL_FADD comp32_39 (
    .a(sum_31[39]),
    .b(net_nb32_39),
    .c(cout_32[38]),
    .cout(cout_32[39]),
    .sum(sum_32[39]));
  AL_FADD comp32_4 (
    .a(sum_31[4]),
    .b(net_nb32_4),
    .c(cout_32[3]),
    .cout(cout_32[4]),
    .sum(sum_32[4]));
  AL_FADD comp32_40 (
    .a(sum_31[40]),
    .b(net_nb32_40),
    .c(cout_32[39]),
    .cout(cout_32[40]),
    .sum(sum_32[40]));
  AL_FADD comp32_41 (
    .a(sum_31[41]),
    .b(net_nb32_41),
    .c(cout_32[40]),
    .cout(cout_32[41]),
    .sum(sum_32[41]));
  AL_FADD comp32_42 (
    .a(sum_31[42]),
    .b(net_nb32_42),
    .c(cout_32[41]),
    .cout(cout_32[42]),
    .sum(sum_32[42]));
  AL_FADD comp32_43 (
    .a(sum_31[43]),
    .b(net_nb32_43),
    .c(cout_32[42]),
    .cout(cout_32[43]),
    .sum(sum_32[43]));
  AL_FADD comp32_44 (
    .a(sum_31[44]),
    .b(net_nb32_44),
    .c(cout_32[43]),
    .cout(cout_32[44]),
    .sum(sum_32[44]));
  AL_FADD comp32_45 (
    .a(sum_31[45]),
    .b(net_nb32_45),
    .c(cout_32[44]),
    .cout(cout_32[45]),
    .sum(sum_32[45]));
  AL_FADD comp32_46 (
    .a(sum_31[46]),
    .b(net_nb32_46),
    .c(cout_32[45]),
    .cout(cout_32[46]),
    .sum(sum_32[46]));
  AL_FADD comp32_47 (
    .a(sum_31[47]),
    .b(net_nb32_47),
    .c(cout_32[46]),
    .cout(cout_32[47]),
    .sum(sum_32[47]));
  AL_FADD comp32_48 (
    .a(sum_31[48]),
    .b(net_nb32_48),
    .c(cout_32[47]),
    .cout(cout_32[48]),
    .sum(sum_32[48]));
  AL_FADD comp32_49 (
    .a(sum_31[49]),
    .b(net_nb32_49),
    .c(cout_32[48]),
    .cout(cout_32[49]),
    .sum(sum_32[49]));
  AL_FADD comp32_5 (
    .a(sum_31[5]),
    .b(net_nb32_5),
    .c(cout_32[4]),
    .cout(cout_32[5]),
    .sum(sum_32[5]));
  AL_FADD comp32_50 (
    .a(sum_31[50]),
    .b(net_nb32_50),
    .c(cout_32[49]),
    .cout(cout_32[50]),
    .sum(sum_32[50]));
  AL_FADD comp32_51 (
    .a(sum_31[51]),
    .b(net_nb32_51),
    .c(cout_32[50]),
    .cout(cout_32[51]),
    .sum(sum_32[51]));
  AL_FADD comp32_52 (
    .a(sum_31[52]),
    .b(net_nb32_52),
    .c(cout_32[51]),
    .cout(cout_32[52]),
    .sum(sum_32[52]));
  AL_FADD comp32_53 (
    .a(sum_31[53]),
    .b(net_nb32_53),
    .c(cout_32[52]),
    .cout(cout_32[53]),
    .sum(sum_32[53]));
  AL_FADD comp32_54 (
    .a(sum_31[54]),
    .b(net_nb32_54),
    .c(cout_32[53]),
    .cout(cout_32[54]),
    .sum(sum_32[54]));
  AL_FADD comp32_55 (
    .a(sum_31[55]),
    .b(net_nb32_55),
    .c(cout_32[54]),
    .cout(cout_32[55]),
    .sum(sum_32[55]));
  AL_FADD comp32_56 (
    .a(sum_31[56]),
    .b(net_nb32_56),
    .c(cout_32[55]),
    .cout(cout_32[56]),
    .sum(sum_32[56]));
  AL_FADD comp32_57 (
    .a(sum_31[57]),
    .b(net_nb32_57),
    .c(cout_32[56]),
    .cout(cout_32[57]),
    .sum(sum_32[57]));
  AL_FADD comp32_58 (
    .a(sum_31[58]),
    .b(net_nb32_58),
    .c(cout_32[57]),
    .cout(cout_32[58]),
    .sum(sum_32[58]));
  AL_FADD comp32_59 (
    .a(sum_31[59]),
    .b(net_nb32_59),
    .c(cout_32[58]),
    .cout(cout_32[59]),
    .sum(sum_32[59]));
  AL_FADD comp32_6 (
    .a(sum_31[6]),
    .b(net_nb32_6),
    .c(cout_32[5]),
    .cout(cout_32[6]),
    .sum(sum_32[6]));
  AL_FADD comp32_60 (
    .a(sum_31[60]),
    .b(net_nb32_60),
    .c(cout_32[59]),
    .cout(cout_32[60]),
    .sum(sum_32[60]));
  AL_FADD comp32_61 (
    .a(sum_31[61]),
    .b(net_nb32_61),
    .c(cout_32[60]),
    .cout(cout_32[61]),
    .sum(sum_32[61]));
  AL_FADD comp32_62 (
    .a(sum_31[62]),
    .b(net_nb32_62),
    .c(cout_32[61]),
    .cout(cout_32[62]),
    .sum(sum_32[62]));
  AL_FADD comp32_63 (
    .a(sum_31[63]),
    .b(net_nb32_63),
    .c(cout_32[62]),
    .cout(cout_32[63]),
    .sum(sum_32[63]));
  AL_FADD comp32_7 (
    .a(sum_31[7]),
    .b(net_nb32_7),
    .c(cout_32[6]),
    .cout(cout_32[7]),
    .sum(sum_32[7]));
  AL_FADD comp32_8 (
    .a(sum_31[8]),
    .b(net_nb32_8),
    .c(cout_32[7]),
    .cout(cout_32[8]),
    .sum(sum_32[8]));
  AL_FADD comp32_9 (
    .a(sum_31[9]),
    .b(net_nb32_9),
    .c(cout_32[8]),
    .cout(cout_32[9]),
    .sum(sum_32[9]));
  AL_FADD comp3_0 (
    .a(i3[0]),
    .b(sum_2[0]),
    .c(1'b0),
    .cout(cout_3[0]),
    .sum(sum_3[0]));
  AL_FADD comp3_1 (
    .a(i3[1]),
    .b(sum_2[1]),
    .c(cout_3[0]),
    .cout(cout_3[1]),
    .sum(sum_3[1]));
  AL_FADD comp3_10 (
    .a(i3[10]),
    .b(sum_2[10]),
    .c(cout_3[9]),
    .cout(cout_3[10]),
    .sum(sum_3[10]));
  AL_FADD comp3_11 (
    .a(i3[11]),
    .b(sum_2[11]),
    .c(cout_3[10]),
    .cout(cout_3[11]),
    .sum(sum_3[11]));
  AL_FADD comp3_12 (
    .a(i3[12]),
    .b(sum_2[12]),
    .c(cout_3[11]),
    .cout(cout_3[12]),
    .sum(sum_3[12]));
  AL_FADD comp3_13 (
    .a(i3[13]),
    .b(sum_2[13]),
    .c(cout_3[12]),
    .cout(cout_3[13]),
    .sum(sum_3[13]));
  AL_FADD comp3_14 (
    .a(i3[14]),
    .b(sum_2[14]),
    .c(cout_3[13]),
    .cout(cout_3[14]),
    .sum(sum_3[14]));
  AL_FADD comp3_15 (
    .a(i3[15]),
    .b(sum_2[15]),
    .c(cout_3[14]),
    .cout(cout_3[15]),
    .sum(sum_3[15]));
  AL_FADD comp3_16 (
    .a(i3[16]),
    .b(sum_2[16]),
    .c(cout_3[15]),
    .cout(cout_3[16]),
    .sum(sum_3[16]));
  AL_FADD comp3_17 (
    .a(i3[17]),
    .b(sum_2[17]),
    .c(cout_3[16]),
    .cout(cout_3[17]),
    .sum(sum_3[17]));
  AL_FADD comp3_18 (
    .a(i3[18]),
    .b(sum_2[18]),
    .c(cout_3[17]),
    .cout(cout_3[18]),
    .sum(sum_3[18]));
  AL_FADD comp3_19 (
    .a(i3[19]),
    .b(sum_2[19]),
    .c(cout_3[18]),
    .cout(cout_3[19]),
    .sum(sum_3[19]));
  AL_FADD comp3_2 (
    .a(i3[2]),
    .b(sum_2[2]),
    .c(cout_3[1]),
    .cout(cout_3[2]),
    .sum(sum_3[2]));
  AL_FADD comp3_20 (
    .a(i3[20]),
    .b(sum_2[20]),
    .c(cout_3[19]),
    .cout(cout_3[20]),
    .sum(sum_3[20]));
  AL_FADD comp3_21 (
    .a(i3[21]),
    .b(sum_2[21]),
    .c(cout_3[20]),
    .cout(cout_3[21]),
    .sum(sum_3[21]));
  AL_FADD comp3_22 (
    .a(i3[22]),
    .b(sum_2[22]),
    .c(cout_3[21]),
    .cout(cout_3[22]),
    .sum(sum_3[22]));
  AL_FADD comp3_23 (
    .a(i3[23]),
    .b(sum_2[23]),
    .c(cout_3[22]),
    .cout(cout_3[23]),
    .sum(sum_3[23]));
  AL_FADD comp3_24 (
    .a(i3[24]),
    .b(sum_2[24]),
    .c(cout_3[23]),
    .cout(cout_3[24]),
    .sum(sum_3[24]));
  AL_FADD comp3_25 (
    .a(i3[25]),
    .b(sum_2[25]),
    .c(cout_3[24]),
    .cout(cout_3[25]),
    .sum(sum_3[25]));
  AL_FADD comp3_26 (
    .a(i3[26]),
    .b(sum_2[26]),
    .c(cout_3[25]),
    .cout(cout_3[26]),
    .sum(sum_3[26]));
  AL_FADD comp3_27 (
    .a(i3[27]),
    .b(sum_2[27]),
    .c(cout_3[26]),
    .cout(cout_3[27]),
    .sum(sum_3[27]));
  AL_FADD comp3_28 (
    .a(i3[28]),
    .b(sum_2[28]),
    .c(cout_3[27]),
    .cout(cout_3[28]),
    .sum(sum_3[28]));
  AL_FADD comp3_29 (
    .a(i3[29]),
    .b(sum_2[29]),
    .c(cout_3[28]),
    .cout(cout_3[29]),
    .sum(sum_3[29]));
  AL_FADD comp3_3 (
    .a(i3[3]),
    .b(sum_2[3]),
    .c(cout_3[2]),
    .cout(cout_3[3]),
    .sum(sum_3[3]));
  AL_FADD comp3_30 (
    .a(i3[30]),
    .b(sum_2[30]),
    .c(cout_3[29]),
    .cout(cout_3[30]),
    .sum(sum_3[30]));
  AL_FADD comp3_31 (
    .a(i3[31]),
    .b(sum_2[31]),
    .c(cout_3[30]),
    .cout(cout_3[31]),
    .sum(sum_3[31]));
  AL_FADD comp3_32 (
    .a(i3[32]),
    .b(sum_2[32]),
    .c(cout_3[31]),
    .cout(cout_3[32]),
    .sum(sum_3[32]));
  AL_FADD comp3_33 (
    .a(i3[33]),
    .b(sum_2[33]),
    .c(cout_3[32]),
    .cout(cout_3[33]),
    .sum(sum_3[33]));
  AL_FADD comp3_34 (
    .a(i3[34]),
    .b(sum_2[34]),
    .c(cout_3[33]),
    .cout(cout_3[34]),
    .sum(sum_3[34]));
  AL_FADD comp3_35 (
    .a(i3[35]),
    .b(sum_2[35]),
    .c(cout_3[34]),
    .cout(cout_3[35]),
    .sum(sum_3[35]));
  AL_FADD comp3_36 (
    .a(i3[36]),
    .b(sum_2[36]),
    .c(cout_3[35]),
    .cout(cout_3[36]),
    .sum(sum_3[36]));
  AL_FADD comp3_37 (
    .a(i3[37]),
    .b(sum_2[37]),
    .c(cout_3[36]),
    .cout(cout_3[37]),
    .sum(sum_3[37]));
  AL_FADD comp3_38 (
    .a(i3[38]),
    .b(sum_2[38]),
    .c(cout_3[37]),
    .cout(cout_3[38]),
    .sum(sum_3[38]));
  AL_FADD comp3_39 (
    .a(i3[39]),
    .b(sum_2[39]),
    .c(cout_3[38]),
    .cout(cout_3[39]),
    .sum(sum_3[39]));
  AL_FADD comp3_4 (
    .a(i3[4]),
    .b(sum_2[4]),
    .c(cout_3[3]),
    .cout(cout_3[4]),
    .sum(sum_3[4]));
  AL_FADD comp3_40 (
    .a(i3[40]),
    .b(sum_2[40]),
    .c(cout_3[39]),
    .cout(cout_3[40]),
    .sum(sum_3[40]));
  AL_FADD comp3_41 (
    .a(i3[41]),
    .b(sum_2[41]),
    .c(cout_3[40]),
    .cout(cout_3[41]),
    .sum(sum_3[41]));
  AL_FADD comp3_42 (
    .a(i3[42]),
    .b(sum_2[42]),
    .c(cout_3[41]),
    .cout(cout_3[42]),
    .sum(sum_3[42]));
  AL_FADD comp3_43 (
    .a(i3[43]),
    .b(sum_2[43]),
    .c(cout_3[42]),
    .cout(cout_3[43]),
    .sum(sum_3[43]));
  AL_FADD comp3_44 (
    .a(i3[44]),
    .b(sum_2[44]),
    .c(cout_3[43]),
    .cout(cout_3[44]),
    .sum(sum_3[44]));
  AL_FADD comp3_45 (
    .a(i3[45]),
    .b(sum_2[45]),
    .c(cout_3[44]),
    .cout(cout_3[45]),
    .sum(sum_3[45]));
  AL_FADD comp3_46 (
    .a(i3[46]),
    .b(sum_2[46]),
    .c(cout_3[45]),
    .cout(cout_3[46]),
    .sum(sum_3[46]));
  AL_FADD comp3_47 (
    .a(i3[47]),
    .b(sum_2[47]),
    .c(cout_3[46]),
    .cout(cout_3[47]),
    .sum(sum_3[47]));
  AL_FADD comp3_48 (
    .a(i3[48]),
    .b(sum_2[48]),
    .c(cout_3[47]),
    .cout(cout_3[48]),
    .sum(sum_3[48]));
  AL_FADD comp3_49 (
    .a(i3[49]),
    .b(sum_2[49]),
    .c(cout_3[48]),
    .cout(cout_3[49]),
    .sum(sum_3[49]));
  AL_FADD comp3_5 (
    .a(i3[5]),
    .b(sum_2[5]),
    .c(cout_3[4]),
    .cout(cout_3[5]),
    .sum(sum_3[5]));
  AL_FADD comp3_50 (
    .a(i3[50]),
    .b(sum_2[50]),
    .c(cout_3[49]),
    .cout(cout_3[50]),
    .sum(sum_3[50]));
  AL_FADD comp3_51 (
    .a(i3[51]),
    .b(sum_2[51]),
    .c(cout_3[50]),
    .cout(cout_3[51]),
    .sum(sum_3[51]));
  AL_FADD comp3_52 (
    .a(i3[52]),
    .b(sum_2[52]),
    .c(cout_3[51]),
    .cout(cout_3[52]),
    .sum(sum_3[52]));
  AL_FADD comp3_53 (
    .a(i3[53]),
    .b(sum_2[53]),
    .c(cout_3[52]),
    .cout(cout_3[53]),
    .sum(sum_3[53]));
  AL_FADD comp3_54 (
    .a(i3[54]),
    .b(sum_2[54]),
    .c(cout_3[53]),
    .cout(cout_3[54]),
    .sum(sum_3[54]));
  AL_FADD comp3_55 (
    .a(i3[55]),
    .b(sum_2[55]),
    .c(cout_3[54]),
    .cout(cout_3[55]),
    .sum(sum_3[55]));
  AL_FADD comp3_56 (
    .a(i3[56]),
    .b(sum_2[56]),
    .c(cout_3[55]),
    .cout(cout_3[56]),
    .sum(sum_3[56]));
  AL_FADD comp3_57 (
    .a(i3[57]),
    .b(sum_2[57]),
    .c(cout_3[56]),
    .cout(cout_3[57]),
    .sum(sum_3[57]));
  AL_FADD comp3_58 (
    .a(i3[58]),
    .b(sum_2[58]),
    .c(cout_3[57]),
    .cout(cout_3[58]),
    .sum(sum_3[58]));
  AL_FADD comp3_59 (
    .a(1'b0),
    .b(sum_2[59]),
    .c(cout_3[58]),
    .cout(cout_3[59]),
    .sum(sum_3[59]));
  AL_FADD comp3_6 (
    .a(i3[6]),
    .b(sum_2[6]),
    .c(cout_3[5]),
    .cout(cout_3[6]),
    .sum(sum_3[6]));
  AL_FADD comp3_60 (
    .a(1'b0),
    .b(sum_2[60]),
    .c(cout_3[59]),
    .cout(cout_3[60]),
    .sum(sum_3[60]));
  AL_FADD comp3_61 (
    .a(1'b0),
    .b(sum_2[61]),
    .c(cout_3[60]),
    .cout(cout_3[61]),
    .sum(sum_3[61]));
  AL_FADD comp3_62 (
    .a(1'b0),
    .b(sum_2[62]),
    .c(cout_3[61]),
    .cout(cout_3[62]),
    .sum(sum_3[62]));
  AL_FADD comp3_63 (
    .a(1'b0),
    .b(sum_2[63]),
    .c(cout_3[62]),
    .cout(cout_3[63]),
    .sum(sum_3[63]));
  AL_FADD comp3_7 (
    .a(i3[7]),
    .b(sum_2[7]),
    .c(cout_3[6]),
    .cout(cout_3[7]),
    .sum(sum_3[7]));
  AL_FADD comp3_8 (
    .a(i3[8]),
    .b(sum_2[8]),
    .c(cout_3[7]),
    .cout(cout_3[8]),
    .sum(sum_3[8]));
  AL_FADD comp3_9 (
    .a(i3[9]),
    .b(sum_2[9]),
    .c(cout_3[8]),
    .cout(cout_3[9]),
    .sum(sum_3[9]));
  AL_FADD comp4_0 (
    .a(i4[0]),
    .b(sum_3[0]),
    .c(1'b0),
    .cout(cout_4[0]),
    .sum(sum_4[0]));
  AL_FADD comp4_1 (
    .a(i4[1]),
    .b(sum_3[1]),
    .c(cout_4[0]),
    .cout(cout_4[1]),
    .sum(sum_4[1]));
  AL_FADD comp4_10 (
    .a(i4[10]),
    .b(sum_3[10]),
    .c(cout_4[9]),
    .cout(cout_4[10]),
    .sum(sum_4[10]));
  AL_FADD comp4_11 (
    .a(i4[11]),
    .b(sum_3[11]),
    .c(cout_4[10]),
    .cout(cout_4[11]),
    .sum(sum_4[11]));
  AL_FADD comp4_12 (
    .a(i4[12]),
    .b(sum_3[12]),
    .c(cout_4[11]),
    .cout(cout_4[12]),
    .sum(sum_4[12]));
  AL_FADD comp4_13 (
    .a(i4[13]),
    .b(sum_3[13]),
    .c(cout_4[12]),
    .cout(cout_4[13]),
    .sum(sum_4[13]));
  AL_FADD comp4_14 (
    .a(i4[14]),
    .b(sum_3[14]),
    .c(cout_4[13]),
    .cout(cout_4[14]),
    .sum(sum_4[14]));
  AL_FADD comp4_15 (
    .a(i4[15]),
    .b(sum_3[15]),
    .c(cout_4[14]),
    .cout(cout_4[15]),
    .sum(sum_4[15]));
  AL_FADD comp4_16 (
    .a(i4[16]),
    .b(sum_3[16]),
    .c(cout_4[15]),
    .cout(cout_4[16]),
    .sum(sum_4[16]));
  AL_FADD comp4_17 (
    .a(i4[17]),
    .b(sum_3[17]),
    .c(cout_4[16]),
    .cout(cout_4[17]),
    .sum(sum_4[17]));
  AL_FADD comp4_18 (
    .a(i4[18]),
    .b(sum_3[18]),
    .c(cout_4[17]),
    .cout(cout_4[18]),
    .sum(sum_4[18]));
  AL_FADD comp4_19 (
    .a(i4[19]),
    .b(sum_3[19]),
    .c(cout_4[18]),
    .cout(cout_4[19]),
    .sum(sum_4[19]));
  AL_FADD comp4_2 (
    .a(i4[2]),
    .b(sum_3[2]),
    .c(cout_4[1]),
    .cout(cout_4[2]),
    .sum(sum_4[2]));
  AL_FADD comp4_20 (
    .a(i4[20]),
    .b(sum_3[20]),
    .c(cout_4[19]),
    .cout(cout_4[20]),
    .sum(sum_4[20]));
  AL_FADD comp4_21 (
    .a(i4[21]),
    .b(sum_3[21]),
    .c(cout_4[20]),
    .cout(cout_4[21]),
    .sum(sum_4[21]));
  AL_FADD comp4_22 (
    .a(i4[22]),
    .b(sum_3[22]),
    .c(cout_4[21]),
    .cout(cout_4[22]),
    .sum(sum_4[22]));
  AL_FADD comp4_23 (
    .a(i4[23]),
    .b(sum_3[23]),
    .c(cout_4[22]),
    .cout(cout_4[23]),
    .sum(sum_4[23]));
  AL_FADD comp4_24 (
    .a(i4[24]),
    .b(sum_3[24]),
    .c(cout_4[23]),
    .cout(cout_4[24]),
    .sum(sum_4[24]));
  AL_FADD comp4_25 (
    .a(i4[25]),
    .b(sum_3[25]),
    .c(cout_4[24]),
    .cout(cout_4[25]),
    .sum(sum_4[25]));
  AL_FADD comp4_26 (
    .a(i4[26]),
    .b(sum_3[26]),
    .c(cout_4[25]),
    .cout(cout_4[26]),
    .sum(sum_4[26]));
  AL_FADD comp4_27 (
    .a(i4[27]),
    .b(sum_3[27]),
    .c(cout_4[26]),
    .cout(cout_4[27]),
    .sum(sum_4[27]));
  AL_FADD comp4_28 (
    .a(i4[28]),
    .b(sum_3[28]),
    .c(cout_4[27]),
    .cout(cout_4[28]),
    .sum(sum_4[28]));
  AL_FADD comp4_29 (
    .a(i4[29]),
    .b(sum_3[29]),
    .c(cout_4[28]),
    .cout(cout_4[29]),
    .sum(sum_4[29]));
  AL_FADD comp4_3 (
    .a(i4[3]),
    .b(sum_3[3]),
    .c(cout_4[2]),
    .cout(cout_4[3]),
    .sum(sum_4[3]));
  AL_FADD comp4_30 (
    .a(i4[30]),
    .b(sum_3[30]),
    .c(cout_4[29]),
    .cout(cout_4[30]),
    .sum(sum_4[30]));
  AL_FADD comp4_31 (
    .a(i4[31]),
    .b(sum_3[31]),
    .c(cout_4[30]),
    .cout(cout_4[31]),
    .sum(sum_4[31]));
  AL_FADD comp4_32 (
    .a(i4[32]),
    .b(sum_3[32]),
    .c(cout_4[31]),
    .cout(cout_4[32]),
    .sum(sum_4[32]));
  AL_FADD comp4_33 (
    .a(i4[33]),
    .b(sum_3[33]),
    .c(cout_4[32]),
    .cout(cout_4[33]),
    .sum(sum_4[33]));
  AL_FADD comp4_34 (
    .a(i4[34]),
    .b(sum_3[34]),
    .c(cout_4[33]),
    .cout(cout_4[34]),
    .sum(sum_4[34]));
  AL_FADD comp4_35 (
    .a(i4[35]),
    .b(sum_3[35]),
    .c(cout_4[34]),
    .cout(cout_4[35]),
    .sum(sum_4[35]));
  AL_FADD comp4_36 (
    .a(i4[36]),
    .b(sum_3[36]),
    .c(cout_4[35]),
    .cout(cout_4[36]),
    .sum(sum_4[36]));
  AL_FADD comp4_37 (
    .a(i4[37]),
    .b(sum_3[37]),
    .c(cout_4[36]),
    .cout(cout_4[37]),
    .sum(sum_4[37]));
  AL_FADD comp4_38 (
    .a(i4[38]),
    .b(sum_3[38]),
    .c(cout_4[37]),
    .cout(cout_4[38]),
    .sum(sum_4[38]));
  AL_FADD comp4_39 (
    .a(i4[39]),
    .b(sum_3[39]),
    .c(cout_4[38]),
    .cout(cout_4[39]),
    .sum(sum_4[39]));
  AL_FADD comp4_4 (
    .a(i4[4]),
    .b(sum_3[4]),
    .c(cout_4[3]),
    .cout(cout_4[4]),
    .sum(sum_4[4]));
  AL_FADD comp4_40 (
    .a(i4[40]),
    .b(sum_3[40]),
    .c(cout_4[39]),
    .cout(cout_4[40]),
    .sum(sum_4[40]));
  AL_FADD comp4_41 (
    .a(i4[41]),
    .b(sum_3[41]),
    .c(cout_4[40]),
    .cout(cout_4[41]),
    .sum(sum_4[41]));
  AL_FADD comp4_42 (
    .a(i4[42]),
    .b(sum_3[42]),
    .c(cout_4[41]),
    .cout(cout_4[42]),
    .sum(sum_4[42]));
  AL_FADD comp4_43 (
    .a(i4[43]),
    .b(sum_3[43]),
    .c(cout_4[42]),
    .cout(cout_4[43]),
    .sum(sum_4[43]));
  AL_FADD comp4_44 (
    .a(i4[44]),
    .b(sum_3[44]),
    .c(cout_4[43]),
    .cout(cout_4[44]),
    .sum(sum_4[44]));
  AL_FADD comp4_45 (
    .a(i4[45]),
    .b(sum_3[45]),
    .c(cout_4[44]),
    .cout(cout_4[45]),
    .sum(sum_4[45]));
  AL_FADD comp4_46 (
    .a(i4[46]),
    .b(sum_3[46]),
    .c(cout_4[45]),
    .cout(cout_4[46]),
    .sum(sum_4[46]));
  AL_FADD comp4_47 (
    .a(i4[47]),
    .b(sum_3[47]),
    .c(cout_4[46]),
    .cout(cout_4[47]),
    .sum(sum_4[47]));
  AL_FADD comp4_48 (
    .a(i4[48]),
    .b(sum_3[48]),
    .c(cout_4[47]),
    .cout(cout_4[48]),
    .sum(sum_4[48]));
  AL_FADD comp4_49 (
    .a(i4[49]),
    .b(sum_3[49]),
    .c(cout_4[48]),
    .cout(cout_4[49]),
    .sum(sum_4[49]));
  AL_FADD comp4_5 (
    .a(i4[5]),
    .b(sum_3[5]),
    .c(cout_4[4]),
    .cout(cout_4[5]),
    .sum(sum_4[5]));
  AL_FADD comp4_50 (
    .a(i4[50]),
    .b(sum_3[50]),
    .c(cout_4[49]),
    .cout(cout_4[50]),
    .sum(sum_4[50]));
  AL_FADD comp4_51 (
    .a(i4[51]),
    .b(sum_3[51]),
    .c(cout_4[50]),
    .cout(cout_4[51]),
    .sum(sum_4[51]));
  AL_FADD comp4_52 (
    .a(i4[52]),
    .b(sum_3[52]),
    .c(cout_4[51]),
    .cout(cout_4[52]),
    .sum(sum_4[52]));
  AL_FADD comp4_53 (
    .a(i4[53]),
    .b(sum_3[53]),
    .c(cout_4[52]),
    .cout(cout_4[53]),
    .sum(sum_4[53]));
  AL_FADD comp4_54 (
    .a(i4[54]),
    .b(sum_3[54]),
    .c(cout_4[53]),
    .cout(cout_4[54]),
    .sum(sum_4[54]));
  AL_FADD comp4_55 (
    .a(i4[55]),
    .b(sum_3[55]),
    .c(cout_4[54]),
    .cout(cout_4[55]),
    .sum(sum_4[55]));
  AL_FADD comp4_56 (
    .a(i4[56]),
    .b(sum_3[56]),
    .c(cout_4[55]),
    .cout(cout_4[56]),
    .sum(sum_4[56]));
  AL_FADD comp4_57 (
    .a(i4[57]),
    .b(sum_3[57]),
    .c(cout_4[56]),
    .cout(cout_4[57]),
    .sum(sum_4[57]));
  AL_FADD comp4_58 (
    .a(1'b0),
    .b(sum_3[58]),
    .c(cout_4[57]),
    .cout(cout_4[58]),
    .sum(sum_4[58]));
  AL_FADD comp4_59 (
    .a(1'b0),
    .b(sum_3[59]),
    .c(cout_4[58]),
    .cout(cout_4[59]),
    .sum(sum_4[59]));
  AL_FADD comp4_6 (
    .a(i4[6]),
    .b(sum_3[6]),
    .c(cout_4[5]),
    .cout(cout_4[6]),
    .sum(sum_4[6]));
  AL_FADD comp4_60 (
    .a(1'b0),
    .b(sum_3[60]),
    .c(cout_4[59]),
    .cout(cout_4[60]),
    .sum(sum_4[60]));
  AL_FADD comp4_61 (
    .a(1'b0),
    .b(sum_3[61]),
    .c(cout_4[60]),
    .cout(cout_4[61]),
    .sum(sum_4[61]));
  AL_FADD comp4_62 (
    .a(1'b0),
    .b(sum_3[62]),
    .c(cout_4[61]),
    .cout(cout_4[62]),
    .sum(sum_4[62]));
  AL_FADD comp4_63 (
    .a(1'b0),
    .b(sum_3[63]),
    .c(cout_4[62]),
    .cout(cout_4[63]),
    .sum(sum_4[63]));
  AL_FADD comp4_7 (
    .a(i4[7]),
    .b(sum_3[7]),
    .c(cout_4[6]),
    .cout(cout_4[7]),
    .sum(sum_4[7]));
  AL_FADD comp4_8 (
    .a(i4[8]),
    .b(sum_3[8]),
    .c(cout_4[7]),
    .cout(cout_4[8]),
    .sum(sum_4[8]));
  AL_FADD comp4_9 (
    .a(i4[9]),
    .b(sum_3[9]),
    .c(cout_4[8]),
    .cout(cout_4[9]),
    .sum(sum_4[9]));
  AL_FADD comp5_0 (
    .a(i5[0]),
    .b(sum_4[0]),
    .c(1'b0),
    .cout(cout_5[0]),
    .sum(sum_5[0]));
  AL_FADD comp5_1 (
    .a(i5[1]),
    .b(sum_4[1]),
    .c(cout_5[0]),
    .cout(cout_5[1]),
    .sum(sum_5[1]));
  AL_FADD comp5_10 (
    .a(i5[10]),
    .b(sum_4[10]),
    .c(cout_5[9]),
    .cout(cout_5[10]),
    .sum(sum_5[10]));
  AL_FADD comp5_11 (
    .a(i5[11]),
    .b(sum_4[11]),
    .c(cout_5[10]),
    .cout(cout_5[11]),
    .sum(sum_5[11]));
  AL_FADD comp5_12 (
    .a(i5[12]),
    .b(sum_4[12]),
    .c(cout_5[11]),
    .cout(cout_5[12]),
    .sum(sum_5[12]));
  AL_FADD comp5_13 (
    .a(i5[13]),
    .b(sum_4[13]),
    .c(cout_5[12]),
    .cout(cout_5[13]),
    .sum(sum_5[13]));
  AL_FADD comp5_14 (
    .a(i5[14]),
    .b(sum_4[14]),
    .c(cout_5[13]),
    .cout(cout_5[14]),
    .sum(sum_5[14]));
  AL_FADD comp5_15 (
    .a(i5[15]),
    .b(sum_4[15]),
    .c(cout_5[14]),
    .cout(cout_5[15]),
    .sum(sum_5[15]));
  AL_FADD comp5_16 (
    .a(i5[16]),
    .b(sum_4[16]),
    .c(cout_5[15]),
    .cout(cout_5[16]),
    .sum(sum_5[16]));
  AL_FADD comp5_17 (
    .a(i5[17]),
    .b(sum_4[17]),
    .c(cout_5[16]),
    .cout(cout_5[17]),
    .sum(sum_5[17]));
  AL_FADD comp5_18 (
    .a(i5[18]),
    .b(sum_4[18]),
    .c(cout_5[17]),
    .cout(cout_5[18]),
    .sum(sum_5[18]));
  AL_FADD comp5_19 (
    .a(i5[19]),
    .b(sum_4[19]),
    .c(cout_5[18]),
    .cout(cout_5[19]),
    .sum(sum_5[19]));
  AL_FADD comp5_2 (
    .a(i5[2]),
    .b(sum_4[2]),
    .c(cout_5[1]),
    .cout(cout_5[2]),
    .sum(sum_5[2]));
  AL_FADD comp5_20 (
    .a(i5[20]),
    .b(sum_4[20]),
    .c(cout_5[19]),
    .cout(cout_5[20]),
    .sum(sum_5[20]));
  AL_FADD comp5_21 (
    .a(i5[21]),
    .b(sum_4[21]),
    .c(cout_5[20]),
    .cout(cout_5[21]),
    .sum(sum_5[21]));
  AL_FADD comp5_22 (
    .a(i5[22]),
    .b(sum_4[22]),
    .c(cout_5[21]),
    .cout(cout_5[22]),
    .sum(sum_5[22]));
  AL_FADD comp5_23 (
    .a(i5[23]),
    .b(sum_4[23]),
    .c(cout_5[22]),
    .cout(cout_5[23]),
    .sum(sum_5[23]));
  AL_FADD comp5_24 (
    .a(i5[24]),
    .b(sum_4[24]),
    .c(cout_5[23]),
    .cout(cout_5[24]),
    .sum(sum_5[24]));
  AL_FADD comp5_25 (
    .a(i5[25]),
    .b(sum_4[25]),
    .c(cout_5[24]),
    .cout(cout_5[25]),
    .sum(sum_5[25]));
  AL_FADD comp5_26 (
    .a(i5[26]),
    .b(sum_4[26]),
    .c(cout_5[25]),
    .cout(cout_5[26]),
    .sum(sum_5[26]));
  AL_FADD comp5_27 (
    .a(i5[27]),
    .b(sum_4[27]),
    .c(cout_5[26]),
    .cout(cout_5[27]),
    .sum(sum_5[27]));
  AL_FADD comp5_28 (
    .a(i5[28]),
    .b(sum_4[28]),
    .c(cout_5[27]),
    .cout(cout_5[28]),
    .sum(sum_5[28]));
  AL_FADD comp5_29 (
    .a(i5[29]),
    .b(sum_4[29]),
    .c(cout_5[28]),
    .cout(cout_5[29]),
    .sum(sum_5[29]));
  AL_FADD comp5_3 (
    .a(i5[3]),
    .b(sum_4[3]),
    .c(cout_5[2]),
    .cout(cout_5[3]),
    .sum(sum_5[3]));
  AL_FADD comp5_30 (
    .a(i5[30]),
    .b(sum_4[30]),
    .c(cout_5[29]),
    .cout(cout_5[30]),
    .sum(sum_5[30]));
  AL_FADD comp5_31 (
    .a(i5[31]),
    .b(sum_4[31]),
    .c(cout_5[30]),
    .cout(cout_5[31]),
    .sum(sum_5[31]));
  AL_FADD comp5_32 (
    .a(i5[32]),
    .b(sum_4[32]),
    .c(cout_5[31]),
    .cout(cout_5[32]),
    .sum(sum_5[32]));
  AL_FADD comp5_33 (
    .a(i5[33]),
    .b(sum_4[33]),
    .c(cout_5[32]),
    .cout(cout_5[33]),
    .sum(sum_5[33]));
  AL_FADD comp5_34 (
    .a(i5[34]),
    .b(sum_4[34]),
    .c(cout_5[33]),
    .cout(cout_5[34]),
    .sum(sum_5[34]));
  AL_FADD comp5_35 (
    .a(i5[35]),
    .b(sum_4[35]),
    .c(cout_5[34]),
    .cout(cout_5[35]),
    .sum(sum_5[35]));
  AL_FADD comp5_36 (
    .a(i5[36]),
    .b(sum_4[36]),
    .c(cout_5[35]),
    .cout(cout_5[36]),
    .sum(sum_5[36]));
  AL_FADD comp5_37 (
    .a(i5[37]),
    .b(sum_4[37]),
    .c(cout_5[36]),
    .cout(cout_5[37]),
    .sum(sum_5[37]));
  AL_FADD comp5_38 (
    .a(i5[38]),
    .b(sum_4[38]),
    .c(cout_5[37]),
    .cout(cout_5[38]),
    .sum(sum_5[38]));
  AL_FADD comp5_39 (
    .a(i5[39]),
    .b(sum_4[39]),
    .c(cout_5[38]),
    .cout(cout_5[39]),
    .sum(sum_5[39]));
  AL_FADD comp5_4 (
    .a(i5[4]),
    .b(sum_4[4]),
    .c(cout_5[3]),
    .cout(cout_5[4]),
    .sum(sum_5[4]));
  AL_FADD comp5_40 (
    .a(i5[40]),
    .b(sum_4[40]),
    .c(cout_5[39]),
    .cout(cout_5[40]),
    .sum(sum_5[40]));
  AL_FADD comp5_41 (
    .a(i5[41]),
    .b(sum_4[41]),
    .c(cout_5[40]),
    .cout(cout_5[41]),
    .sum(sum_5[41]));
  AL_FADD comp5_42 (
    .a(i5[42]),
    .b(sum_4[42]),
    .c(cout_5[41]),
    .cout(cout_5[42]),
    .sum(sum_5[42]));
  AL_FADD comp5_43 (
    .a(i5[43]),
    .b(sum_4[43]),
    .c(cout_5[42]),
    .cout(cout_5[43]),
    .sum(sum_5[43]));
  AL_FADD comp5_44 (
    .a(i5[44]),
    .b(sum_4[44]),
    .c(cout_5[43]),
    .cout(cout_5[44]),
    .sum(sum_5[44]));
  AL_FADD comp5_45 (
    .a(i5[45]),
    .b(sum_4[45]),
    .c(cout_5[44]),
    .cout(cout_5[45]),
    .sum(sum_5[45]));
  AL_FADD comp5_46 (
    .a(i5[46]),
    .b(sum_4[46]),
    .c(cout_5[45]),
    .cout(cout_5[46]),
    .sum(sum_5[46]));
  AL_FADD comp5_47 (
    .a(i5[47]),
    .b(sum_4[47]),
    .c(cout_5[46]),
    .cout(cout_5[47]),
    .sum(sum_5[47]));
  AL_FADD comp5_48 (
    .a(i5[48]),
    .b(sum_4[48]),
    .c(cout_5[47]),
    .cout(cout_5[48]),
    .sum(sum_5[48]));
  AL_FADD comp5_49 (
    .a(i5[49]),
    .b(sum_4[49]),
    .c(cout_5[48]),
    .cout(cout_5[49]),
    .sum(sum_5[49]));
  AL_FADD comp5_5 (
    .a(i5[5]),
    .b(sum_4[5]),
    .c(cout_5[4]),
    .cout(cout_5[5]),
    .sum(sum_5[5]));
  AL_FADD comp5_50 (
    .a(i5[50]),
    .b(sum_4[50]),
    .c(cout_5[49]),
    .cout(cout_5[50]),
    .sum(sum_5[50]));
  AL_FADD comp5_51 (
    .a(i5[51]),
    .b(sum_4[51]),
    .c(cout_5[50]),
    .cout(cout_5[51]),
    .sum(sum_5[51]));
  AL_FADD comp5_52 (
    .a(i5[52]),
    .b(sum_4[52]),
    .c(cout_5[51]),
    .cout(cout_5[52]),
    .sum(sum_5[52]));
  AL_FADD comp5_53 (
    .a(i5[53]),
    .b(sum_4[53]),
    .c(cout_5[52]),
    .cout(cout_5[53]),
    .sum(sum_5[53]));
  AL_FADD comp5_54 (
    .a(i5[54]),
    .b(sum_4[54]),
    .c(cout_5[53]),
    .cout(cout_5[54]),
    .sum(sum_5[54]));
  AL_FADD comp5_55 (
    .a(i5[55]),
    .b(sum_4[55]),
    .c(cout_5[54]),
    .cout(cout_5[55]),
    .sum(sum_5[55]));
  AL_FADD comp5_56 (
    .a(i5[56]),
    .b(sum_4[56]),
    .c(cout_5[55]),
    .cout(cout_5[56]),
    .sum(sum_5[56]));
  AL_FADD comp5_57 (
    .a(1'b0),
    .b(sum_4[57]),
    .c(cout_5[56]),
    .cout(cout_5[57]),
    .sum(sum_5[57]));
  AL_FADD comp5_58 (
    .a(1'b0),
    .b(sum_4[58]),
    .c(cout_5[57]),
    .cout(cout_5[58]),
    .sum(sum_5[58]));
  AL_FADD comp5_59 (
    .a(1'b0),
    .b(sum_4[59]),
    .c(cout_5[58]),
    .cout(cout_5[59]),
    .sum(sum_5[59]));
  AL_FADD comp5_6 (
    .a(i5[6]),
    .b(sum_4[6]),
    .c(cout_5[5]),
    .cout(cout_5[6]),
    .sum(sum_5[6]));
  AL_FADD comp5_60 (
    .a(1'b0),
    .b(sum_4[60]),
    .c(cout_5[59]),
    .cout(cout_5[60]),
    .sum(sum_5[60]));
  AL_FADD comp5_61 (
    .a(1'b0),
    .b(sum_4[61]),
    .c(cout_5[60]),
    .cout(cout_5[61]),
    .sum(sum_5[61]));
  AL_FADD comp5_62 (
    .a(1'b0),
    .b(sum_4[62]),
    .c(cout_5[61]),
    .cout(cout_5[62]),
    .sum(sum_5[62]));
  AL_FADD comp5_63 (
    .a(1'b0),
    .b(sum_4[63]),
    .c(cout_5[62]),
    .cout(cout_5[63]),
    .sum(sum_5[63]));
  AL_FADD comp5_7 (
    .a(i5[7]),
    .b(sum_4[7]),
    .c(cout_5[6]),
    .cout(cout_5[7]),
    .sum(sum_5[7]));
  AL_FADD comp5_8 (
    .a(i5[8]),
    .b(sum_4[8]),
    .c(cout_5[7]),
    .cout(cout_5[8]),
    .sum(sum_5[8]));
  AL_FADD comp5_9 (
    .a(i5[9]),
    .b(sum_4[9]),
    .c(cout_5[8]),
    .cout(cout_5[9]),
    .sum(sum_5[9]));
  AL_FADD comp6_0 (
    .a(i6[0]),
    .b(sum_5[0]),
    .c(1'b0),
    .cout(cout_6[0]),
    .sum(sum_6[0]));
  AL_FADD comp6_1 (
    .a(i6[1]),
    .b(sum_5[1]),
    .c(cout_6[0]),
    .cout(cout_6[1]),
    .sum(sum_6[1]));
  AL_FADD comp6_10 (
    .a(i6[10]),
    .b(sum_5[10]),
    .c(cout_6[9]),
    .cout(cout_6[10]),
    .sum(sum_6[10]));
  AL_FADD comp6_11 (
    .a(i6[11]),
    .b(sum_5[11]),
    .c(cout_6[10]),
    .cout(cout_6[11]),
    .sum(sum_6[11]));
  AL_FADD comp6_12 (
    .a(i6[12]),
    .b(sum_5[12]),
    .c(cout_6[11]),
    .cout(cout_6[12]),
    .sum(sum_6[12]));
  AL_FADD comp6_13 (
    .a(i6[13]),
    .b(sum_5[13]),
    .c(cout_6[12]),
    .cout(cout_6[13]),
    .sum(sum_6[13]));
  AL_FADD comp6_14 (
    .a(i6[14]),
    .b(sum_5[14]),
    .c(cout_6[13]),
    .cout(cout_6[14]),
    .sum(sum_6[14]));
  AL_FADD comp6_15 (
    .a(i6[15]),
    .b(sum_5[15]),
    .c(cout_6[14]),
    .cout(cout_6[15]),
    .sum(sum_6[15]));
  AL_FADD comp6_16 (
    .a(i6[16]),
    .b(sum_5[16]),
    .c(cout_6[15]),
    .cout(cout_6[16]),
    .sum(sum_6[16]));
  AL_FADD comp6_17 (
    .a(i6[17]),
    .b(sum_5[17]),
    .c(cout_6[16]),
    .cout(cout_6[17]),
    .sum(sum_6[17]));
  AL_FADD comp6_18 (
    .a(i6[18]),
    .b(sum_5[18]),
    .c(cout_6[17]),
    .cout(cout_6[18]),
    .sum(sum_6[18]));
  AL_FADD comp6_19 (
    .a(i6[19]),
    .b(sum_5[19]),
    .c(cout_6[18]),
    .cout(cout_6[19]),
    .sum(sum_6[19]));
  AL_FADD comp6_2 (
    .a(i6[2]),
    .b(sum_5[2]),
    .c(cout_6[1]),
    .cout(cout_6[2]),
    .sum(sum_6[2]));
  AL_FADD comp6_20 (
    .a(i6[20]),
    .b(sum_5[20]),
    .c(cout_6[19]),
    .cout(cout_6[20]),
    .sum(sum_6[20]));
  AL_FADD comp6_21 (
    .a(i6[21]),
    .b(sum_5[21]),
    .c(cout_6[20]),
    .cout(cout_6[21]),
    .sum(sum_6[21]));
  AL_FADD comp6_22 (
    .a(i6[22]),
    .b(sum_5[22]),
    .c(cout_6[21]),
    .cout(cout_6[22]),
    .sum(sum_6[22]));
  AL_FADD comp6_23 (
    .a(i6[23]),
    .b(sum_5[23]),
    .c(cout_6[22]),
    .cout(cout_6[23]),
    .sum(sum_6[23]));
  AL_FADD comp6_24 (
    .a(i6[24]),
    .b(sum_5[24]),
    .c(cout_6[23]),
    .cout(cout_6[24]),
    .sum(sum_6[24]));
  AL_FADD comp6_25 (
    .a(i6[25]),
    .b(sum_5[25]),
    .c(cout_6[24]),
    .cout(cout_6[25]),
    .sum(sum_6[25]));
  AL_FADD comp6_26 (
    .a(i6[26]),
    .b(sum_5[26]),
    .c(cout_6[25]),
    .cout(cout_6[26]),
    .sum(sum_6[26]));
  AL_FADD comp6_27 (
    .a(i6[27]),
    .b(sum_5[27]),
    .c(cout_6[26]),
    .cout(cout_6[27]),
    .sum(sum_6[27]));
  AL_FADD comp6_28 (
    .a(i6[28]),
    .b(sum_5[28]),
    .c(cout_6[27]),
    .cout(cout_6[28]),
    .sum(sum_6[28]));
  AL_FADD comp6_29 (
    .a(i6[29]),
    .b(sum_5[29]),
    .c(cout_6[28]),
    .cout(cout_6[29]),
    .sum(sum_6[29]));
  AL_FADD comp6_3 (
    .a(i6[3]),
    .b(sum_5[3]),
    .c(cout_6[2]),
    .cout(cout_6[3]),
    .sum(sum_6[3]));
  AL_FADD comp6_30 (
    .a(i6[30]),
    .b(sum_5[30]),
    .c(cout_6[29]),
    .cout(cout_6[30]),
    .sum(sum_6[30]));
  AL_FADD comp6_31 (
    .a(i6[31]),
    .b(sum_5[31]),
    .c(cout_6[30]),
    .cout(cout_6[31]),
    .sum(sum_6[31]));
  AL_FADD comp6_32 (
    .a(i6[32]),
    .b(sum_5[32]),
    .c(cout_6[31]),
    .cout(cout_6[32]),
    .sum(sum_6[32]));
  AL_FADD comp6_33 (
    .a(i6[33]),
    .b(sum_5[33]),
    .c(cout_6[32]),
    .cout(cout_6[33]),
    .sum(sum_6[33]));
  AL_FADD comp6_34 (
    .a(i6[34]),
    .b(sum_5[34]),
    .c(cout_6[33]),
    .cout(cout_6[34]),
    .sum(sum_6[34]));
  AL_FADD comp6_35 (
    .a(i6[35]),
    .b(sum_5[35]),
    .c(cout_6[34]),
    .cout(cout_6[35]),
    .sum(sum_6[35]));
  AL_FADD comp6_36 (
    .a(i6[36]),
    .b(sum_5[36]),
    .c(cout_6[35]),
    .cout(cout_6[36]),
    .sum(sum_6[36]));
  AL_FADD comp6_37 (
    .a(i6[37]),
    .b(sum_5[37]),
    .c(cout_6[36]),
    .cout(cout_6[37]),
    .sum(sum_6[37]));
  AL_FADD comp6_38 (
    .a(i6[38]),
    .b(sum_5[38]),
    .c(cout_6[37]),
    .cout(cout_6[38]),
    .sum(sum_6[38]));
  AL_FADD comp6_39 (
    .a(i6[39]),
    .b(sum_5[39]),
    .c(cout_6[38]),
    .cout(cout_6[39]),
    .sum(sum_6[39]));
  AL_FADD comp6_4 (
    .a(i6[4]),
    .b(sum_5[4]),
    .c(cout_6[3]),
    .cout(cout_6[4]),
    .sum(sum_6[4]));
  AL_FADD comp6_40 (
    .a(i6[40]),
    .b(sum_5[40]),
    .c(cout_6[39]),
    .cout(cout_6[40]),
    .sum(sum_6[40]));
  AL_FADD comp6_41 (
    .a(i6[41]),
    .b(sum_5[41]),
    .c(cout_6[40]),
    .cout(cout_6[41]),
    .sum(sum_6[41]));
  AL_FADD comp6_42 (
    .a(i6[42]),
    .b(sum_5[42]),
    .c(cout_6[41]),
    .cout(cout_6[42]),
    .sum(sum_6[42]));
  AL_FADD comp6_43 (
    .a(i6[43]),
    .b(sum_5[43]),
    .c(cout_6[42]),
    .cout(cout_6[43]),
    .sum(sum_6[43]));
  AL_FADD comp6_44 (
    .a(i6[44]),
    .b(sum_5[44]),
    .c(cout_6[43]),
    .cout(cout_6[44]),
    .sum(sum_6[44]));
  AL_FADD comp6_45 (
    .a(i6[45]),
    .b(sum_5[45]),
    .c(cout_6[44]),
    .cout(cout_6[45]),
    .sum(sum_6[45]));
  AL_FADD comp6_46 (
    .a(i6[46]),
    .b(sum_5[46]),
    .c(cout_6[45]),
    .cout(cout_6[46]),
    .sum(sum_6[46]));
  AL_FADD comp6_47 (
    .a(i6[47]),
    .b(sum_5[47]),
    .c(cout_6[46]),
    .cout(cout_6[47]),
    .sum(sum_6[47]));
  AL_FADD comp6_48 (
    .a(i6[48]),
    .b(sum_5[48]),
    .c(cout_6[47]),
    .cout(cout_6[48]),
    .sum(sum_6[48]));
  AL_FADD comp6_49 (
    .a(i6[49]),
    .b(sum_5[49]),
    .c(cout_6[48]),
    .cout(cout_6[49]),
    .sum(sum_6[49]));
  AL_FADD comp6_5 (
    .a(i6[5]),
    .b(sum_5[5]),
    .c(cout_6[4]),
    .cout(cout_6[5]),
    .sum(sum_6[5]));
  AL_FADD comp6_50 (
    .a(i6[50]),
    .b(sum_5[50]),
    .c(cout_6[49]),
    .cout(cout_6[50]),
    .sum(sum_6[50]));
  AL_FADD comp6_51 (
    .a(i6[51]),
    .b(sum_5[51]),
    .c(cout_6[50]),
    .cout(cout_6[51]),
    .sum(sum_6[51]));
  AL_FADD comp6_52 (
    .a(i6[52]),
    .b(sum_5[52]),
    .c(cout_6[51]),
    .cout(cout_6[52]),
    .sum(sum_6[52]));
  AL_FADD comp6_53 (
    .a(i6[53]),
    .b(sum_5[53]),
    .c(cout_6[52]),
    .cout(cout_6[53]),
    .sum(sum_6[53]));
  AL_FADD comp6_54 (
    .a(i6[54]),
    .b(sum_5[54]),
    .c(cout_6[53]),
    .cout(cout_6[54]),
    .sum(sum_6[54]));
  AL_FADD comp6_55 (
    .a(i6[55]),
    .b(sum_5[55]),
    .c(cout_6[54]),
    .cout(cout_6[55]),
    .sum(sum_6[55]));
  AL_FADD comp6_56 (
    .a(1'b0),
    .b(sum_5[56]),
    .c(cout_6[55]),
    .cout(cout_6[56]),
    .sum(sum_6[56]));
  AL_FADD comp6_57 (
    .a(1'b0),
    .b(sum_5[57]),
    .c(cout_6[56]),
    .cout(cout_6[57]),
    .sum(sum_6[57]));
  AL_FADD comp6_58 (
    .a(1'b0),
    .b(sum_5[58]),
    .c(cout_6[57]),
    .cout(cout_6[58]),
    .sum(sum_6[58]));
  AL_FADD comp6_59 (
    .a(1'b0),
    .b(sum_5[59]),
    .c(cout_6[58]),
    .cout(cout_6[59]),
    .sum(sum_6[59]));
  AL_FADD comp6_6 (
    .a(i6[6]),
    .b(sum_5[6]),
    .c(cout_6[5]),
    .cout(cout_6[6]),
    .sum(sum_6[6]));
  AL_FADD comp6_60 (
    .a(1'b0),
    .b(sum_5[60]),
    .c(cout_6[59]),
    .cout(cout_6[60]),
    .sum(sum_6[60]));
  AL_FADD comp6_61 (
    .a(1'b0),
    .b(sum_5[61]),
    .c(cout_6[60]),
    .cout(cout_6[61]),
    .sum(sum_6[61]));
  AL_FADD comp6_62 (
    .a(1'b0),
    .b(sum_5[62]),
    .c(cout_6[61]),
    .cout(cout_6[62]),
    .sum(sum_6[62]));
  AL_FADD comp6_63 (
    .a(1'b0),
    .b(sum_5[63]),
    .c(cout_6[62]),
    .cout(cout_6[63]),
    .sum(sum_6[63]));
  AL_FADD comp6_7 (
    .a(i6[7]),
    .b(sum_5[7]),
    .c(cout_6[6]),
    .cout(cout_6[7]),
    .sum(sum_6[7]));
  AL_FADD comp6_8 (
    .a(i6[8]),
    .b(sum_5[8]),
    .c(cout_6[7]),
    .cout(cout_6[8]),
    .sum(sum_6[8]));
  AL_FADD comp6_9 (
    .a(i6[9]),
    .b(sum_5[9]),
    .c(cout_6[8]),
    .cout(cout_6[9]),
    .sum(sum_6[9]));
  AL_FADD comp7_0 (
    .a(i7[0]),
    .b(sum_6[0]),
    .c(1'b0),
    .cout(cout_7[0]),
    .sum(sum_7[0]));
  AL_FADD comp7_1 (
    .a(i7[1]),
    .b(sum_6[1]),
    .c(cout_7[0]),
    .cout(cout_7[1]),
    .sum(sum_7[1]));
  AL_FADD comp7_10 (
    .a(i7[10]),
    .b(sum_6[10]),
    .c(cout_7[9]),
    .cout(cout_7[10]),
    .sum(sum_7[10]));
  AL_FADD comp7_11 (
    .a(i7[11]),
    .b(sum_6[11]),
    .c(cout_7[10]),
    .cout(cout_7[11]),
    .sum(sum_7[11]));
  AL_FADD comp7_12 (
    .a(i7[12]),
    .b(sum_6[12]),
    .c(cout_7[11]),
    .cout(cout_7[12]),
    .sum(sum_7[12]));
  AL_FADD comp7_13 (
    .a(i7[13]),
    .b(sum_6[13]),
    .c(cout_7[12]),
    .cout(cout_7[13]),
    .sum(sum_7[13]));
  AL_FADD comp7_14 (
    .a(i7[14]),
    .b(sum_6[14]),
    .c(cout_7[13]),
    .cout(cout_7[14]),
    .sum(sum_7[14]));
  AL_FADD comp7_15 (
    .a(i7[15]),
    .b(sum_6[15]),
    .c(cout_7[14]),
    .cout(cout_7[15]),
    .sum(sum_7[15]));
  AL_FADD comp7_16 (
    .a(i7[16]),
    .b(sum_6[16]),
    .c(cout_7[15]),
    .cout(cout_7[16]),
    .sum(sum_7[16]));
  AL_FADD comp7_17 (
    .a(i7[17]),
    .b(sum_6[17]),
    .c(cout_7[16]),
    .cout(cout_7[17]),
    .sum(sum_7[17]));
  AL_FADD comp7_18 (
    .a(i7[18]),
    .b(sum_6[18]),
    .c(cout_7[17]),
    .cout(cout_7[18]),
    .sum(sum_7[18]));
  AL_FADD comp7_19 (
    .a(i7[19]),
    .b(sum_6[19]),
    .c(cout_7[18]),
    .cout(cout_7[19]),
    .sum(sum_7[19]));
  AL_FADD comp7_2 (
    .a(i7[2]),
    .b(sum_6[2]),
    .c(cout_7[1]),
    .cout(cout_7[2]),
    .sum(sum_7[2]));
  AL_FADD comp7_20 (
    .a(i7[20]),
    .b(sum_6[20]),
    .c(cout_7[19]),
    .cout(cout_7[20]),
    .sum(sum_7[20]));
  AL_FADD comp7_21 (
    .a(i7[21]),
    .b(sum_6[21]),
    .c(cout_7[20]),
    .cout(cout_7[21]),
    .sum(sum_7[21]));
  AL_FADD comp7_22 (
    .a(i7[22]),
    .b(sum_6[22]),
    .c(cout_7[21]),
    .cout(cout_7[22]),
    .sum(sum_7[22]));
  AL_FADD comp7_23 (
    .a(i7[23]),
    .b(sum_6[23]),
    .c(cout_7[22]),
    .cout(cout_7[23]),
    .sum(sum_7[23]));
  AL_FADD comp7_24 (
    .a(i7[24]),
    .b(sum_6[24]),
    .c(cout_7[23]),
    .cout(cout_7[24]),
    .sum(sum_7[24]));
  AL_FADD comp7_25 (
    .a(i7[25]),
    .b(sum_6[25]),
    .c(cout_7[24]),
    .cout(cout_7[25]),
    .sum(sum_7[25]));
  AL_FADD comp7_26 (
    .a(i7[26]),
    .b(sum_6[26]),
    .c(cout_7[25]),
    .cout(cout_7[26]),
    .sum(sum_7[26]));
  AL_FADD comp7_27 (
    .a(i7[27]),
    .b(sum_6[27]),
    .c(cout_7[26]),
    .cout(cout_7[27]),
    .sum(sum_7[27]));
  AL_FADD comp7_28 (
    .a(i7[28]),
    .b(sum_6[28]),
    .c(cout_7[27]),
    .cout(cout_7[28]),
    .sum(sum_7[28]));
  AL_FADD comp7_29 (
    .a(i7[29]),
    .b(sum_6[29]),
    .c(cout_7[28]),
    .cout(cout_7[29]),
    .sum(sum_7[29]));
  AL_FADD comp7_3 (
    .a(i7[3]),
    .b(sum_6[3]),
    .c(cout_7[2]),
    .cout(cout_7[3]),
    .sum(sum_7[3]));
  AL_FADD comp7_30 (
    .a(i7[30]),
    .b(sum_6[30]),
    .c(cout_7[29]),
    .cout(cout_7[30]),
    .sum(sum_7[30]));
  AL_FADD comp7_31 (
    .a(i7[31]),
    .b(sum_6[31]),
    .c(cout_7[30]),
    .cout(cout_7[31]),
    .sum(sum_7[31]));
  AL_FADD comp7_32 (
    .a(i7[32]),
    .b(sum_6[32]),
    .c(cout_7[31]),
    .cout(cout_7[32]),
    .sum(sum_7[32]));
  AL_FADD comp7_33 (
    .a(i7[33]),
    .b(sum_6[33]),
    .c(cout_7[32]),
    .cout(cout_7[33]),
    .sum(sum_7[33]));
  AL_FADD comp7_34 (
    .a(i7[34]),
    .b(sum_6[34]),
    .c(cout_7[33]),
    .cout(cout_7[34]),
    .sum(sum_7[34]));
  AL_FADD comp7_35 (
    .a(i7[35]),
    .b(sum_6[35]),
    .c(cout_7[34]),
    .cout(cout_7[35]),
    .sum(sum_7[35]));
  AL_FADD comp7_36 (
    .a(i7[36]),
    .b(sum_6[36]),
    .c(cout_7[35]),
    .cout(cout_7[36]),
    .sum(sum_7[36]));
  AL_FADD comp7_37 (
    .a(i7[37]),
    .b(sum_6[37]),
    .c(cout_7[36]),
    .cout(cout_7[37]),
    .sum(sum_7[37]));
  AL_FADD comp7_38 (
    .a(i7[38]),
    .b(sum_6[38]),
    .c(cout_7[37]),
    .cout(cout_7[38]),
    .sum(sum_7[38]));
  AL_FADD comp7_39 (
    .a(i7[39]),
    .b(sum_6[39]),
    .c(cout_7[38]),
    .cout(cout_7[39]),
    .sum(sum_7[39]));
  AL_FADD comp7_4 (
    .a(i7[4]),
    .b(sum_6[4]),
    .c(cout_7[3]),
    .cout(cout_7[4]),
    .sum(sum_7[4]));
  AL_FADD comp7_40 (
    .a(i7[40]),
    .b(sum_6[40]),
    .c(cout_7[39]),
    .cout(cout_7[40]),
    .sum(sum_7[40]));
  AL_FADD comp7_41 (
    .a(i7[41]),
    .b(sum_6[41]),
    .c(cout_7[40]),
    .cout(cout_7[41]),
    .sum(sum_7[41]));
  AL_FADD comp7_42 (
    .a(i7[42]),
    .b(sum_6[42]),
    .c(cout_7[41]),
    .cout(cout_7[42]),
    .sum(sum_7[42]));
  AL_FADD comp7_43 (
    .a(i7[43]),
    .b(sum_6[43]),
    .c(cout_7[42]),
    .cout(cout_7[43]),
    .sum(sum_7[43]));
  AL_FADD comp7_44 (
    .a(i7[44]),
    .b(sum_6[44]),
    .c(cout_7[43]),
    .cout(cout_7[44]),
    .sum(sum_7[44]));
  AL_FADD comp7_45 (
    .a(i7[45]),
    .b(sum_6[45]),
    .c(cout_7[44]),
    .cout(cout_7[45]),
    .sum(sum_7[45]));
  AL_FADD comp7_46 (
    .a(i7[46]),
    .b(sum_6[46]),
    .c(cout_7[45]),
    .cout(cout_7[46]),
    .sum(sum_7[46]));
  AL_FADD comp7_47 (
    .a(i7[47]),
    .b(sum_6[47]),
    .c(cout_7[46]),
    .cout(cout_7[47]),
    .sum(sum_7[47]));
  AL_FADD comp7_48 (
    .a(i7[48]),
    .b(sum_6[48]),
    .c(cout_7[47]),
    .cout(cout_7[48]),
    .sum(sum_7[48]));
  AL_FADD comp7_49 (
    .a(i7[49]),
    .b(sum_6[49]),
    .c(cout_7[48]),
    .cout(cout_7[49]),
    .sum(sum_7[49]));
  AL_FADD comp7_5 (
    .a(i7[5]),
    .b(sum_6[5]),
    .c(cout_7[4]),
    .cout(cout_7[5]),
    .sum(sum_7[5]));
  AL_FADD comp7_50 (
    .a(i7[50]),
    .b(sum_6[50]),
    .c(cout_7[49]),
    .cout(cout_7[50]),
    .sum(sum_7[50]));
  AL_FADD comp7_51 (
    .a(i7[51]),
    .b(sum_6[51]),
    .c(cout_7[50]),
    .cout(cout_7[51]),
    .sum(sum_7[51]));
  AL_FADD comp7_52 (
    .a(i7[52]),
    .b(sum_6[52]),
    .c(cout_7[51]),
    .cout(cout_7[52]),
    .sum(sum_7[52]));
  AL_FADD comp7_53 (
    .a(i7[53]),
    .b(sum_6[53]),
    .c(cout_7[52]),
    .cout(cout_7[53]),
    .sum(sum_7[53]));
  AL_FADD comp7_54 (
    .a(i7[54]),
    .b(sum_6[54]),
    .c(cout_7[53]),
    .cout(cout_7[54]),
    .sum(sum_7[54]));
  AL_FADD comp7_55 (
    .a(1'b0),
    .b(sum_6[55]),
    .c(cout_7[54]),
    .cout(cout_7[55]),
    .sum(sum_7[55]));
  AL_FADD comp7_56 (
    .a(1'b0),
    .b(sum_6[56]),
    .c(cout_7[55]),
    .cout(cout_7[56]),
    .sum(sum_7[56]));
  AL_FADD comp7_57 (
    .a(1'b0),
    .b(sum_6[57]),
    .c(cout_7[56]),
    .cout(cout_7[57]),
    .sum(sum_7[57]));
  AL_FADD comp7_58 (
    .a(1'b0),
    .b(sum_6[58]),
    .c(cout_7[57]),
    .cout(cout_7[58]),
    .sum(sum_7[58]));
  AL_FADD comp7_59 (
    .a(1'b0),
    .b(sum_6[59]),
    .c(cout_7[58]),
    .cout(cout_7[59]),
    .sum(sum_7[59]));
  AL_FADD comp7_6 (
    .a(i7[6]),
    .b(sum_6[6]),
    .c(cout_7[5]),
    .cout(cout_7[6]),
    .sum(sum_7[6]));
  AL_FADD comp7_60 (
    .a(1'b0),
    .b(sum_6[60]),
    .c(cout_7[59]),
    .cout(cout_7[60]),
    .sum(sum_7[60]));
  AL_FADD comp7_61 (
    .a(1'b0),
    .b(sum_6[61]),
    .c(cout_7[60]),
    .cout(cout_7[61]),
    .sum(sum_7[61]));
  AL_FADD comp7_62 (
    .a(1'b0),
    .b(sum_6[62]),
    .c(cout_7[61]),
    .cout(cout_7[62]),
    .sum(sum_7[62]));
  AL_FADD comp7_63 (
    .a(1'b0),
    .b(sum_6[63]),
    .c(cout_7[62]),
    .cout(cout_7[63]),
    .sum(sum_7[63]));
  AL_FADD comp7_7 (
    .a(i7[7]),
    .b(sum_6[7]),
    .c(cout_7[6]),
    .cout(cout_7[7]),
    .sum(sum_7[7]));
  AL_FADD comp7_8 (
    .a(i7[8]),
    .b(sum_6[8]),
    .c(cout_7[7]),
    .cout(cout_7[8]),
    .sum(sum_7[8]));
  AL_FADD comp7_9 (
    .a(i7[9]),
    .b(sum_6[9]),
    .c(cout_7[8]),
    .cout(cout_7[9]),
    .sum(sum_7[9]));
  AL_FADD comp8_0 (
    .a(i8[0]),
    .b(sum_7[0]),
    .c(1'b0),
    .cout(cout_8[0]),
    .sum(sum_8[0]));
  AL_FADD comp8_1 (
    .a(i8[1]),
    .b(sum_7[1]),
    .c(cout_8[0]),
    .cout(cout_8[1]),
    .sum(sum_8[1]));
  AL_FADD comp8_10 (
    .a(i8[10]),
    .b(sum_7[10]),
    .c(cout_8[9]),
    .cout(cout_8[10]),
    .sum(sum_8[10]));
  AL_FADD comp8_11 (
    .a(i8[11]),
    .b(sum_7[11]),
    .c(cout_8[10]),
    .cout(cout_8[11]),
    .sum(sum_8[11]));
  AL_FADD comp8_12 (
    .a(i8[12]),
    .b(sum_7[12]),
    .c(cout_8[11]),
    .cout(cout_8[12]),
    .sum(sum_8[12]));
  AL_FADD comp8_13 (
    .a(i8[13]),
    .b(sum_7[13]),
    .c(cout_8[12]),
    .cout(cout_8[13]),
    .sum(sum_8[13]));
  AL_FADD comp8_14 (
    .a(i8[14]),
    .b(sum_7[14]),
    .c(cout_8[13]),
    .cout(cout_8[14]),
    .sum(sum_8[14]));
  AL_FADD comp8_15 (
    .a(i8[15]),
    .b(sum_7[15]),
    .c(cout_8[14]),
    .cout(cout_8[15]),
    .sum(sum_8[15]));
  AL_FADD comp8_16 (
    .a(i8[16]),
    .b(sum_7[16]),
    .c(cout_8[15]),
    .cout(cout_8[16]),
    .sum(sum_8[16]));
  AL_FADD comp8_17 (
    .a(i8[17]),
    .b(sum_7[17]),
    .c(cout_8[16]),
    .cout(cout_8[17]),
    .sum(sum_8[17]));
  AL_FADD comp8_18 (
    .a(i8[18]),
    .b(sum_7[18]),
    .c(cout_8[17]),
    .cout(cout_8[18]),
    .sum(sum_8[18]));
  AL_FADD comp8_19 (
    .a(i8[19]),
    .b(sum_7[19]),
    .c(cout_8[18]),
    .cout(cout_8[19]),
    .sum(sum_8[19]));
  AL_FADD comp8_2 (
    .a(i8[2]),
    .b(sum_7[2]),
    .c(cout_8[1]),
    .cout(cout_8[2]),
    .sum(sum_8[2]));
  AL_FADD comp8_20 (
    .a(i8[20]),
    .b(sum_7[20]),
    .c(cout_8[19]),
    .cout(cout_8[20]),
    .sum(sum_8[20]));
  AL_FADD comp8_21 (
    .a(i8[21]),
    .b(sum_7[21]),
    .c(cout_8[20]),
    .cout(cout_8[21]),
    .sum(sum_8[21]));
  AL_FADD comp8_22 (
    .a(i8[22]),
    .b(sum_7[22]),
    .c(cout_8[21]),
    .cout(cout_8[22]),
    .sum(sum_8[22]));
  AL_FADD comp8_23 (
    .a(i8[23]),
    .b(sum_7[23]),
    .c(cout_8[22]),
    .cout(cout_8[23]),
    .sum(sum_8[23]));
  AL_FADD comp8_24 (
    .a(i8[24]),
    .b(sum_7[24]),
    .c(cout_8[23]),
    .cout(cout_8[24]),
    .sum(sum_8[24]));
  AL_FADD comp8_25 (
    .a(i8[25]),
    .b(sum_7[25]),
    .c(cout_8[24]),
    .cout(cout_8[25]),
    .sum(sum_8[25]));
  AL_FADD comp8_26 (
    .a(i8[26]),
    .b(sum_7[26]),
    .c(cout_8[25]),
    .cout(cout_8[26]),
    .sum(sum_8[26]));
  AL_FADD comp8_27 (
    .a(i8[27]),
    .b(sum_7[27]),
    .c(cout_8[26]),
    .cout(cout_8[27]),
    .sum(sum_8[27]));
  AL_FADD comp8_28 (
    .a(i8[28]),
    .b(sum_7[28]),
    .c(cout_8[27]),
    .cout(cout_8[28]),
    .sum(sum_8[28]));
  AL_FADD comp8_29 (
    .a(i8[29]),
    .b(sum_7[29]),
    .c(cout_8[28]),
    .cout(cout_8[29]),
    .sum(sum_8[29]));
  AL_FADD comp8_3 (
    .a(i8[3]),
    .b(sum_7[3]),
    .c(cout_8[2]),
    .cout(cout_8[3]),
    .sum(sum_8[3]));
  AL_FADD comp8_30 (
    .a(i8[30]),
    .b(sum_7[30]),
    .c(cout_8[29]),
    .cout(cout_8[30]),
    .sum(sum_8[30]));
  AL_FADD comp8_31 (
    .a(i8[31]),
    .b(sum_7[31]),
    .c(cout_8[30]),
    .cout(cout_8[31]),
    .sum(sum_8[31]));
  AL_FADD comp8_32 (
    .a(i8[32]),
    .b(sum_7[32]),
    .c(cout_8[31]),
    .cout(cout_8[32]),
    .sum(sum_8[32]));
  AL_FADD comp8_33 (
    .a(i8[33]),
    .b(sum_7[33]),
    .c(cout_8[32]),
    .cout(cout_8[33]),
    .sum(sum_8[33]));
  AL_FADD comp8_34 (
    .a(i8[34]),
    .b(sum_7[34]),
    .c(cout_8[33]),
    .cout(cout_8[34]),
    .sum(sum_8[34]));
  AL_FADD comp8_35 (
    .a(i8[35]),
    .b(sum_7[35]),
    .c(cout_8[34]),
    .cout(cout_8[35]),
    .sum(sum_8[35]));
  AL_FADD comp8_36 (
    .a(i8[36]),
    .b(sum_7[36]),
    .c(cout_8[35]),
    .cout(cout_8[36]),
    .sum(sum_8[36]));
  AL_FADD comp8_37 (
    .a(i8[37]),
    .b(sum_7[37]),
    .c(cout_8[36]),
    .cout(cout_8[37]),
    .sum(sum_8[37]));
  AL_FADD comp8_38 (
    .a(i8[38]),
    .b(sum_7[38]),
    .c(cout_8[37]),
    .cout(cout_8[38]),
    .sum(sum_8[38]));
  AL_FADD comp8_39 (
    .a(i8[39]),
    .b(sum_7[39]),
    .c(cout_8[38]),
    .cout(cout_8[39]),
    .sum(sum_8[39]));
  AL_FADD comp8_4 (
    .a(i8[4]),
    .b(sum_7[4]),
    .c(cout_8[3]),
    .cout(cout_8[4]),
    .sum(sum_8[4]));
  AL_FADD comp8_40 (
    .a(i8[40]),
    .b(sum_7[40]),
    .c(cout_8[39]),
    .cout(cout_8[40]),
    .sum(sum_8[40]));
  AL_FADD comp8_41 (
    .a(i8[41]),
    .b(sum_7[41]),
    .c(cout_8[40]),
    .cout(cout_8[41]),
    .sum(sum_8[41]));
  AL_FADD comp8_42 (
    .a(i8[42]),
    .b(sum_7[42]),
    .c(cout_8[41]),
    .cout(cout_8[42]),
    .sum(sum_8[42]));
  AL_FADD comp8_43 (
    .a(i8[43]),
    .b(sum_7[43]),
    .c(cout_8[42]),
    .cout(cout_8[43]),
    .sum(sum_8[43]));
  AL_FADD comp8_44 (
    .a(i8[44]),
    .b(sum_7[44]),
    .c(cout_8[43]),
    .cout(cout_8[44]),
    .sum(sum_8[44]));
  AL_FADD comp8_45 (
    .a(i8[45]),
    .b(sum_7[45]),
    .c(cout_8[44]),
    .cout(cout_8[45]),
    .sum(sum_8[45]));
  AL_FADD comp8_46 (
    .a(i8[46]),
    .b(sum_7[46]),
    .c(cout_8[45]),
    .cout(cout_8[46]),
    .sum(sum_8[46]));
  AL_FADD comp8_47 (
    .a(i8[47]),
    .b(sum_7[47]),
    .c(cout_8[46]),
    .cout(cout_8[47]),
    .sum(sum_8[47]));
  AL_FADD comp8_48 (
    .a(i8[48]),
    .b(sum_7[48]),
    .c(cout_8[47]),
    .cout(cout_8[48]),
    .sum(sum_8[48]));
  AL_FADD comp8_49 (
    .a(i8[49]),
    .b(sum_7[49]),
    .c(cout_8[48]),
    .cout(cout_8[49]),
    .sum(sum_8[49]));
  AL_FADD comp8_5 (
    .a(i8[5]),
    .b(sum_7[5]),
    .c(cout_8[4]),
    .cout(cout_8[5]),
    .sum(sum_8[5]));
  AL_FADD comp8_50 (
    .a(i8[50]),
    .b(sum_7[50]),
    .c(cout_8[49]),
    .cout(cout_8[50]),
    .sum(sum_8[50]));
  AL_FADD comp8_51 (
    .a(i8[51]),
    .b(sum_7[51]),
    .c(cout_8[50]),
    .cout(cout_8[51]),
    .sum(sum_8[51]));
  AL_FADD comp8_52 (
    .a(i8[52]),
    .b(sum_7[52]),
    .c(cout_8[51]),
    .cout(cout_8[52]),
    .sum(sum_8[52]));
  AL_FADD comp8_53 (
    .a(i8[53]),
    .b(sum_7[53]),
    .c(cout_8[52]),
    .cout(cout_8[53]),
    .sum(sum_8[53]));
  AL_FADD comp8_54 (
    .a(1'b0),
    .b(sum_7[54]),
    .c(cout_8[53]),
    .cout(cout_8[54]),
    .sum(sum_8[54]));
  AL_FADD comp8_55 (
    .a(1'b0),
    .b(sum_7[55]),
    .c(cout_8[54]),
    .cout(cout_8[55]),
    .sum(sum_8[55]));
  AL_FADD comp8_56 (
    .a(1'b0),
    .b(sum_7[56]),
    .c(cout_8[55]),
    .cout(cout_8[56]),
    .sum(sum_8[56]));
  AL_FADD comp8_57 (
    .a(1'b0),
    .b(sum_7[57]),
    .c(cout_8[56]),
    .cout(cout_8[57]),
    .sum(sum_8[57]));
  AL_FADD comp8_58 (
    .a(1'b0),
    .b(sum_7[58]),
    .c(cout_8[57]),
    .cout(cout_8[58]),
    .sum(sum_8[58]));
  AL_FADD comp8_59 (
    .a(1'b0),
    .b(sum_7[59]),
    .c(cout_8[58]),
    .cout(cout_8[59]),
    .sum(sum_8[59]));
  AL_FADD comp8_6 (
    .a(i8[6]),
    .b(sum_7[6]),
    .c(cout_8[5]),
    .cout(cout_8[6]),
    .sum(sum_8[6]));
  AL_FADD comp8_60 (
    .a(1'b0),
    .b(sum_7[60]),
    .c(cout_8[59]),
    .cout(cout_8[60]),
    .sum(sum_8[60]));
  AL_FADD comp8_61 (
    .a(1'b0),
    .b(sum_7[61]),
    .c(cout_8[60]),
    .cout(cout_8[61]),
    .sum(sum_8[61]));
  AL_FADD comp8_62 (
    .a(1'b0),
    .b(sum_7[62]),
    .c(cout_8[61]),
    .cout(cout_8[62]),
    .sum(sum_8[62]));
  AL_FADD comp8_63 (
    .a(1'b0),
    .b(sum_7[63]),
    .c(cout_8[62]),
    .cout(cout_8[63]),
    .sum(sum_8[63]));
  AL_FADD comp8_7 (
    .a(i8[7]),
    .b(sum_7[7]),
    .c(cout_8[6]),
    .cout(cout_8[7]),
    .sum(sum_8[7]));
  AL_FADD comp8_8 (
    .a(i8[8]),
    .b(sum_7[8]),
    .c(cout_8[7]),
    .cout(cout_8[8]),
    .sum(sum_8[8]));
  AL_FADD comp8_9 (
    .a(i8[9]),
    .b(sum_7[9]),
    .c(cout_8[8]),
    .cout(cout_8[9]),
    .sum(sum_8[9]));
  AL_FADD comp9_0 (
    .a(i9[0]),
    .b(sum_8[0]),
    .c(1'b0),
    .cout(cout_9[0]),
    .sum(sum_9[0]));
  AL_FADD comp9_1 (
    .a(i9[1]),
    .b(sum_8[1]),
    .c(cout_9[0]),
    .cout(cout_9[1]),
    .sum(sum_9[1]));
  AL_FADD comp9_10 (
    .a(i9[10]),
    .b(sum_8[10]),
    .c(cout_9[9]),
    .cout(cout_9[10]),
    .sum(sum_9[10]));
  AL_FADD comp9_11 (
    .a(i9[11]),
    .b(sum_8[11]),
    .c(cout_9[10]),
    .cout(cout_9[11]),
    .sum(sum_9[11]));
  AL_FADD comp9_12 (
    .a(i9[12]),
    .b(sum_8[12]),
    .c(cout_9[11]),
    .cout(cout_9[12]),
    .sum(sum_9[12]));
  AL_FADD comp9_13 (
    .a(i9[13]),
    .b(sum_8[13]),
    .c(cout_9[12]),
    .cout(cout_9[13]),
    .sum(sum_9[13]));
  AL_FADD comp9_14 (
    .a(i9[14]),
    .b(sum_8[14]),
    .c(cout_9[13]),
    .cout(cout_9[14]),
    .sum(sum_9[14]));
  AL_FADD comp9_15 (
    .a(i9[15]),
    .b(sum_8[15]),
    .c(cout_9[14]),
    .cout(cout_9[15]),
    .sum(sum_9[15]));
  AL_FADD comp9_16 (
    .a(i9[16]),
    .b(sum_8[16]),
    .c(cout_9[15]),
    .cout(cout_9[16]),
    .sum(sum_9[16]));
  AL_FADD comp9_17 (
    .a(i9[17]),
    .b(sum_8[17]),
    .c(cout_9[16]),
    .cout(cout_9[17]),
    .sum(sum_9[17]));
  AL_FADD comp9_18 (
    .a(i9[18]),
    .b(sum_8[18]),
    .c(cout_9[17]),
    .cout(cout_9[18]),
    .sum(sum_9[18]));
  AL_FADD comp9_19 (
    .a(i9[19]),
    .b(sum_8[19]),
    .c(cout_9[18]),
    .cout(cout_9[19]),
    .sum(sum_9[19]));
  AL_FADD comp9_2 (
    .a(i9[2]),
    .b(sum_8[2]),
    .c(cout_9[1]),
    .cout(cout_9[2]),
    .sum(sum_9[2]));
  AL_FADD comp9_20 (
    .a(i9[20]),
    .b(sum_8[20]),
    .c(cout_9[19]),
    .cout(cout_9[20]),
    .sum(sum_9[20]));
  AL_FADD comp9_21 (
    .a(i9[21]),
    .b(sum_8[21]),
    .c(cout_9[20]),
    .cout(cout_9[21]),
    .sum(sum_9[21]));
  AL_FADD comp9_22 (
    .a(i9[22]),
    .b(sum_8[22]),
    .c(cout_9[21]),
    .cout(cout_9[22]),
    .sum(sum_9[22]));
  AL_FADD comp9_23 (
    .a(i9[23]),
    .b(sum_8[23]),
    .c(cout_9[22]),
    .cout(cout_9[23]),
    .sum(sum_9[23]));
  AL_FADD comp9_24 (
    .a(i9[24]),
    .b(sum_8[24]),
    .c(cout_9[23]),
    .cout(cout_9[24]),
    .sum(sum_9[24]));
  AL_FADD comp9_25 (
    .a(i9[25]),
    .b(sum_8[25]),
    .c(cout_9[24]),
    .cout(cout_9[25]),
    .sum(sum_9[25]));
  AL_FADD comp9_26 (
    .a(i9[26]),
    .b(sum_8[26]),
    .c(cout_9[25]),
    .cout(cout_9[26]),
    .sum(sum_9[26]));
  AL_FADD comp9_27 (
    .a(i9[27]),
    .b(sum_8[27]),
    .c(cout_9[26]),
    .cout(cout_9[27]),
    .sum(sum_9[27]));
  AL_FADD comp9_28 (
    .a(i9[28]),
    .b(sum_8[28]),
    .c(cout_9[27]),
    .cout(cout_9[28]),
    .sum(sum_9[28]));
  AL_FADD comp9_29 (
    .a(i9[29]),
    .b(sum_8[29]),
    .c(cout_9[28]),
    .cout(cout_9[29]),
    .sum(sum_9[29]));
  AL_FADD comp9_3 (
    .a(i9[3]),
    .b(sum_8[3]),
    .c(cout_9[2]),
    .cout(cout_9[3]),
    .sum(sum_9[3]));
  AL_FADD comp9_30 (
    .a(i9[30]),
    .b(sum_8[30]),
    .c(cout_9[29]),
    .cout(cout_9[30]),
    .sum(sum_9[30]));
  AL_FADD comp9_31 (
    .a(i9[31]),
    .b(sum_8[31]),
    .c(cout_9[30]),
    .cout(cout_9[31]),
    .sum(sum_9[31]));
  AL_FADD comp9_32 (
    .a(i9[32]),
    .b(sum_8[32]),
    .c(cout_9[31]),
    .cout(cout_9[32]),
    .sum(sum_9[32]));
  AL_FADD comp9_33 (
    .a(i9[33]),
    .b(sum_8[33]),
    .c(cout_9[32]),
    .cout(cout_9[33]),
    .sum(sum_9[33]));
  AL_FADD comp9_34 (
    .a(i9[34]),
    .b(sum_8[34]),
    .c(cout_9[33]),
    .cout(cout_9[34]),
    .sum(sum_9[34]));
  AL_FADD comp9_35 (
    .a(i9[35]),
    .b(sum_8[35]),
    .c(cout_9[34]),
    .cout(cout_9[35]),
    .sum(sum_9[35]));
  AL_FADD comp9_36 (
    .a(i9[36]),
    .b(sum_8[36]),
    .c(cout_9[35]),
    .cout(cout_9[36]),
    .sum(sum_9[36]));
  AL_FADD comp9_37 (
    .a(i9[37]),
    .b(sum_8[37]),
    .c(cout_9[36]),
    .cout(cout_9[37]),
    .sum(sum_9[37]));
  AL_FADD comp9_38 (
    .a(i9[38]),
    .b(sum_8[38]),
    .c(cout_9[37]),
    .cout(cout_9[38]),
    .sum(sum_9[38]));
  AL_FADD comp9_39 (
    .a(i9[39]),
    .b(sum_8[39]),
    .c(cout_9[38]),
    .cout(cout_9[39]),
    .sum(sum_9[39]));
  AL_FADD comp9_4 (
    .a(i9[4]),
    .b(sum_8[4]),
    .c(cout_9[3]),
    .cout(cout_9[4]),
    .sum(sum_9[4]));
  AL_FADD comp9_40 (
    .a(i9[40]),
    .b(sum_8[40]),
    .c(cout_9[39]),
    .cout(cout_9[40]),
    .sum(sum_9[40]));
  AL_FADD comp9_41 (
    .a(i9[41]),
    .b(sum_8[41]),
    .c(cout_9[40]),
    .cout(cout_9[41]),
    .sum(sum_9[41]));
  AL_FADD comp9_42 (
    .a(i9[42]),
    .b(sum_8[42]),
    .c(cout_9[41]),
    .cout(cout_9[42]),
    .sum(sum_9[42]));
  AL_FADD comp9_43 (
    .a(i9[43]),
    .b(sum_8[43]),
    .c(cout_9[42]),
    .cout(cout_9[43]),
    .sum(sum_9[43]));
  AL_FADD comp9_44 (
    .a(i9[44]),
    .b(sum_8[44]),
    .c(cout_9[43]),
    .cout(cout_9[44]),
    .sum(sum_9[44]));
  AL_FADD comp9_45 (
    .a(i9[45]),
    .b(sum_8[45]),
    .c(cout_9[44]),
    .cout(cout_9[45]),
    .sum(sum_9[45]));
  AL_FADD comp9_46 (
    .a(i9[46]),
    .b(sum_8[46]),
    .c(cout_9[45]),
    .cout(cout_9[46]),
    .sum(sum_9[46]));
  AL_FADD comp9_47 (
    .a(i9[47]),
    .b(sum_8[47]),
    .c(cout_9[46]),
    .cout(cout_9[47]),
    .sum(sum_9[47]));
  AL_FADD comp9_48 (
    .a(i9[48]),
    .b(sum_8[48]),
    .c(cout_9[47]),
    .cout(cout_9[48]),
    .sum(sum_9[48]));
  AL_FADD comp9_49 (
    .a(i9[49]),
    .b(sum_8[49]),
    .c(cout_9[48]),
    .cout(cout_9[49]),
    .sum(sum_9[49]));
  AL_FADD comp9_5 (
    .a(i9[5]),
    .b(sum_8[5]),
    .c(cout_9[4]),
    .cout(cout_9[5]),
    .sum(sum_9[5]));
  AL_FADD comp9_50 (
    .a(i9[50]),
    .b(sum_8[50]),
    .c(cout_9[49]),
    .cout(cout_9[50]),
    .sum(sum_9[50]));
  AL_FADD comp9_51 (
    .a(i9[51]),
    .b(sum_8[51]),
    .c(cout_9[50]),
    .cout(cout_9[51]),
    .sum(sum_9[51]));
  AL_FADD comp9_52 (
    .a(i9[52]),
    .b(sum_8[52]),
    .c(cout_9[51]),
    .cout(cout_9[52]),
    .sum(sum_9[52]));
  AL_FADD comp9_53 (
    .a(1'b0),
    .b(sum_8[53]),
    .c(cout_9[52]),
    .cout(cout_9[53]),
    .sum(sum_9[53]));
  AL_FADD comp9_54 (
    .a(1'b0),
    .b(sum_8[54]),
    .c(cout_9[53]),
    .cout(cout_9[54]),
    .sum(sum_9[54]));
  AL_FADD comp9_55 (
    .a(1'b0),
    .b(sum_8[55]),
    .c(cout_9[54]),
    .cout(cout_9[55]),
    .sum(sum_9[55]));
  AL_FADD comp9_56 (
    .a(1'b0),
    .b(sum_8[56]),
    .c(cout_9[55]),
    .cout(cout_9[56]),
    .sum(sum_9[56]));
  AL_FADD comp9_57 (
    .a(1'b0),
    .b(sum_8[57]),
    .c(cout_9[56]),
    .cout(cout_9[57]),
    .sum(sum_9[57]));
  AL_FADD comp9_58 (
    .a(1'b0),
    .b(sum_8[58]),
    .c(cout_9[57]),
    .cout(cout_9[58]),
    .sum(sum_9[58]));
  AL_FADD comp9_59 (
    .a(1'b0),
    .b(sum_8[59]),
    .c(cout_9[58]),
    .cout(cout_9[59]),
    .sum(sum_9[59]));
  AL_FADD comp9_6 (
    .a(i9[6]),
    .b(sum_8[6]),
    .c(cout_9[5]),
    .cout(cout_9[6]),
    .sum(sum_9[6]));
  AL_FADD comp9_60 (
    .a(1'b0),
    .b(sum_8[60]),
    .c(cout_9[59]),
    .cout(cout_9[60]),
    .sum(sum_9[60]));
  AL_FADD comp9_61 (
    .a(1'b0),
    .b(sum_8[61]),
    .c(cout_9[60]),
    .cout(cout_9[61]),
    .sum(sum_9[61]));
  AL_FADD comp9_62 (
    .a(1'b0),
    .b(sum_8[62]),
    .c(cout_9[61]),
    .cout(cout_9[62]),
    .sum(sum_9[62]));
  AL_FADD comp9_63 (
    .a(1'b0),
    .b(sum_8[63]),
    .c(cout_9[62]),
    .cout(cout_9[63]),
    .sum(sum_9[63]));
  AL_FADD comp9_7 (
    .a(i9[7]),
    .b(sum_8[7]),
    .c(cout_9[6]),
    .cout(cout_9[7]),
    .sum(sum_9[7]));
  AL_FADD comp9_8 (
    .a(i9[8]),
    .b(sum_8[8]),
    .c(cout_9[7]),
    .cout(cout_9[8]),
    .sum(sum_9[8]));
  AL_FADD comp9_9 (
    .a(i9[9]),
    .b(sum_8[9]),
    .c(cout_9[8]),
    .cout(cout_9[9]),
    .sum(sum_9[9]));
  not inv_b31_0 (net_nb31_0, i31[0]);
  not inv_b31_1 (net_nb31_1, i31[1]);
  not inv_b31_10 (net_nb31_10, i31[10]);
  not inv_b31_11 (net_nb31_11, i31[11]);
  not inv_b31_12 (net_nb31_12, i31[12]);
  not inv_b31_13 (net_nb31_13, i31[13]);
  not inv_b31_14 (net_nb31_14, i31[14]);
  not inv_b31_15 (net_nb31_15, i31[15]);
  not inv_b31_16 (net_nb31_16, i31[16]);
  not inv_b31_17 (net_nb31_17, i31[17]);
  not inv_b31_18 (net_nb31_18, i31[18]);
  not inv_b31_19 (net_nb31_19, i31[19]);
  not inv_b31_2 (net_nb31_2, i31[2]);
  not inv_b31_20 (net_nb31_20, i31[20]);
  not inv_b31_21 (net_nb31_21, i31[21]);
  not inv_b31_22 (net_nb31_22, i31[22]);
  not inv_b31_23 (net_nb31_23, i31[23]);
  not inv_b31_24 (net_nb31_24, i31[24]);
  not inv_b31_25 (net_nb31_25, i31[25]);
  not inv_b31_26 (net_nb31_26, i31[26]);
  not inv_b31_27 (net_nb31_27, i31[27]);
  not inv_b31_28 (net_nb31_28, i31[28]);
  not inv_b31_29 (net_nb31_29, i31[29]);
  not inv_b31_3 (net_nb31_3, i31[3]);
  not inv_b31_30 (net_nb31_30, i31[30]);
  not inv_b31_31 (net_nb31_31, i31[31]);
  not inv_b31_32 (net_nb31_32, i31[32]);
  not inv_b31_33 (net_nb31_33, i31[33]);
  not inv_b31_34 (net_nb31_34, i31[34]);
  not inv_b31_35 (net_nb31_35, i31[35]);
  not inv_b31_36 (net_nb31_36, i31[36]);
  not inv_b31_37 (net_nb31_37, i31[37]);
  not inv_b31_38 (net_nb31_38, i31[38]);
  not inv_b31_39 (net_nb31_39, i31[39]);
  not inv_b31_4 (net_nb31_4, i31[4]);
  not inv_b31_40 (net_nb31_40, i31[40]);
  not inv_b31_41 (net_nb31_41, i31[41]);
  not inv_b31_42 (net_nb31_42, i31[42]);
  not inv_b31_43 (net_nb31_43, i31[43]);
  not inv_b31_44 (net_nb31_44, i31[44]);
  not inv_b31_45 (net_nb31_45, i31[45]);
  not inv_b31_46 (net_nb31_46, i31[46]);
  not inv_b31_47 (net_nb31_47, i31[47]);
  not inv_b31_48 (net_nb31_48, i31[48]);
  not inv_b31_49 (net_nb31_49, i31[49]);
  not inv_b31_5 (net_nb31_5, i31[5]);
  not inv_b31_50 (net_nb31_50, i31[50]);
  not inv_b31_51 (net_nb31_51, i31[51]);
  not inv_b31_52 (net_nb31_52, i31[52]);
  not inv_b31_53 (net_nb31_53, i31[53]);
  not inv_b31_54 (net_nb31_54, i31[54]);
  not inv_b31_55 (net_nb31_55, i31[55]);
  not inv_b31_56 (net_nb31_56, i31[56]);
  not inv_b31_57 (net_nb31_57, i31[57]);
  not inv_b31_58 (net_nb31_58, i31[58]);
  not inv_b31_59 (net_nb31_59, i31[59]);
  not inv_b31_6 (net_nb31_6, i31[6]);
  not inv_b31_60 (net_nb31_60, i31[60]);
  not inv_b31_61 (net_nb31_61, i31[61]);
  not inv_b31_62 (net_nb31_62, i31[62]);
  not inv_b31_63 (net_nb31_63, 1'b0);
  not inv_b31_7 (net_nb31_7, i31[7]);
  not inv_b31_8 (net_nb31_8, i31[8]);
  not inv_b31_9 (net_nb31_9, i31[9]);
  not inv_b32_0 (net_nb32_0, i32[0]);
  not inv_b32_1 (net_nb32_1, i32[1]);
  not inv_b32_10 (net_nb32_10, i32[10]);
  not inv_b32_11 (net_nb32_11, i32[11]);
  not inv_b32_12 (net_nb32_12, i32[12]);
  not inv_b32_13 (net_nb32_13, i32[13]);
  not inv_b32_14 (net_nb32_14, i32[14]);
  not inv_b32_15 (net_nb32_15, i32[15]);
  not inv_b32_16 (net_nb32_16, i32[16]);
  not inv_b32_17 (net_nb32_17, i32[17]);
  not inv_b32_18 (net_nb32_18, i32[18]);
  not inv_b32_19 (net_nb32_19, i32[19]);
  not inv_b32_2 (net_nb32_2, i32[2]);
  not inv_b32_20 (net_nb32_20, i32[20]);
  not inv_b32_21 (net_nb32_21, i32[21]);
  not inv_b32_22 (net_nb32_22, i32[22]);
  not inv_b32_23 (net_nb32_23, i32[23]);
  not inv_b32_24 (net_nb32_24, i32[24]);
  not inv_b32_25 (net_nb32_25, i32[25]);
  not inv_b32_26 (net_nb32_26, i32[26]);
  not inv_b32_27 (net_nb32_27, i32[27]);
  not inv_b32_28 (net_nb32_28, i32[28]);
  not inv_b32_29 (net_nb32_29, i32[29]);
  not inv_b32_3 (net_nb32_3, i32[3]);
  not inv_b32_30 (net_nb32_30, i32[30]);
  not inv_b32_31 (net_nb32_31, i32[31]);
  not inv_b32_32 (net_nb32_32, i32[32]);
  not inv_b32_33 (net_nb32_33, i32[33]);
  not inv_b32_34 (net_nb32_34, i32[34]);
  not inv_b32_35 (net_nb32_35, i32[35]);
  not inv_b32_36 (net_nb32_36, i32[36]);
  not inv_b32_37 (net_nb32_37, i32[37]);
  not inv_b32_38 (net_nb32_38, i32[38]);
  not inv_b32_39 (net_nb32_39, i32[39]);
  not inv_b32_4 (net_nb32_4, i32[4]);
  not inv_b32_40 (net_nb32_40, i32[40]);
  not inv_b32_41 (net_nb32_41, i32[41]);
  not inv_b32_42 (net_nb32_42, i32[42]);
  not inv_b32_43 (net_nb32_43, i32[43]);
  not inv_b32_44 (net_nb32_44, i32[44]);
  not inv_b32_45 (net_nb32_45, i32[45]);
  not inv_b32_46 (net_nb32_46, i32[46]);
  not inv_b32_47 (net_nb32_47, i32[47]);
  not inv_b32_48 (net_nb32_48, i32[48]);
  not inv_b32_49 (net_nb32_49, i32[49]);
  not inv_b32_5 (net_nb32_5, i32[5]);
  not inv_b32_50 (net_nb32_50, i32[50]);
  not inv_b32_51 (net_nb32_51, i32[51]);
  not inv_b32_52 (net_nb32_52, i32[52]);
  not inv_b32_53 (net_nb32_53, i32[53]);
  not inv_b32_54 (net_nb32_54, i32[54]);
  not inv_b32_55 (net_nb32_55, i32[55]);
  not inv_b32_56 (net_nb32_56, i32[56]);
  not inv_b32_57 (net_nb32_57, i32[57]);
  not inv_b32_58 (net_nb32_58, i32[58]);
  not inv_b32_59 (net_nb32_59, i32[59]);
  not inv_b32_6 (net_nb32_6, i32[6]);
  not inv_b32_60 (net_nb32_60, i32[60]);
  not inv_b32_61 (net_nb32_61, i32[61]);
  not inv_b32_62 (net_nb32_62, i32[62]);
  not inv_b32_63 (net_nb32_63, 1'b0);
  not inv_b32_7 (net_nb32_7, i32[7]);
  not inv_b32_8 (net_nb32_8, i32[8]);
  not inv_b32_9 (net_nb32_9, i32[9]);
  not inv_cout31_63 (net_ncout31_63, cout_31[63]);
  not inv_cout32_63 (net_ncout32_63, cout_32[63]);

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  // synthesis translate_off
  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end
  // synthesis translate_on

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

module AL_FADD
  (
  input a,
  input b,
  input c,
  output sum,
  output cout
  );

  wire prop;
  wire not_prop;
  wire sel_i0;
  wire sel_i1;

  xor u0 (prop, a, b);
  xor u1 (sum, prop, c);
  not u2 (not_prop, prop);
  and u3 (sel_i1, prop, c);
  and u4 (sel_i0, not_prop, a);
  or  u5 (cout, sel_i0, sel_i1);

endmodule

module AL_LATCH
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  // synthesis translate_off
  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end
  // synthesis translate_on

  always @(reset or set or clk or d)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else if (clk)
      q <= d;
  end

endmodule

