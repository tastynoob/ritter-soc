// Verilog netlist created by TD v5.0.38657
// Thu Jan 27 23:49:07 2022

`timescale 1ns / 1ps
module TEST_TOP  // ../simulation/tb.v(6)
  (
  );




endmodule 

