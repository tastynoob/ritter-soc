// Verilog netlist created by TD v5.0.38657
// Fri Feb 25 00:19:08 2022

`timescale 1ns / 1ps
module SOC_TOP  // ../RTL/soc_top/soc_top.v(5)
  (
  i_clk,
  i_io_rx,
  i_rstn,
  o_io_tx
  );

  input i_clk;  // ../RTL/soc_top/soc_top.v(6)
  input i_io_rx;  // ../RTL/soc_top/soc_top.v(9)
  input i_rstn;  // ../RTL/soc_top/soc_top.v(7)
  output o_io_tx;  // ../RTL/soc_top/soc_top.v(10)

  wire [31:0] periph_addr;  // ../RTL/soc_top/soc_top.v(40)
  wire [31:0] periph_rdata;  // ../RTL/soc_top/soc_top.v(44)
  wire [31:0] periph_wdata;  // ../RTL/soc_top/soc_top.v(43)
  wire [31:0] \u_PERIPH_TOP/timer_ribs_rdata ;  // ../RTL/periph/periph_top.v(65)
  wire [1:0] \u_PERIPH_TOP/u_SLAVE_SEL/sel_tag ;  // ../RTL/core/rib.v(78)
  wire [7:0] \u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id ;  // ../RTL/core/rib.v(113)
  wire [63:0] \u_PERIPH_TOP/u_TIMER2RIB/n12 ;
  wire [63:0] \u_PERIPH_TOP/u_TIMER2RIB/n13 ;
  wire [63:0] \u_PERIPH_TOP/u_TIMER2RIB/n14 ;
  wire [63:0] \u_PERIPH_TOP/u_TIMER2RIB/n18 ;
  wire [63:0] \u_PERIPH_TOP/u_TIMER2RIB/timer_cnt ;  // ../RTL/periph/timer2rib.v(30)
  wire [31:0] \u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl ;  // ../RTL/periph/timer2rib.v(29)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/rx_data ;  // ../RTL/periph/usart2rib.v(34)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/tx_buffer ;  // ../RTL/periph/usart2rib.v(30)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 ;  // al_ip/usart_gate.v(45)
  wire [5:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 ;  // al_ip/usart_gate.v(46)
  wire [5:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 ;  // al_ip/usart_gate.v(49)
  wire [5:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 ;  // al_ip/usart_gate.v(48)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 ;  // al_ip/usart_gate.v(47)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 ;  // al_ip/usart_gate.v(50)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 ;  // al_ip/usart_gate.v(52)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 ;  // al_ip/usart_gate.v(51)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 ;  // al_ip/usart_gate.v(55)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 ;  // al_ip/usart_gate.v(56)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 ;  // al_ip/usart_gate.v(57)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 ;  // al_ip/usart_gate.v(60)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 ;  // al_ip/usart_gate.v(59)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 ;  // al_ip/usart_gate.v(58)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 ;  // al_ip/usart_gate.v(61)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 ;  // al_ip/usart_gate.v(67)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A68B0 ;  // al_ip/usart_gate.v(69)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A7020 ;  // al_ip/usart_gate.v(68)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 ;  // al_ip/usart_gate.v(70)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 ;  // al_ip/usart_gate.v(71)
  wire [2:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 ;  // al_ip/usart_gate.v(72)
  wire [3:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 ;  // al_ip/usart_gate.v(73)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 ;  // al_ip/usart_gate.v(74)
  wire [7:0] \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 ;  // al_ip/usart_gate.v(75)
  wire [31:0] \u_PERIPH_TOP/usart_rib_rdata ;  // ../RTL/periph/periph_top.v(35)
  wire [4:0] \u_internal_reset/synch_regs_q ;  // ../RTL/core/reset.v(13)
  wire _al_u582_o;
  wire _al_u583_o;
  wire _al_u585_o;
  wire _al_u587_o;
  wire _al_u589_o;
  wire _al_u591_o;
  wire _al_u593_o;
  wire _al_u595_o;
  wire _al_u597_o;
  wire _al_u599_o;
  wire _al_u601_o;
  wire _al_u603_o;
  wire _al_u605_o;
  wire _al_u607_o;
  wire _al_u609_o;
  wire _al_u611_o;
  wire _al_u613_o;
  wire _al_u615_o;
  wire _al_u617_o;
  wire _al_u619_o;
  wire _al_u621_o;
  wire _al_u623_o;
  wire _al_u625_o;
  wire _al_u627_o;
  wire _al_u629_o;
  wire _al_u631_o;
  wire _al_u633_o;
  wire _al_u635_o;
  wire _al_u637_o;
  wire _al_u639_o;
  wire _al_u641_o;
  wire _al_u643_o;
  wire _al_u645_o;
  wire _al_u647_o;
  wire _al_u649_o;
  wire _al_u651_o;
  wire _al_u653_o;
  wire _al_u655_o;
  wire _al_u657_o;
  wire _al_u659_o;
  wire _al_u661_o;
  wire _al_u663_o;
  wire _al_u664_o;
  wire _al_u672_o;
  wire _al_u673_o;
  wire _al_u674_o;
  wire _al_u773_o;
  wire _al_u774_o;
  wire _al_u776_o;
  wire clk_84mhz;  // ../RTL/soc_top/soc_top.v(16)
  wire clk_84mhz_keep;
  wire extlock;  // ../RTL/soc_top/soc_top.v(15)
  wire i_clk_pad;  // ../RTL/soc_top/soc_top.v(6)
  wire i_io_rx_pad;  // ../RTL/soc_top/soc_top.v(9)
  wire i_rstn_pad;  // ../RTL/soc_top/soc_top.v(7)
  wire n0;
  wire n1;
  wire o_io_tx_pad;  // ../RTL/soc_top/soc_top.v(10)
  wire periph_req;  // ../RTL/soc_top/soc_top.v(45)
  wire periph_wrcs;  // ../RTL/soc_top/soc_top.v(41)
  wire reset;  // ../RTL/soc_top/soc_top.v(31)
  wire \u_PERIPH_TOP/timer_ribs_req ;  // ../RTL/periph/periph_top.v(66)
  wire \u_PERIPH_TOP/timer_ribs_rsp ;  // ../RTL/periph/periph_top.v(68)
  wire \u_PERIPH_TOP/u_SLAVE_SEL/default_cs ;  // ../RTL/core/rib.v(112)
  wire \u_PERIPH_TOP/u_SLAVE_SEL/handshake_rdy_last ;  // ../RTL/core/rib.v(117)
  wire \u_PERIPH_TOP/u_SLAVE_SEL/n0 ;
  wire \u_PERIPH_TOP/u_SLAVE_SEL/n1 ;
  wire \u_PERIPH_TOP/u_SLAVE_SEL/n3 ;
  wire \u_PERIPH_TOP/u_SLAVE_SEL/n6 ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c11 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c15 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c19 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c23 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c27 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c3 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c31 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c35 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c39 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c43 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c47 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c51 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c55 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c59 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c63 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/add0/c7 ;  // ../RTL/periph/timer2rib.v(73)
  wire \u_PERIPH_TOP/u_TIMER2RIB/mux3_b0_sel_is_3_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_8_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b10_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b11_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b12_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b13_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b14_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b15_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b16_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b17_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b18_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b19_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b1_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b20_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b21_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b22_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b23_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b24_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b25_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b26_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b27_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b28_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b29_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b2_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b30_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b31_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b3_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b4_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b5_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b6_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b7_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b8_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel1_b9_var_o ;
  wire \u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/n16 ;
  wire \u_PERIPH_TOP/u_USART2RIB/rx_err ;  // ../RTL/periph/usart2rib.v(35)
  wire \u_PERIPH_TOP/u_USART2RIB/rx_vld ;  // ../RTL/periph/usart2rib.v(33)
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b0_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b1_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b2_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b3_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b4_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b5_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b6_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/sel0_b7_var_o ;
  wire \u_PERIPH_TOP/u_USART2RIB/tx_en ;  // ../RTL/periph/usart2rib.v(37)
  wire \u_PERIPH_TOP/u_USART2RIB/tx_rdy ;  // ../RTL/periph/usart2rib.v(36)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533120 ;  // al_ip/usart_gate.v(160)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5335F0 ;  // al_ip/usart_gate.v(158)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533EE0 ;  // al_ip/usart_gate.v(168)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534250 ;  // al_ip/usart_gate.v(181)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534510 ;  // al_ip/usart_gate.v(164)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534880 ;  // al_ip/usart_gate.v(162)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534B40 ;  // al_ip/usart_gate.v(175)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534BF0 ;  // al_ip/usart_gate.v(177)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535380 ;  // al_ip/usart_gate.v(166)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535430 ;  // al_ip/usart_gate.v(170)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535590 ;  // al_ip/usart_gate.v(172)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535640 ;  // al_ip/usart_gate.v(179)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A340 ;  // al_ip/usart_gate.v(200)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A550 ;  // al_ip/usart_gate.v(199)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A550340 ;  // al_ip/usart_gate.v(53)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ;  // al_ip/usart_gate.v(213)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ;  // al_ip/usart_gate.v(214)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E4A0 ;  // al_ip/usart_gate.v(144)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E600 ;  // al_ip/usart_gate.v(148)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82ECE0 ;  // al_ip/usart_gate.v(142)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FB50 ;  // al_ip/usart_gate.v(146)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FCB0 ;  // al_ip/usart_gate.v(150)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830390 ;  // al_ip/usart_gate.v(152)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830C80 ;  // al_ip/usart_gate.v(156)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ;  // al_ip/usart_gate.v(154)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A832AC0 ;  // al_ip/usart_gate.v(183)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A832EE0 ;  // al_ip/usart_gate.v(155)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ;  // al_ip/usart_gate.v(184)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ;  // al_ip/usart_gate.v(187)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C9110 ;  // al_ip/usart_gate.v(186)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C93D0 ;  // al_ip/usart_gate.v(188)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C95E0 ;  // al_ip/usart_gate.v(185)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB2C0 ;  // al_ip/usart_gate.v(189)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB420 ;  // al_ip/usart_gate.v(190)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB6E0 ;  // al_ip/usart_gate.v(192)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB790 ;  // al_ip/usart_gate.v(196)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB840 ;  // al_ip/usart_gate.v(191)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CBF20 ;  // al_ip/usart_gate.v(197)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CC810 ;  // al_ip/usart_gate.v(198)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCA20 ;  // al_ip/usart_gate.v(195)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCD90 ;  // al_ip/usart_gate.v(193)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD470 ;  // al_ip/usart_gate.v(194)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD890 ;  // al_ip/usart_gate.v(201)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ;  // al_ip/usart_gate.v(202)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2010 ;  // al_ip/usart_gate.v(204)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2F30 ;  // al_ip/usart_gate.v(203)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D3FB0 ;  // al_ip/usart_gate.v(211)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4320 ;  // al_ip/usart_gate.v(205)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4480 ;  // al_ip/usart_gate.v(209)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4C10 ;  // al_ip/usart_gate.v(207)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D50E0 ;  // al_ip/usart_gate.v(206)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5A80 ;  // al_ip/usart_gate.v(210)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5B30 ;  // al_ip/usart_gate.v(212)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5BE0 ;  // al_ip/usart_gate.v(208)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5BBF0 ;  // al_ip/usart_gate.v(54)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5D780 ;  // al_ip/usart_gate.v(62)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5F070 ;  // al_ip/usart_gate.v(63)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA60730 ;  // al_ip/usart_gate.v(64)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA63600 ;  // al_ip/usart_gate.v(65)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9D8A0 ;  // al_ip/usart_gate.v(139)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9D950 ;  // al_ip/usart_gate.v(80)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DA00 ;  // al_ip/usart_gate.v(135)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DAB0 ;  // al_ip/usart_gate.v(118)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DB60 ;  // al_ip/usart_gate.v(119)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DC10 ;  // al_ip/usart_gate.v(126)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DCC0 ;  // al_ip/usart_gate.v(136)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ;  // al_ip/usart_gate.v(121)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DE20 ;  // al_ip/usart_gate.v(76)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DED0 ;  // al_ip/usart_gate.v(78)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DF80 ;  // al_ip/usart_gate.v(92)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ;  // al_ip/usart_gate.v(96)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E0E0 ;  // al_ip/usart_gate.v(97)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E190 ;  // al_ip/usart_gate.v(101)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E240 ;  // al_ip/usart_gate.v(87)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ;  // al_ip/usart_gate.v(127)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E500 ;  // al_ip/usart_gate.v(116)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ;  // al_ip/usart_gate.v(128)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E710 ;  // al_ip/usart_gate.v(138)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E7C0 ;  // al_ip/usart_gate.v(91)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ;  // al_ip/usart_gate.v(79)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E920 ;  // al_ip/usart_gate.v(93)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E9D0 ;  // al_ip/usart_gate.v(103)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EA80 ;  // al_ip/usart_gate.v(102)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EB30 ;  // al_ip/usart_gate.v(104)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EBE0 ;  // al_ip/usart_gate.v(105)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EC90 ;  // al_ip/usart_gate.v(106)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EDF0 ;  // al_ip/usart_gate.v(140)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EEA0 ;  // al_ip/usart_gate.v(107)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EF50 ;  // al_ip/usart_gate.v(108)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F000 ;  // al_ip/usart_gate.v(89)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ;  // al_ip/usart_gate.v(134)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F160 ;  // al_ip/usart_gate.v(125)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F210 ;  // al_ip/usart_gate.v(122)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ;  // al_ip/usart_gate.v(77)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F370 ;  // al_ip/usart_gate.v(81)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F420 ;  // al_ip/usart_gate.v(123)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F4D0 ;  // al_ip/usart_gate.v(84)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F580 ;  // al_ip/usart_gate.v(131)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F630 ;  // al_ip/usart_gate.v(85)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F6E0 ;  // al_ip/usart_gate.v(94)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F790 ;  // al_ip/usart_gate.v(98)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ;  // al_ip/usart_gate.v(124)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F8F0 ;  // al_ip/usart_gate.v(82)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F9A0 ;  // al_ip/usart_gate.v(88)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FA50 ;  // al_ip/usart_gate.v(83)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FB00 ;  // al_ip/usart_gate.v(90)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ;  // al_ip/usart_gate.v(117)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FC60 ;  // al_ip/usart_gate.v(95)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FD10 ;  // al_ip/usart_gate.v(99)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FDC0 ;  // al_ip/usart_gate.v(100)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FF20 ;  // al_ip/usart_gate.v(132)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FFD0 ;  // al_ip/usart_gate.v(129)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0080 ;  // al_ip/usart_gate.v(133)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA01E0 ;  // al_ip/usart_gate.v(137)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0290 ;  // al_ip/usart_gate.v(130)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0340 ;  // al_ip/usart_gate.v(86)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA03F0 ;  // al_ip/usart_gate.v(120)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0760 ;  // al_ip/usart_gate.v(115)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0A20 ;  // al_ip/usart_gate.v(114)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1100 ;  // al_ip/usart_gate.v(110)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1940 ;  // al_ip/usart_gate.v(112)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1AA0 ;  // al_ip/usart_gate.v(109)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1F70 ;  // al_ip/usart_gate.v(113)
  wire \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA22E0 ;  // al_ip/usart_gate.v(111)
  wire \u_PERIPH_TOP/usart_rib_req ;  // ../RTL/periph/periph_top.v(36)
  wire \u_PERIPH_TOP/usart_rib_rsp ;  // ../RTL/periph/periph_top.v(38)
  wire \u_pll/clk0_buf ;  // al_ip/pll.v(32)

  EG_PHY_PAD #(
    //.HYSTERESIS("OFF"),
    //.LOCATION("K14"),
    //.PCICLAMP("OFF"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u539 (
    .ipad(i_clk),
    .di(i_clk_pad));  // ../RTL/soc_top/soc_top.v(6)
  EG_PHY_PAD #(
    //.CLKSRC("CLK"),
    //.HYSTERESIS("OFF"),
    //.LOCATION("L12"),
    //.PCICLAMP("OFF"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .SRMODE("ASYNC"),
    .TSMUX("1"))
    _al_u540 (
    .ipad(i_io_rx),
    .di(i_io_rx_pad));  // ../RTL/soc_top/soc_top.v(9)
  EG_PHY_PAD #(
    //.HYSTERESIS("OFF"),
    //.LOCATION("K16"),
    //.PCICLAMP("OFF"),
    //.PULLMODE("PULLUP"),
    .IOTYPE("LVCMOS25"),
    .MODE("IN"),
    .TSMUX("1"))
    _al_u541 (
    .ipad(i_rstn),
    .di(i_rstn_pad));  // ../RTL/soc_top/soc_top.v(7)
  EG_PHY_PAD #(
    //.LOCATION("J11"),
    //.PCICLAMP("OFF"),
    //.PULLMODE("NONE"),
    //.SLEWRATE("SLOW"),
    .DRIVE("8"),
    .IOTYPE("LVCMOS25"),
    .MODE("OUT"),
    .TSMUX("0"))
    _al_u542 (
    .do({open_n52,open_n53,open_n54,o_io_tx_pad}),
    .opad(o_io_tx));  // ../RTL/soc_top/soc_top.v(10)
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u547 (
    .a(\u_PERIPH_TOP/timer_ribs_rsp ),
    .b(\u_PERIPH_TOP/usart_rib_rsp ),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u548 (
    .a(i_rstn_pad),
    .b(extlock),
    .o(n1));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u549 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/n1 ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/handshake_rdy_last ),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/n6 ));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h5140))
    _al_u550 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .o(periph_rdata[0]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h5140))
    _al_u551 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .o(periph_rdata[1]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h5140))
    _al_u552 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .o(periph_rdata[2]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h5140))
    _al_u553 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .o(periph_rdata[3]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h5140))
    _al_u554 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .o(periph_rdata[4]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h5140))
    _al_u555 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .o(periph_rdata[5]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h5140))
    _al_u556 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .o(periph_rdata[6]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'h5140))
    _al_u557 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .o(periph_rdata[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u558 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .o(periph_rdata[9]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u559 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .o(periph_rdata[8]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u560 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .o(periph_rdata[31]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u561 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .o(periph_rdata[30]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u562 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .o(periph_rdata[29]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u563 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .o(periph_rdata[28]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u564 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .o(periph_rdata[27]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u565 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .o(periph_rdata[26]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u566 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .o(periph_rdata[25]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u567 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .o(periph_rdata[24]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u568 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .o(periph_rdata[23]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u569 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .o(periph_rdata[22]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u570 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .o(periph_rdata[21]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u571 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .o(periph_rdata[20]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u572 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .o(periph_rdata[19]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u573 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .o(periph_rdata[18]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u574 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .o(periph_rdata[17]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u575 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .o(periph_rdata[16]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u576 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .o(periph_rdata[15]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u577 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .o(periph_rdata[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u578 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .o(periph_rdata[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u579 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .o(periph_rdata[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u580 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .o(periph_rdata[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u581 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]),
    .c(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .o(periph_rdata[10]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u582 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .o(_al_u582_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u583 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [1]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .o(_al_u583_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u584 (
    .a(_al_u583_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [33]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b1_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u585 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [10]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .o(_al_u585_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u586 (
    .a(_al_u585_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [42]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [10]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b10_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u587 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [11]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .o(_al_u587_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u588 (
    .a(_al_u587_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [43]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [11]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b11_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u589 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [12]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .o(_al_u589_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u590 (
    .a(_al_u589_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [44]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [12]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b12_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u591 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [13]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .o(_al_u591_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u592 (
    .a(_al_u591_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [45]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [13]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b13_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u593 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [14]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .o(_al_u593_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u594 (
    .a(_al_u593_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [46]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [14]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b14_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u595 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [15]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .o(_al_u595_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u596 (
    .a(_al_u595_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [47]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [15]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b15_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u597 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [16]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .o(_al_u597_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u598 (
    .a(_al_u597_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [48]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [16]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b16_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u599 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [17]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .o(_al_u599_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u600 (
    .a(_al_u599_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [49]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [17]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b17_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u601 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [18]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .o(_al_u601_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u602 (
    .a(_al_u601_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [50]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [18]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b18_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u603 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [19]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .o(_al_u603_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u604 (
    .a(_al_u603_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [51]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [19]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b19_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u605 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [2]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .o(_al_u605_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u606 (
    .a(_al_u605_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [34]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [2]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b2_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u607 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [20]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .o(_al_u607_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u608 (
    .a(_al_u607_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [52]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [20]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b20_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u609 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [21]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .o(_al_u609_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u610 (
    .a(_al_u609_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [53]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [21]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b21_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u611 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [22]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .o(_al_u611_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u612 (
    .a(_al_u611_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [54]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [22]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b22_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u613 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [23]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .o(_al_u613_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u614 (
    .a(_al_u613_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [55]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [23]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b23_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u615 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [24]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .o(_al_u615_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u616 (
    .a(_al_u615_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [56]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [24]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b24_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u617 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [25]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .o(_al_u617_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u618 (
    .a(_al_u617_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [57]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [25]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b25_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u619 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [26]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .o(_al_u619_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u620 (
    .a(_al_u619_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [58]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [26]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b26_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u621 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [27]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .o(_al_u621_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u622 (
    .a(_al_u621_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [59]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [27]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b27_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u623 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [28]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .o(_al_u623_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u624 (
    .a(_al_u623_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [60]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [28]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b28_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u625 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [29]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .o(_al_u625_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u626 (
    .a(_al_u625_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [61]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [29]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b29_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u627 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [3]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .o(_al_u627_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u628 (
    .a(_al_u627_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [35]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [3]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b3_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u629 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [30]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .o(_al_u629_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u630 (
    .a(_al_u629_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [62]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [30]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b30_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u631 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [31]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .o(_al_u631_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u632 (
    .a(_al_u631_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [63]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [31]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b31_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u633 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [4]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .o(_al_u633_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u634 (
    .a(_al_u633_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [36]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [4]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b4_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u635 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [5]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .o(_al_u635_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u636 (
    .a(_al_u635_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [37]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [5]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b5_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u637 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [6]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .o(_al_u637_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u638 (
    .a(_al_u637_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [38]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [6]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b6_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u639 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [7]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .o(_al_u639_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u640 (
    .a(_al_u639_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [39]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [7]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b7_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u641 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [8]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .o(_al_u641_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u642 (
    .a(_al_u641_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [40]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [8]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b8_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((C*A)*~(D)*~(B)+(C*A)*D*~(B)+~((C*A))*D*B+(C*A)*D*B)"),
    .INIT(16'h13df))
    _al_u643 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [9]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .o(_al_u643_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u644 (
    .a(_al_u643_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [41]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [9]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b9_var_o ));
  AL_MAP_LUT5 #(
    .EQN("~((E*~(C)*~(A)+E*C*~(A)+~(E)*C*A+E*C*A)*~(D)*~(B)+(E*~(C)*~(A)+E*C*~(A)+~(E)*C*A+E*C*A)*D*~(B)+~((E*~(C)*~(A)+E*C*~(A)+~(E)*C*A+E*C*A))*D*B+(E*~(C)*~(A)+E*C*~(A)+~(E)*C*A+E*C*A)*D*B)"),
    .INIT(32'h02ce13df))
    _al_u645 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [0]),
    .d(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .e(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(_al_u645_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*~(C)+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(C)+~(~A)*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C+~A*(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*C)"),
    .INIT(32'hf535c505))
    _al_u646 (
    .a(_al_u645_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [32]),
    .e(\u_PERIPH_TOP/timer_ribs_rdata [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_var_o ));
  AL_MAP_LUT5 #(
    .EQN("~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'h0c2e1d3f))
    _al_u647 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/tx_rdy ),
    .o(_al_u647_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(~A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'hf5c53505))
    _al_u648 (
    .a(_al_u647_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/rx_data [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b0_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    .INIT(16'h1d3f))
    _al_u649 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [3]),
    .o(_al_u649_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(~A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'hf5c53505))
    _al_u650 (
    .a(_al_u649_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [3]),
    .e(\u_PERIPH_TOP/u_USART2RIB/rx_data [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b3_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    .INIT(16'h1d3f))
    _al_u651 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [4]),
    .o(_al_u651_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(~A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'hf5c53505))
    _al_u652 (
    .a(_al_u651_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [4]),
    .e(\u_PERIPH_TOP/u_USART2RIB/rx_data [4]),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b4_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    .INIT(16'h1d3f))
    _al_u653 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [5]),
    .o(_al_u653_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(~A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'hf5c53505))
    _al_u654 (
    .a(_al_u653_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [5]),
    .e(\u_PERIPH_TOP/u_USART2RIB/rx_data [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b5_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    .INIT(16'h1d3f))
    _al_u655 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [7]),
    .o(_al_u655_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(~A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'hf5c53505))
    _al_u656 (
    .a(_al_u655_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [7]),
    .e(\u_PERIPH_TOP/u_USART2RIB/rx_data [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b7_var_o ));
  AL_MAP_LUT4 #(
    .EQN("~((D*A)*~(C)*~(B)+(D*A)*C*~(B)+~((D*A))*C*B+(D*A)*C*B)"),
    .INIT(16'h1d3f))
    _al_u657 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [6]),
    .o(_al_u657_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(~A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'hf5c53505))
    _al_u658 (
    .a(_al_u657_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [6]),
    .e(\u_PERIPH_TOP/u_USART2RIB/rx_data [6]),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b6_var_o ));
  AL_MAP_LUT5 #(
    .EQN("~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'h0c2e1d3f))
    _al_u659 (
    .a(periph_addr[2]),
    .b(periph_wrcs),
    .c(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/rx_vld ),
    .o(_al_u659_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(~A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'hf5c53505))
    _al_u660 (
    .a(_al_u659_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/rx_data [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b1_var_o ));
  AL_MAP_LUT5 #(
    .EQN("~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*~(D)*~(C)+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*D*~(C)+~((A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B))*D*C+(A*~(E)*~(B)+A*E*~(B)+~(A)*E*B+A*E*B)*D*C)"),
    .INIT(32'h01f10dfd))
    _al_u661 (
    .a(\u_PERIPH_TOP/u_USART2RIB/rx_err ),
    .b(periph_addr[2]),
    .c(periph_wrcs),
    .d(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [2]),
    .o(_al_u661_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(~A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+~A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'hf5c53505))
    _al_u662 (
    .a(_al_u661_o),
    .b(_al_u582_o),
    .c(periph_addr[3]),
    .d(\u_PERIPH_TOP/usart_rib_rdata [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/rx_data [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/sel0_b2_var_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u663 (
    .a(periph_addr[31]),
    .b(periph_addr[30]),
    .c(periph_addr[29]),
    .d(periph_addr[28]),
    .o(_al_u663_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u664 (
    .a(periph_addr[27]),
    .b(periph_addr[26]),
    .o(_al_u664_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u665 (
    .a(_al_u663_o),
    .b(_al_u664_o),
    .c(periph_addr[25]),
    .d(periph_addr[24]),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u666 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/timer_ribs_req ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u667 (
    .a(_al_u663_o),
    .b(_al_u664_o),
    .c(periph_addr[25]),
    .d(periph_addr[24]),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u668 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [0]),
    .o(\u_PERIPH_TOP/usart_rib_req ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u669 (
    .a(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [0]),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/n3 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u670 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/n3 ),
    .o(\u_PERIPH_TOP/u_SLAVE_SEL/n0 ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u671 (
    .a(periph_addr[7]),
    .b(periph_addr[6]),
    .c(periph_addr[5]),
    .d(periph_addr[4]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_8_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u672 (
    .a(periph_addr[15]),
    .b(periph_addr[14]),
    .c(periph_addr[13]),
    .d(periph_addr[12]),
    .o(_al_u672_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u673 (
    .a(_al_u672_o),
    .b(periph_addr[11]),
    .c(periph_addr[10]),
    .d(periph_addr[9]),
    .e(periph_addr[8]),
    .o(_al_u673_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u674 (
    .a(periph_addr[3]),
    .b(periph_addr[2]),
    .c(periph_wrcs),
    .o(_al_u674_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u675 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .c(_al_u673_o),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_8_sel_is_2_o ),
    .e(_al_u674_o),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/mux3_b0_sel_is_3_o ));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*A)"),
    .INIT(32'h00800000))
    _al_u676 (
    .a(_al_u673_o),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_8_sel_is_2_o ),
    .c(periph_addr[3]),
    .d(periph_addr[2]),
    .e(periph_wrcs),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u677 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[31]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [63]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [63]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u678 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [63]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [63]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [63]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((D*A))+B*C*~((D*A))+~(B)*C*(D*A)+B*C*(D*A))"),
    .INIT(16'he4cc))
    _al_u679 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n14 [63]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n12 [63]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [63]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u680 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[30]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [62]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [62]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u681 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [62]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [62]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [62]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u682 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [62]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [62]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [62]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u683 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[29]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [61]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [61]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u684 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [61]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [61]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [61]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u685 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [61]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [61]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [61]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u686 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[28]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [60]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [60]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u687 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [60]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [60]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [60]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u688 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [60]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [60]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [60]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u689 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[27]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [59]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [59]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u690 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [59]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [59]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [59]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u691 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [59]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [59]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [59]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u692 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[26]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [58]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [58]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u693 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [58]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [58]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [58]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u694 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [58]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [58]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [58]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u695 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[25]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [57]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [57]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u696 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [57]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [57]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [57]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u697 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [57]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [57]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [57]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u698 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[24]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [56]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [56]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u699 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [56]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [56]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [56]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u700 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [56]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [56]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [56]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u701 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[23]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [55]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [55]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u702 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [55]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [55]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [55]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u703 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [55]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [55]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [55]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u704 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[22]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [54]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [54]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u705 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [54]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [54]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [54]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u706 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [54]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [54]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [54]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u707 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[21]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [53]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [53]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u708 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [53]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [53]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [53]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u709 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [53]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [53]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [53]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u710 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[20]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [52]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [52]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u711 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [52]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [52]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [52]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u712 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [52]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [52]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [52]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u713 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[19]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [51]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [51]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u714 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [51]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [51]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [51]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u715 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [51]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [51]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [51]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u716 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[18]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [50]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [50]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u717 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [50]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [50]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [50]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u718 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [50]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [50]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [50]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u719 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[17]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [49]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [49]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u720 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [49]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [49]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [49]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u721 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [49]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [49]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [49]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u722 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[16]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [48]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [48]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u723 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [48]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [48]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [48]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u724 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [48]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [48]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [48]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u725 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[15]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [47]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [47]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u726 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [47]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [47]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [47]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u727 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [47]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [47]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [47]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u728 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[14]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [46]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [46]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u729 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [46]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [46]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [46]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u730 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [46]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [46]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [46]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u731 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[13]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [45]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [45]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u732 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [45]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [45]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [45]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u733 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [45]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [45]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [45]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u734 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[12]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [44]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [44]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u735 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [44]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [44]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [44]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u736 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [44]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [44]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [44]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u737 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[11]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [43]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [43]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u738 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [43]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [43]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [43]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u739 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [43]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [43]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [43]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u740 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[10]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [42]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [42]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u741 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [42]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [42]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [42]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u742 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [42]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [42]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [42]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u743 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[9]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [41]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [41]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u744 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [41]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [41]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [41]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u745 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [41]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [41]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [41]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u746 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[8]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [40]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [40]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u747 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [40]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [40]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [40]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u748 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [40]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [40]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [40]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u749 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[7]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [39]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [39]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u750 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [39]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [39]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [39]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u751 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [39]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [39]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [39]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u752 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[6]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [38]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [38]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u753 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [38]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [38]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [38]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u754 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [38]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [38]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [38]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u755 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[5]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [37]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [37]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u756 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [37]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [37]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [37]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u757 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [37]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [37]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [37]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u758 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[4]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [36]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [36]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u759 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [36]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [36]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [36]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u760 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [36]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [36]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [36]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u761 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[3]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [35]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [35]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u762 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [35]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [35]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [35]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u763 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [35]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [35]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [35]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u764 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[2]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [34]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [34]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u765 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [34]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [34]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [34]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u766 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [34]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [34]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [34]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u767 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[1]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [33]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [33]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u768 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [33]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [33]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [33]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u769 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [33]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [33]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [33]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u770 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/sel2_b32_sel_is_3_o ),
    .b(periph_wdata[0]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [32]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [32]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u771 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [32]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [32]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [32]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u772 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [32]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [32]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [32]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u773 (
    .a(periph_addr[3]),
    .b(periph_addr[2]),
    .c(periph_wrcs),
    .o(_al_u773_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u774 (
    .a(_al_u673_o),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_8_sel_is_2_o ),
    .c(_al_u773_o),
    .o(_al_u774_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*~B))"),
    .INIT(16'ha080))
    _al_u775 (
    .a(periph_req),
    .b(_al_u774_o),
    .c(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_en ),
    .o(\u_PERIPH_TOP/u_USART2RIB/n16 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u776 (
    .a(_al_u673_o),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_def_8_sel_is_2_o ),
    .c(reset),
    .o(_al_u776_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u777 (
    .a(periph_req),
    .b(_al_u776_o),
    .c(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u778 (
    .a(periph_req),
    .b(_al_u776_o),
    .c(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [0]),
    .d(_al_u773_o),
    .o(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u779 (
    .a(_al_u774_o),
    .b(periph_wdata[9]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [9]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u780 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [9]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [9]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [9]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u781 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [9]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [9]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [9]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u782 (
    .a(_al_u774_o),
    .b(periph_wdata[8]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [8]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u783 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [8]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [8]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [8]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u784 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [8]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [8]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u785 (
    .a(_al_u774_o),
    .b(periph_wdata[7]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [7]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u786 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [7]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [7]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [7]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u787 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [7]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [7]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u788 (
    .a(_al_u774_o),
    .b(periph_wdata[6]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [6]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u789 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [6]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [6]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [6]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u790 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [6]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [6]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u791 (
    .a(_al_u774_o),
    .b(periph_wdata[5]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [5]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u792 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [5]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [5]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [5]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u793 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [5]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [5]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u794 (
    .a(_al_u774_o),
    .b(periph_wdata[4]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [4]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u795 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [4]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [4]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [4]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u796 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [4]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [4]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u797 (
    .a(_al_u774_o),
    .b(periph_wdata[3]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [3]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u798 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [3]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [3]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [3]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u799 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [3]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [3]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u800 (
    .a(_al_u774_o),
    .b(periph_wdata[31]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [31]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u801 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [31]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [31]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [31]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u802 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [31]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [31]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u803 (
    .a(_al_u774_o),
    .b(periph_wdata[30]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [30]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u804 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [30]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [30]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [30]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u805 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [30]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [30]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [30]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u806 (
    .a(_al_u774_o),
    .b(periph_wdata[2]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [2]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u807 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [2]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [2]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [2]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'hdf80))
    _al_u808 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [2]),
    .c(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n14 [2]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u809 (
    .a(_al_u774_o),
    .b(periph_wdata[29]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [29]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u810 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [29]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [29]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [29]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u811 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [29]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [29]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [29]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u812 (
    .a(_al_u774_o),
    .b(periph_wdata[28]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [28]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u813 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [28]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [28]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [28]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u814 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [28]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [28]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [28]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u815 (
    .a(_al_u774_o),
    .b(periph_wdata[27]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [27]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u816 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [27]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [27]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [27]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u817 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [27]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [27]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [27]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u818 (
    .a(_al_u774_o),
    .b(periph_wdata[26]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [26]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u819 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [26]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [26]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [26]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u820 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [26]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [26]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [26]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u821 (
    .a(_al_u774_o),
    .b(periph_wdata[25]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [25]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u822 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [25]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [25]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [25]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u823 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [25]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [25]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [25]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u824 (
    .a(_al_u774_o),
    .b(periph_wdata[24]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [24]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u825 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [24]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [24]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [24]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u826 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [24]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [24]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [24]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u827 (
    .a(_al_u774_o),
    .b(periph_wdata[23]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [23]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u828 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [23]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [23]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [23]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u829 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [23]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [23]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [23]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u830 (
    .a(_al_u774_o),
    .b(periph_wdata[22]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [22]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u831 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [22]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [22]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [22]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u832 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [22]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [22]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [22]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u833 (
    .a(_al_u774_o),
    .b(periph_wdata[21]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [21]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u834 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [21]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [21]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [21]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u835 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [21]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [21]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [21]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u836 (
    .a(_al_u774_o),
    .b(periph_wdata[20]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [20]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u837 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [20]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [20]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [20]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u838 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [20]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [20]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [20]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u839 (
    .a(_al_u774_o),
    .b(periph_wdata[1]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [1]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u840 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [1]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [1]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [1]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'hdf80))
    _al_u841 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [1]),
    .c(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n14 [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u842 (
    .a(_al_u774_o),
    .b(periph_wdata[19]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [19]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u843 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [19]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [19]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [19]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u844 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [19]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [19]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [19]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u845 (
    .a(_al_u774_o),
    .b(periph_wdata[18]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [18]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u846 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [18]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [18]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [18]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u847 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [18]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [18]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [18]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u848 (
    .a(_al_u774_o),
    .b(periph_wdata[17]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [17]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u849 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [17]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [17]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [17]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u850 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [17]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [17]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [17]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u851 (
    .a(_al_u774_o),
    .b(periph_wdata[16]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [16]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u852 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [16]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [16]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [16]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u853 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [16]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [16]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [16]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u854 (
    .a(_al_u774_o),
    .b(periph_wdata[15]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [15]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u855 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [15]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [15]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [15]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u856 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [15]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [15]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u857 (
    .a(_al_u774_o),
    .b(periph_wdata[14]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [14]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u858 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [14]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [14]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [14]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u859 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [14]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [14]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u860 (
    .a(_al_u774_o),
    .b(periph_wdata[13]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [13]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u861 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [13]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [13]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [13]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u862 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [13]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [13]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u863 (
    .a(_al_u774_o),
    .b(periph_wdata[12]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [12]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u864 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [12]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [12]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [12]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u865 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [12]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [12]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u866 (
    .a(_al_u774_o),
    .b(periph_wdata[11]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [11]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u867 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [11]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [11]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [11]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u868 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [11]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [11]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u869 (
    .a(_al_u774_o),
    .b(periph_wdata[10]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [10]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u870 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [10]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [10]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [10]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B)*~((D*A))+C*B*~((D*A))+~(C)*B*(D*A)+C*B*(D*A))"),
    .INIT(16'hd8f0))
    _al_u871 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [10]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/n14 [10]),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u872 (
    .a(_al_u774_o),
    .b(periph_wdata[0]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n12 [0]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u873 (
    .a(\u_PERIPH_TOP/u_TIMER2RIB/n13 [0]),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [0]),
    .c(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n14 [0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'hdf80))
    _al_u874 (
    .a(periph_req),
    .b(\u_PERIPH_TOP/u_TIMER2RIB/n12 [0]),
    .c(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n14 [0]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/n18 [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u875 (
    .a(periph_req),
    .b(_al_u776_o),
    .c(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .o(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ));
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'h1))
    _al_u876 (
    .a(i_rstn_pad),
    .o(n0));
  AL_BUFKEEP #(
    .KEEP("OUT"))
    _bufkeep_clk_84mhz (
    .i(clk_84mhz_keep),
    .o(clk_84mhz));  // ../RTL/soc_top/soc_top.v(16)
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  CORE_TOP u_CORE_TOP (
    .i_clk(clk_84mhz),
    .i_ribp_gnt(\u_PERIPH_TOP/u_SLAVE_SEL/n0 ),
    .i_ribp_rdata(periph_rdata),
    .i_ribp_rsp(\u_PERIPH_TOP/u_SLAVE_SEL/n1 ),
    .i_ribx_gnt(1'b0),
    .i_ribx_rdata(32'b00000000000000000000000000000000),
    .i_ribx_rsp(1'b0),
    .i_rstn(reset),
    .o_ribp_addr({periph_addr[31:24],open_n115,open_n116,open_n117,open_n118,open_n119,open_n120,open_n121,open_n122,periph_addr[15:2],open_n123,open_n124}),
    .o_ribp_req(periph_req),
    .o_ribp_wdata(periph_wdata),
    .o_ribp_wrcs(periph_wrcs));  // ../RTL/soc_top/soc_top.v(51)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("SET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_SLAVE_SEL/default_cs_reg  (
    .ce(\u_PERIPH_TOP/u_SLAVE_SEL/n6 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/n3 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_SLAVE_SEL/default_cs ));  // ../RTL/core/rib.v(121)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_SLAVE_SEL/handshake_rdy_last_reg  (
    .ce(\u_PERIPH_TOP/u_SLAVE_SEL/n6 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/n0 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_SLAVE_SEL/handshake_rdy_last ));  // ../RTL/core/rib.v(121)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_SLAVE_SEL/reg0_b0  (
    .ce(\u_PERIPH_TOP/u_SLAVE_SEL/n6 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_SLAVE_SEL/sel_tag_id [0]));  // ../RTL/core/rib.v(121)
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u11_al_u880  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [13],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [11]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [14],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [12]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c11 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [13],\u_PERIPH_TOP/u_TIMER2RIB/n13 [11]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c15 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [14],\u_PERIPH_TOP/u_TIMER2RIB/n13 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u15_al_u881  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [17],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [15]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [18],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [16]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c15 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [17],\u_PERIPH_TOP/u_TIMER2RIB/n13 [15]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c19 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [18],\u_PERIPH_TOP/u_TIMER2RIB/n13 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u19_al_u882  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [21],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [19]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [22],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [20]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c19 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [21],\u_PERIPH_TOP/u_TIMER2RIB/n13 [19]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c23 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [22],\u_PERIPH_TOP/u_TIMER2RIB/n13 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u23_al_u883  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [25],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [23]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [26],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [24]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c23 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [25],\u_PERIPH_TOP/u_TIMER2RIB/n13 [23]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c27 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [26],\u_PERIPH_TOP/u_TIMER2RIB/n13 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u27_al_u884  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [29],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [27]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [30],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [28]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c27 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [29],\u_PERIPH_TOP/u_TIMER2RIB/n13 [27]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c31 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [30],\u_PERIPH_TOP/u_TIMER2RIB/n13 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u31_al_u885  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [33],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [31]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [34],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [32]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c31 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [33],\u_PERIPH_TOP/u_TIMER2RIB/n13 [31]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c35 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [34],\u_PERIPH_TOP/u_TIMER2RIB/n13 [32]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u35_al_u886  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [37],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [35]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [38],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [36]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c35 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [37],\u_PERIPH_TOP/u_TIMER2RIB/n13 [35]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c39 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [38],\u_PERIPH_TOP/u_TIMER2RIB/n13 [36]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u39_al_u887  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [41],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [39]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [42],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [40]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c39 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [41],\u_PERIPH_TOP/u_TIMER2RIB/n13 [39]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c43 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [42],\u_PERIPH_TOP/u_TIMER2RIB/n13 [40]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u3_al_u878  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [5],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [3]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [6],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [4]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c3 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [5],\u_PERIPH_TOP/u_TIMER2RIB/n13 [3]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c7 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [6],\u_PERIPH_TOP/u_TIMER2RIB/n13 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u43_al_u888  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [45],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [43]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [46],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [44]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c43 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [45],\u_PERIPH_TOP/u_TIMER2RIB/n13 [43]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c47 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [46],\u_PERIPH_TOP/u_TIMER2RIB/n13 [44]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y6Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u47_al_u889  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [49],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [47]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [50],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [48]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c47 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [49],\u_PERIPH_TOP/u_TIMER2RIB/n13 [47]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c51 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [50],\u_PERIPH_TOP/u_TIMER2RIB/n13 [48]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y6Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u51_al_u890  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [53],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [51]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [54],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [52]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c51 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [53],\u_PERIPH_TOP/u_TIMER2RIB/n13 [51]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c55 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [54],\u_PERIPH_TOP/u_TIMER2RIB/n13 [52]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y7Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u55_al_u891  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [57],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [55]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [58],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [56]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c55 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [57],\u_PERIPH_TOP/u_TIMER2RIB/n13 [55]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c59 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [58],\u_PERIPH_TOP/u_TIMER2RIB/n13 [56]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y7Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u59_al_u892  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [61],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [59]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [62],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [60]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c59 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [61],\u_PERIPH_TOP/u_TIMER2RIB/n13 [59]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c63 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [62],\u_PERIPH_TOP/u_TIMER2RIB/n13 [60]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y8Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u63_al_u893  (
    .a({open_n453,\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [63]}),
    .c(2'b00),
    .d({open_n458,1'b0}),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c63 ),
    .f({open_n475,\u_PERIPH_TOP/u_TIMER2RIB/n13 [63]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/u7_al_u879  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [9],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [7]}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [10],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [8]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_PERIPH_TOP/u_TIMER2RIB/add0/c7 ),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [9],\u_PERIPH_TOP/u_TIMER2RIB/n13 [7]}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c11 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [10],\u_PERIPH_TOP/u_TIMER2RIB/n13 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_TIMER2RIB/add0/ucin_al_u877  (
    .a({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [1],1'b0}),
    .b({\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [2],\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [0]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({\u_PERIPH_TOP/u_TIMER2RIB/n13 [1],open_n516}),
    .fco(\u_PERIPH_TOP/u_TIMER2RIB/add0/c3 ),
    .fx({\u_PERIPH_TOP/u_TIMER2RIB/n13 [2],\u_PERIPH_TOP/u_TIMER2RIB/n13 [0]}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/o_ribs_rsp_reg  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/timer_ribs_req ),
    .sr(reset),
    .q(\u_PERIPH_TOP/timer_ribs_rsp ));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [0]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b1  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [1]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b10  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [10]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [10]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b11  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [11]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [11]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b12  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [12]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [12]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b13  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [13]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [13]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b14  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [14]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [14]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b15  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [15]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [15]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b16  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [16]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [16]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b17  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [17]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [17]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b18  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [18]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [18]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b19  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [19]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [19]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b2  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [2]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b20  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [20]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [20]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b21  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [21]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [21]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b22  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [22]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [22]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b23  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [23]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [23]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b24  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [24]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [24]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b25  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [25]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [25]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b26  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [26]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [26]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b27  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [27]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [27]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b28  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [28]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [28]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b29  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [29]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [29]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b3  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [3]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [3]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b30  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [30]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [30]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b31  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [31]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [31]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b32  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [32]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [32]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b33  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [33]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [33]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b34  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [34]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [34]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b35  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [35]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [35]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b36  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [36]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [36]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b37  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [37]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [37]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b38  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [38]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [38]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b39  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [39]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [39]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b4  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [4]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [4]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b40  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [40]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [40]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b41  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [41]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [41]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b42  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [42]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [42]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b43  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [43]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [43]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b44  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [44]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [44]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b45  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [45]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [45]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b46  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [46]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [46]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b47  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [47]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [47]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b48  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [48]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [48]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b49  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [49]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [49]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b5  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [5]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [5]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b50  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [50]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [50]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b51  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [51]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [51]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b52  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [52]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [52]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b53  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [53]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [53]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b54  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [54]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [54]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b55  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [55]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [55]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b56  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [56]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [56]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b57  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [57]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [57]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b58  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [58]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [58]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b59  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [59]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [59]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b6  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [6]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [6]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b60  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [60]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [60]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b61  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [61]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [61]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b62  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [62]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [62]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b63  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [63]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [63]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b7  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [7]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [7]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b8  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [8]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [8]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg0_b9  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/n18 [9]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_cnt [9]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b0  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b0_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [0]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b1  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b1_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [1]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b10  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b10_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [10]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b11  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b11_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [11]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b12  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b12_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [12]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b13  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b13_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [13]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b14  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b14_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [14]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b15  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b15_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [15]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b16  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b16_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [16]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b17  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b17_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [17]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b18  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b18_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [18]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b19  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b19_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [19]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b2  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b2_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [2]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b20  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b20_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [20]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b21  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b21_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [21]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b22  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b22_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [22]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b23  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b23_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [23]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b24  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b24_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [24]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b25  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b25_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [25]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b26  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b26_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [26]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b27  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b27_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [27]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b28  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b28_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [28]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b29  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b29_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [29]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b3  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b3_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [3]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b30  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b30_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [30]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b31  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b31_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [31]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b4  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b4_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [4]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b5  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b5_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [5]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b6  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b6_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [6]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b7  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b7_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [7]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b8  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b8_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [8]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg1_b9  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux7_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_TIMER2RIB/sel1_b9_var_o ),
    .q(\u_PERIPH_TOP/timer_ribs_rdata [9]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("SET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_TIMER2RIB/reg2_b0  (
    .ce(\u_PERIPH_TOP/u_TIMER2RIB/mux3_b0_sel_is_3_o ),
    .clk(clk_84mhz),
    .d(periph_wdata[0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_TIMER2RIB/timer_ctrl [0]));  // ../RTL/periph/timer2rib.v(34)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/o_ribs_rsp_reg  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/usart_rib_req ),
    .sr(reset),
    .q(\u_PERIPH_TOP/usart_rib_rsp ));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg0_b0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b0_var_o ),
    .q(\u_PERIPH_TOP/usart_rib_rdata [0]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg0_b1  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b1_var_o ),
    .q(\u_PERIPH_TOP/usart_rib_rdata [1]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg0_b2  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b2_var_o ),
    .q(\u_PERIPH_TOP/usart_rib_rdata [2]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg0_b3  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b3_var_o ),
    .q(\u_PERIPH_TOP/usart_rib_rdata [3]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg0_b4  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b4_var_o ),
    .q(\u_PERIPH_TOP/usart_rib_rdata [4]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg0_b5  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b5_var_o ),
    .q(\u_PERIPH_TOP/usart_rib_rdata [5]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg0_b6  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b6_var_o ),
    .q(\u_PERIPH_TOP/usart_rib_rdata [6]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg0_b7  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux3_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/sel0_b7_var_o ),
    .q(\u_PERIPH_TOP/usart_rib_rdata [7]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg1_b0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(periph_wdata[0]),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [0]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg1_b1  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(periph_wdata[1]),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [1]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg1_b2  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(periph_wdata[2]),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [2]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg1_b3  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(periph_wdata[3]),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [3]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg1_b4  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(periph_wdata[4]),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [4]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg1_b5  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(periph_wdata[5]),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [5]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg1_b6  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(periph_wdata[6]),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [6]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_PERIPH_TOP/u_USART2RIB/reg1_b7  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/mux5_b0_sel_is_2_o ),
    .clk(clk_84mhz),
    .d(periph_wdata[7]),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [7]));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/tx_en_reg  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/n16 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_en ));  // ../RTL/periph/usart2rib.v(48)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A78C4C0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB840 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCD90 ));  // al_ip/usart_gate.v(1818)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A78F160  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A832EE0 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ));  // al_ip/usart_gate.v(1468)
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F940|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F610"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"),
    .REG1_REGSET("RESET"),
    .REG1_SD("F"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A78F490|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A880B50  (
    .a(2'b01),
    .b({1'b1,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [5]}),
    .clk(clk_84mhz),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830390 ),
    .sr(reset),
    .f({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ,open_n652}),
    .q({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ,open_n656}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A826290  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [3]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [3]));  // al_ip/usart_gate.v(1594)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8268F0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [2]));  // al_ip/usart_gate.v(1558)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A826F50  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [1]));  // al_ip/usart_gate.v(1549)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A827060  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [5]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [5]));  // al_ip/usart_gate.v(1612)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("SET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A827390  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D50E0 ),
    .sr(reset),
    .q(o_io_tx_pad));  // al_ip/usart_gate.v(2358)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A827D20  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [4]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [4]));  // al_ip/usart_gate.v(1603)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A827F40  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [1]));  // al_ip/usart_gate.v(1576)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A828380  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 [0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [0]));  // al_ip/usart_gate.v(1540)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8285A0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5BE0 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4480 ));  // al_ip/usart_gate.v(2367)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8298C0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [0]));  // al_ip/usart_gate.v(1567)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A829F20  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD890 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2010 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5A80 ));  // al_ip/usart_gate.v(2376)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82A360  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [2]));  // al_ip/usart_gate.v(1585)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("SET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82CBC0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4320 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/tx_rdy ));  // al_ip/usart_gate.v(2385)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82CCD0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D3FB0 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5B30 ));  // al_ip/usart_gate.v(2394)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A876BF0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [3]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [3]));  // al_ip/usart_gate.v(1854)
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'b0000010010001100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A877360  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0A20 ));  // al_ip/usart_gate.v(785)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A877470  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [2]));  // al_ip/usart_gate.v(1881)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A877580  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [5]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [5]));  // al_ip/usart_gate.v(1971)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~(~C*~B)))"),
    .INIT(32'b10101010101010101010101000000010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8779C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1100 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA22E0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1940 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [3]));  // al_ip/usart_gate.v(765)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A877AD0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [3]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [3]));  // al_ip/usart_gate.v(1953)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A877F10  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]));  // al_ip/usart_gate.v(1908)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878130  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [1]));  // al_ip/usart_gate.v(1935)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878240  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [3]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [3]));  // al_ip/usart_gate.v(1890)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878350  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [6]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [6]));  // al_ip/usart_gate.v(1980)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878460  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [0]));  // al_ip/usart_gate.v(1998)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878570  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [0]));  // al_ip/usart_gate.v(1827)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878680  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]));  // al_ip/usart_gate.v(1917)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878790  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [1]));  // al_ip/usart_gate.v(2007)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878AC0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [1]));  // al_ip/usart_gate.v(1836)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878BD0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 [0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]));  // al_ip/usart_gate.v(1899)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111000010111111011100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878CE0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1F70 ));  // al_ip/usart_gate.v(775)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878DF0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [7]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [7]));  // al_ip/usart_gate.v(1989)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A878F00  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [3]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [2]));  // al_ip/usart_gate.v(2016)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879120  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [1]));  // al_ip/usart_gate.v(1872)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'b0000001000000111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879450  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [2]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0760 ));  // al_ip/usart_gate.v(794)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~(~C*~B)))"),
    .INIT(32'b10101010101010101010101000000010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879560  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1F70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0A20 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0760 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [2]));  // al_ip/usart_gate.v(803)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879670  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0]));  // al_ip/usart_gate.v(1926)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879890  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2]));  // al_ip/usart_gate.v(1944)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879BC0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [0]));  // al_ip/usart_gate.v(1863)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879CD0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [4]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [4]));  // al_ip/usart_gate.v(1962)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879DE0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [4]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [3]));  // al_ip/usart_gate.v(2025)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A879EF0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [5]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [4]));  // al_ip/usart_gate.v(2034)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'b0000001000000111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87A000  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [3]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1940 ));  // al_ip/usart_gate.v(756)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87A110  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [2]));  // al_ip/usart_gate.v(1845)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87A220  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [6]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [5]));  // al_ip/usart_gate.v(2043)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87A440  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCA20 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [7]));  // al_ip/usart_gate.v(2061)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87A550  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_data [7]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_data [6]));  // al_ip/usart_gate.v(2052)
  AL_MAP_LUT1 #(
    .EQN("(~A)"),
    .INIT(2'b01))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87B650  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 [0]));  // al_ip/usart_gate.v(813)
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87D850|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87FD80"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87D850|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87FD80  (
    .a({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [0],1'b0}),
    .b(2'b10),
    .f({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [0],open_n698}),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82ECE0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87D850|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87FD80"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87EC80_al_u894  (
    .a({open_n703,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [5]}),
    .b({open_n704,1'b0}),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FB50 ),
    .f({open_n723,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [5]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87D850|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87FD80"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87EEA0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87D960  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [2:1]),
    .b(2'b00),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82ECE0 ),
    .f(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [2:1]),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E4A0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87D850|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87FD80"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F720|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A881C50  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [4:3]),
    .b(2'b00),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E4A0 ),
    .f(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [4:3]),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FB50 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F940|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F610"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F940|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F610  (
    .a(2'b01),
    .b({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [0],1'b0}),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E600 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F940|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F610"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8800B0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87FFA0  (
    .a(2'b10),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [2:1]),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82E600 ),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FCB0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F940|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A87F610"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8801C0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A880930  (
    .a(2'b01),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54D8D0 [4:3]),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A82FCB0 ),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830390 ));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A881A30  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4C10 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D3FB0 ));  // al_ip/usart_gate.v(2403)
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A932BF0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935230"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9326A0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936770  (
    .a(2'b11),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2:1]),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535380 ),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533EE0 ));
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("SET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9327B0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A832AC0 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [3]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCA20 ));  // al_ip/usart_gate.v(2088)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9328C0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [7]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [7]));  // al_ip/usart_gate.v(2349)
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A932BF0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935230"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A932BF0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935230  (
    .a(2'b11),
    .b({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0],1'b0}),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535380 ));
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A932D00  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [0]));  // al_ip/usart_gate.v(2124)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933140  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [3]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [3]));  // al_ip/usart_gate.v(2313)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933250  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]));  // al_ip/usart_gate.v(2295)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933360  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [0]));  // al_ip/usart_gate.v(2286)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("LATCH"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933580  (
    .clk(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2F30 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 [0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [0]));  // al_ip/usart_gate.v(2223)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9337A0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [1]));  // al_ip/usart_gate.v(2133)
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9338B0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934F00"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9338B0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934F00  (
    .a({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0],1'b0}),
    .b(2'b10),
    .f({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [0],open_n920}),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5335F0 ));
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9339C0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [2]));  // al_ip/usart_gate.v(2142)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933BE0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [5]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [5]));  // al_ip/usart_gate.v(2169)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933CF0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]));  // al_ip/usart_gate.v(2205)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("LATCH"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933E00  (
    .clk(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2F30 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [2]));  // al_ip/usart_gate.v(2241)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933F10  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]));  // al_ip/usart_gate.v(2250)
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9338B0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934F00"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934130|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936110  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [4:3]),
    .b(2'b00),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533120 ),
    .f(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [4:3]),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534880 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9338B0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934F00"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934240_al_u895  (
    .a({open_n950,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [7]}),
    .b({open_n951,1'b0}),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534510 ),
    .f({open_n970,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [7]}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934350  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB2C0 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/rx_vld ));  // al_ip/usart_gate.v(2079)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934460  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [2]));  // al_ip/usart_gate.v(2304)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934570  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB790 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CBF20 ));  // al_ip/usart_gate.v(2097)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934680  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]));  // al_ip/usart_gate.v(2259)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9348A0  (
    .clk(clk_84mhz),
    .d(i_io_rx_pad),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB790 ));  // al_ip/usart_gate.v(2106)
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9338B0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934F00"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934CE0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A933AD0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2:1]),
    .b(2'b00),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A5335F0 ),
    .f(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [2:1]),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533120 ));
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934DF0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [4]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [4]));  // al_ip/usart_gate.v(2160)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935010  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]));  // al_ip/usart_gate.v(2214)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935120  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [4]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [4]));  // al_ip/usart_gate.v(2322)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935340  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [2]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]));  // al_ip/usart_gate.v(2268)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935560  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [6]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [6]));  // al_ip/usart_gate.v(2340)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935670  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [0]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]));  // al_ip/usart_gate.v(2196)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935780  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [3]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [3]));  // al_ip/usart_gate.v(2277)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935890  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [7]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [7]));  // al_ip/usart_gate.v(2187)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935AB0  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB420 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CC810 ));  // al_ip/usart_gate.v(2115)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935CD0  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [3]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [3]));  // al_ip/usart_gate.v(2151)
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A9338B0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A934F00"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935DE0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936660  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [6:5]),
    .b(2'b00),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534880 ),
    .f(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [6:5]),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534510 ));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936000  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [5]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [5]));  // al_ip/usart_gate.v(2331)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936220  (
    .ce(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/tx_buffer [6]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [6]));  // al_ip/usart_gate.v(2178)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("INV"),
    .DFFMODE("LATCH"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936330  (
    .clk(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2F30 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 [1]),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [1]));  // al_ip/usart_gate.v(2232)
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A932BF0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935230"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A937760|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A936BB0  (
    .a(2'b00),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [6:5]),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535430 ),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535590 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A932BF0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935230"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A938640|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A937BA0  (
    .a(2'b00),
    .b({1'b1,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [7]}),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535590 ),
    .f({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ,open_n1076}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A938970  (
    .clk(clk_84mhz),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB6E0 ),
    .sr(reset),
    .q(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD470 ));  // al_ip/usart_gate.v(2070)
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A932BF0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A935230"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A938EC0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A939EB0  (
    .a(2'b01),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [4:3]),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A533EE0 ),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535430 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C710|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A937CB0"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93AD90|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C820  (
    .a(2'b11),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [6:5]),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535640 ),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534250 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C710|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A937CB0"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C0B0|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93DE70  (
    .a(2'b00),
    .b({1'b1,\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [7]}),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534250 ),
    .f({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C93D0 ,open_n1149}));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C710|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A937CB0"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C600|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93B2E0  (
    .a(2'b11),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [4:3]),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534BF0 ),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A535640 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C710|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A937CB0"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C710|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A937CB0  (
    .a(2'b11),
    .b({\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0],1'b0}),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534B40 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C710|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A937CB0"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93D700|u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A93C2D0  (
    .a(2'b11),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2:1]),
    .fci(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534B40 ),
    .fco(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A534BF0 ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(D@C)))"),
    .INIT(16'b1000110011001000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA080  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C9110 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [0]));  // al_ip/usart_gate.v(1186)
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'b00101000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA190  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FFD0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CBF20 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [0]));  // al_ip/usart_gate.v(1236)
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*~B))*~(C)+~A*(D*~B)*~(C)+~(~A)*(D*~B)*C+~A*(D*~B)*C)"),
    .INIT(16'b0011010100000101))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA2A0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0290 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [2]));  // al_ip/usart_gate.v(1270)
  AL_MAP_LUT5 #(
    .EQN("(~B*(~E*~((~D*~A))*~(C)+~E*(~D*~A)*~(C)+~(~E)*(~D*~A)*C+~E*(~D*~A)*C))"),
    .INIT(32'b00000000000100000000001100010011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA3B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FF20 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [0]),
    .e(o_io_tx_pad),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E710 ));  // al_ip/usart_gate.v(1397)
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*B*A))"),
    .INIT(16'b0000000001111111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA4C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F160 ));  // al_ip/usart_gate.v(1109)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*B*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11001000110011111111011111111111),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA5D0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A340 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F580 ));  // al_ip/usart_gate.v(1286)
  AL_MAP_LUT5 #(
    .EQN("(A*~((E*~(B)*~(C)+E*B*~(C)+~(E)*B*C+E*B*C))*~(D)+A*(E*~(B)*~(C)+E*B*~(C)+~(E)*B*C+E*B*C)*~(D)+~(A)*(E*~(B)*~(C)+E*B*~(C)+~(E)*B*C+E*B*C)*D+A*(E*~(B)*~(C)+E*B*~(C)+~(E)*B*C+E*B*C)*D)"),
    .INIT(32'b11001111101010101100000010101010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA6E0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5D780 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A68B0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [0]));  // al_ip/usart_gate.v(266)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA7F0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F370 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F8F0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [6]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [6]));  // al_ip/usart_gate.v(336)
  AL_MAP_LUT5 #(
    .EQN("(A*~((~C*~B))*D*~(E)+A*(~C*~B)*D*~(E)+~(A)*(~C*~B)*~(D)*E+A*(~C*~B)*~(D)*E)"),
    .INIT(32'b00000000000000111010101000000000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACA900  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0080 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 [2]));  // al_ip/usart_gate.v(1332)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACAA10  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F4D0 ));  // al_ip/usart_gate.v(355)
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~(C*~B)*~(A)*~(D)+~(C*~B)*A*~(D)+~(~(C*~B))*A*D+~(C*~B)*A*D))"),
    .INIT(32'b00000000000000000101010100110000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACAB20  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0080 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A68B0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F210 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 [1]));  // al_ip/usart_gate.v(246)
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(C*A)))"),
    .INIT(16'b1110110000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACAC30  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DCC0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .d(reset),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 [0]));  // al_ip/usart_gate.v(1369)
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*~B))*~(C)+~A*(D*~B)*~(C)+~(~A)*(D*~B)*C+~A*(D*~B)*C)"),
    .INIT(16'b0011010100000101))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACAD40  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F420 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [1]));  // al_ip/usart_gate.v(1090)
  AL_MAP_LUT5 #(
    .EQN("(E*A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(32'b10001000101000000000000000000000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACAE50  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C93D0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5BBF0 ));  // al_ip/usart_gate.v(1099)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACAF60  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5A80 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9D8A0 ));  // al_ip/usart_gate.v(1407)
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'b0001))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB070  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ),
    .b(o_io_tx_pad),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DE20 ));  // al_ip/usart_gate.v(229)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB180  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CBF20 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C9110 ));  // al_ip/usart_gate.v(1127)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'b1000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB290  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A550 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A340 ));  // al_ip/usart_gate.v(1279)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB3A0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [6]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [6]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F370 ));  // al_ip/usart_gate.v(320)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB4B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [5]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FA50 ));  // al_ip/usart_gate.v(346)
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(C*A)))"),
    .INIT(16'b1100110010000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB5C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DC10 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [3]));  // al_ip/usart_gate.v(1149)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB6D0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [6]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F8F0 ));  // al_ip/usart_gate.v(329)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB7E0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [7]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DED0 ));  // al_ip/usart_gate.v(286)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'b10101011100010111101111111111111),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACB8F0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F420 ));  // al_ip/usart_gate.v(1072)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACBA00  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [4]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [4]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F630 ));  // al_ip/usart_gate.v(372)
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*(D@A))"),
    .INIT(16'b0101000110100010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACBB10  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA01E0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD470 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB6E0 ));  // al_ip/usart_gate.v(1388)
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'b0001000001010000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACBC20  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DA00 ));  // al_ip/usart_gate.v(1342)
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'b00000010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACBD30  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ));  // al_ip/usart_gate.v(1082)
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'b10000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACBE40  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CBF20 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830C80 ));  // al_ip/usart_gate.v(1202)
  AL_MAP_LUT4 #(
    .EQN("(A*(C@(D*B)))"),
    .INIT(16'b0010100010100000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACBF50  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FFD0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CBF20 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [1]));  // al_ip/usart_gate.v(1227)
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*A)))"),
    .INIT(16'b1100100011000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC060  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FF20 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0080 ));  // al_ip/usart_gate.v(1313)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~(E*~C)*~(B)*~(D)+~(E*~C)*B*~(D)+~(~(E*~C))*B*D+~(E*~C)*B*D))"),
    .INIT(32'b00100010000010100010001000000000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC170  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C93D0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ));  // al_ip/usart_gate.v(276)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC280  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9D950 ));  // al_ip/usart_gate.v(303)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC390  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FA50 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F4D0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [5]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [5]));  // al_ip/usart_gate.v(362)
  AL_MAP_LUT4 #(
    .EQN("(A*(D@(C*B)))"),
    .INIT(16'b0010101010000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC4A0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FFD0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830C80 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [3]));  // al_ip/usart_gate.v(1210)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'b10111010000000001011101010111011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC5B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E710 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9D8A0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .e(o_io_tx_pad),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EDF0 ));  // al_ip/usart_gate.v(1414)
  AL_MAP_LUT5 #(
    .EQN("(A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'b10111011101100001000110010000000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC6C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A68B0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5D780 ));  // al_ip/usart_gate.v(256)
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'b10000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC7D0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C9110 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DC10 ));  // al_ip/usart_gate.v(1134)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC8E0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F630 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0340 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [4]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [4]));  // al_ip/usart_gate.v(388)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACC9F0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F9A0 ));  // al_ip/usart_gate.v(407)
  AL_MAP_LUT4 #(
    .EQN("(B*(A*~(C)*~(D)+~(A)*C*~(D)+A*~(C)*D+~(A)*C*D+A*C*D))"),
    .INIT(16'b1100100001001000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACCB00  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DC10 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [2]));  // al_ip/usart_gate.v(1158)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACCC10  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [4]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0340 ));  // al_ip/usart_gate.v(381)
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*~B))*~(C)+~A*(D*~B)*~(C)+~(~A)*(D*~B)*C+~A*(D*~B)*C)"),
    .INIT(16'b0011010100000101))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACCD20  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F580 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8670 [3]));  // al_ip/usart_gate.v(1296)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACCE30  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [3]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E240 ));  // al_ip/usart_gate.v(398)
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'b00101000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACCF40  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FFD0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830C80 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55B0F0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A772F10 [2]));  // al_ip/usart_gate.v(1219)
  AL_MAP_LUT5 #(
    .EQN("(B*~(~A*~(E@(D*C))))"),
    .INIT(32'b10001100110011001100100010001000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD050  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C9110 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A76D950 [1]));  // al_ip/usart_gate.v(1176)
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'b0000000010000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD160  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C95E0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DAB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A833D50 ));  // al_ip/usart_gate.v(1244)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD270  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E240 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F9A0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [3]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [3]));  // al_ip/usart_gate.v(414)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD380  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F000 ));  // al_ip/usart_gate.v(424)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'b1000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD490  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A550 ));  // al_ip/usart_gate.v(1253)
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*A)"),
    .INIT(32'b00000000100000000000000000000000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD5A0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C95E0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DAB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCA20 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA01E0 ));  // al_ip/usart_gate.v(1378)
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'b0001))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD6B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C95E0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FFD0 ));  // al_ip/usart_gate.v(1195)
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'b00000100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD7C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ));  // al_ip/usart_gate.v(295)
  AL_MAP_LUT5 #(
    .EQN("(~B*~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*~(C)+~B*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)+~(~B)*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C+~B*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C)"),
    .INIT(32'b11110011010100111010001100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD8D0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [0]),
    .e(o_io_tx_pad),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5F070 ));  // al_ip/usart_gate.v(219)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACD9E0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DED0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9D950 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [7]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [7]));  // al_ip/usart_gate.v(310)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'b1000000000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACDAF0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897F10 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ));  // al_ip/usart_gate.v(1167)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~C*~B))"),
    .INIT(32'b10101010101010101010101010101000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACDC00  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ));  // al_ip/usart_gate.v(1322)
  AL_MAP_LUT5 #(
    .EQN("~((~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*~(C)*~(E)+(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*C*~(E)+~((~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))*C*E+(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)*C*E)"),
    .INIT(32'b00001111000011110101010111001100),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACDD10  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EDF0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5F070 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DE20 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D50E0 ));  // al_ip/usart_gate.v(236)
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*~A)"),
    .INIT(16'b0000000000010000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACDE20  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5BBF0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F160 ),
    .c(reset),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 [1]));  // al_ip/usart_gate.v(1118)
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'b0001))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACDF30  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ));  // al_ip/usart_gate.v(1142)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*B*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11001000110011111111011111111111),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE040  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A53A550 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA0290 ));  // al_ip/usart_gate.v(1260)
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'b10000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE150  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FF20 ));  // al_ip/usart_gate.v(1305)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~A*~(D*B)))"),
    .INIT(16'b0000111000001010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE260  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DA00 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F840 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4480 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A5F10 [0]));  // al_ip/usart_gate.v(1351)
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(B*A))"),
    .INIT(16'b0000000001110000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE370  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DCC0 ));  // al_ip/usart_gate.v(1360)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE480  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DF80 ));  // al_ip/usart_gate.v(459)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE590  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E920 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F6E0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [0]));  // al_ip/usart_gate.v(492)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACE7B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FB00 ));  // al_ip/usart_gate.v(433)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'b0000010000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACED00  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FF20 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ));  // al_ip/usart_gate.v(520)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACF580  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F000 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FB00 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [2]));  // al_ip/usart_gate.v(440)
  AL_MAP_LUT5 #(
    .EQN("(D*(B*~((C*~A))*~(E)+B*(C*~A)*~(E)+~(B)*(C*~A)*E+B*(C*~A)*E))"),
    .INIT(32'b01010000000000001100110000000000),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACF690  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FC60 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA5BBF0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E3A0 ),
    .d(reset),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8988B0 [2]));  // al_ip/usart_gate.v(510)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AACF7A0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [1]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A7020 [1]));  // al_ip/usart_gate.v(537)
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'b0100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD0020  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F6E0 ));  // al_ip/usart_gate.v(485)
  AL_MAP_LUT5 #(
    .EQN("~(A*~((~C*~(D*B)))*~(E)+A*(~C*~(D*B))*~(E)+~(A)*(~C*~(D*B))*E+A*(~C*~(D*B))*E)"),
    .INIT(32'b11111100111100000101010101010101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD0680  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E7C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E870 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DF80 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A899100 [1]));  // al_ip/usart_gate.v(466)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD0DF0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E920 ));  // al_ip/usart_gate.v(476)
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'b11001000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD1340  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E5B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FC60 ));  // al_ip/usart_gate.v(502)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD1670  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA63600 ));  // al_ip/usart_gate.v(529)
  AL_MAP_LUT5 #(
    .EQN("(A*~((D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B))*~(C)+A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*~(C)+~(A)*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C+A*(D*~(E)*~(B)+D*E*~(B)+~(D)*E*B+D*E*B)*C)"),
    .INIT(32'b11111010110010100011101000001010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD1780  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A7020 [1]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA60730 ));  // al_ip/usart_gate.v(545)
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'b0100110001011111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD2220  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F2C0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A897880 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E7C0 ));  // al_ip/usart_gate.v(450)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'b10101010000011001111111100111111),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD2BB0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [7]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FDC0 ));  // al_ip/usart_gate.v(603)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111000010111111011100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD2DD0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [0]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E0E0 ));  // al_ip/usart_gate.v(565)
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'b0000010010001100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD3100  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [6]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EA80 ));  // al_ip/usart_gate.v(633)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'b0000001000000111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD3320  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [5]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EC90 ));  // al_ip/usart_gate.v(680)
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'b0000010010001100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD3A90  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [5]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [6]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EBE0 ));  // al_ip/usart_gate.v(671)
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'b0000010010001100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD3CB0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [3]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [4]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA22E0 ));  // al_ip/usart_gate.v(747)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'b0000001000000111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD4530  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [6]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [6]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E9D0 ));  // al_ip/usart_gate.v(642)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~(~C*~B)))"),
    .INIT(32'b10101010101010101010101000000010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD4640  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E190 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EA80 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E9D0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [6]));  // al_ip/usart_gate.v(651)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111001101010000000000000101),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD4860  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FDC0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [7]));  // al_ip/usart_gate.v(613)
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'b0000010010001100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD5740  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F790 ));  // al_ip/usart_gate.v(575)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111000010111111011100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD5960  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [6]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E190 ));  // al_ip/usart_gate.v(623)
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'b0000010010001100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD5A70  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F0B0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [4]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EF50 ));  // al_ip/usart_gate.v(709)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'b0000001000000111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD5C90  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FD10 ));  // al_ip/usart_gate.v(584)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111000010111111011100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD5DA0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [4]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EEA0 ));  // al_ip/usart_gate.v(699)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~(~C*~B)))"),
    .INIT(32'b10101010101010101010101000000010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD5EB0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EB30 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EBE0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EC90 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [5]));  // al_ip/usart_gate.v(689)
  AL_MAP_LUT5 #(
    .EQN("((B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)*~(E)*~(D)+(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)*E*~(D)+~((B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))*E*D+(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)*E*D)"),
    .INIT(32'b11111111101011000000000010101100),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD62F0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA63600 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA60730 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [1]));  // al_ip/usart_gate.v(555)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111000010111111011100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6510  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [5]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [6]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EB30 ));  // al_ip/usart_gate.v(661)
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'b0000001000000111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6620  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [4]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [4]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1AA0 ));  // al_ip/usart_gate.v(718)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~(~C*~B)))"),
    .INIT(32'b10101010101010101010101000000010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6730  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EEA0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9EF50 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1AA0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [4]));  // al_ip/usart_gate.v(727)
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'b11111111000010111111011100000011),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6840  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E030 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [3]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AAAC0 [4]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA1100 ));  // al_ip/usart_gate.v(737)
  AL_MAP_LUT5 #(
    .EQN("(A*~(~E*~D*~(~C*~B)))"),
    .INIT(32'b10101010101010101010101000000010),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6B70  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E0E0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F790 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FD10 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A86E0 [0]));  // al_ip/usart_gate.v(593)
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'b0110))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6C80  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 [1]));  // al_ip/usart_gate.v(861)
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'b00000010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD6FB0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ));  // al_ip/usart_gate.v(954)
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(B*~(D*~C)))"),
    .INIT(16'b1110101011101110))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD72E0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4480 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5B30 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D3FB0 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5BE0 ));  // al_ip/usart_gate.v(918)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'b1000000000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD73F0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A832EE0 ));  // al_ip/usart_gate.v(936)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'b1000000000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7500  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55CB30 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C95E0 ));  // al_ip/usart_gate.v(978)
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'b1000000000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7610  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DAB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C8350 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DB60 ));  // al_ip/usart_gate.v(1003)
  AL_MAP_LUT4 #(
    .EQN("(D*~((~C*B))*~(A)+D*(~C*B)*~(A)+~(D)*(~C*B)*A+D*(~C*B)*A)"),
    .INIT(16'b0101110100001000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7720  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCA20 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CC810 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB420 ));  // al_ip/usart_gate.v(994)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7940  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [0]));  // al_ip/usart_gate.v(854)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'b1000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7A50  (
    .a(\u_PERIPH_TOP/u_USART2RIB/tx_en ),
    .b(\u_PERIPH_TOP/u_USART2RIB/tx_rdy ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D1E00 ));  // al_ip/usart_gate.v(875)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7B60  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [5]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [5]));  // al_ip/usart_gate.v(819)
  AL_MAP_LUT4 #(
    .EQN("~(D@C@B@A)"),
    .INIT(16'b1001011001101001))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7C70  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [6]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [7]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E500 ));  // al_ip/usart_gate.v(890)
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~C)*~(A)*~(B)+~(D*~C)*A*~(B)+~(~(D*~C))*A*B+~(D*~C)*A*B)"),
    .INIT(16'b0100011101000100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7D80  (
    .a(\u_PERIPH_TOP/u_USART2RIB/tx_en ),
    .b(\u_PERIPH_TOP/u_USART2RIB/tx_rdy ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D5B30 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D3FB0 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4320 ));  // al_ip/usart_gate.v(927)
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'b10100010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD7E90  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA03F0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB840 ));  // al_ip/usart_gate.v(1021)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD81C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [4]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [4]));  // al_ip/usart_gate.v(826)
  AL_MAP_LUT4 #(
    .EQN("(B*~((D@C))*~(A)+B*(D@C)*~(A)+~(B)*(D@C)*A+B*(D@C)*A)"),
    .INIT(16'b0100111011100100))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8600  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DB60 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCD90 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD470 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCA20 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAA03F0 ));  // al_ip/usart_gate.v(1012)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'b0000001000000000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8710  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A87C0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4480 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ));  // al_ip/usart_gate.v(1029)
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'b0000000000000001))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8820  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A8980 [3]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A68B0 [0]));  // al_ip/usart_gate.v(1047)
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'b1111101100000010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8930  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D3FB0 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D4C10 ));  // al_ip/usart_gate.v(909)
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'b0101111100001000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8A40  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C93D0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [0]),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_vld ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A550340 ));  // al_ip/usart_gate.v(945)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'b1000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8D70  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702AB0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F210 ));  // al_ip/usart_gate.v(1056)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8E80  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [1]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A55C970 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DAB0 ));  // al_ip/usart_gate.v(962)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'b1000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD8F90  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8C95E0 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A702530 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A832AC0 ));  // al_ip/usart_gate.v(987)
  AL_MAP_LUT5 #(
    .EQN("~(E@D@C@B@A)"),
    .INIT(32'b01101001100101101001011001101001),
    .LOC("UNPLACED"))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD90A0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9E500 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [2]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [3]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [4]),
    .e(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8AA190 [5]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2010 ));  // al_ip/usart_gate.v(899)
  AL_MAP_LUT4 #(
    .EQN("~(~D*C*B*A)"),
    .INIT(16'b1111111101111111))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD91B0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A68B0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9F210 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8D2F30 ));  // al_ip/usart_gate.v(1063)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD92C0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [3]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [3]));  // al_ip/usart_gate.v(833)
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'b0000000000000010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD93D0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DD70 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [0]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [1]),
    .d(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8A4BD0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CD890 ));  // al_ip/usart_gate.v(1038)
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'b01111000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD95F0  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [0]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [1]),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54CDE0 [2]),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54FF50 [2]));  // al_ip/usart_gate.v(882)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD9920  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [1]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [1]));  // al_ip/usart_gate.v(847)
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'b0010))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD9C50  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F770 [2]),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A830D30 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A54F2A0 [2]));  // al_ip/usart_gate.v(840)
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'b1110))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD9D60  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CCD90 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CC810 ),
    .o(\u_PERIPH_TOP/u_USART2RIB/rx_err ));  // al_ip/usart_gate.v(868)
  AL_MAP_LUT4 #(
    .EQN("((D*~B)*~(A)*~(C)+(D*~B)*A*~(C)+~((D*~B))*A*C+(D*~B)*A*C)"),
    .INIT(16'b1010001110100000))
    \u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AAD9E70  (
    .a(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A550340 ),
    .b(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9FBB0 ),
    .c(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673AA9DAB0 ),
    .d(\u_PERIPH_TOP/u_USART2RIB/rx_vld ),
    .o(\u_PERIPH_TOP/u_USART2RIB/u_USART/al_000002673A8CB2C0 ));  // al_ip/usart_gate.v(969)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_internal_reset/reg0_b0  (
    .clk(i_clk_pad),
    .d(1'b1),
    .sr(n1),
    .q(\u_internal_reset/synch_regs_q [0]));  // ../RTL/core/reset.v(16)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_internal_reset/reg0_b1  (
    .clk(i_clk_pad),
    .d(\u_internal_reset/synch_regs_q [0]),
    .sr(n1),
    .q(\u_internal_reset/synch_regs_q [1]));  // ../RTL/core/reset.v(16)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_internal_reset/reg0_b2  (
    .clk(i_clk_pad),
    .d(\u_internal_reset/synch_regs_q [1]),
    .sr(n1),
    .q(\u_internal_reset/synch_regs_q [2]));  // ../RTL/core/reset.v(16)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_internal_reset/reg0_b3  (
    .clk(i_clk_pad),
    .d(\u_internal_reset/synch_regs_q [2]),
    .sr(n1),
    .q(\u_internal_reset/synch_regs_q [3]));  // ../RTL/core/reset.v(16)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_internal_reset/reg0_b4  (
    .clk(i_clk_pad),
    .d(\u_internal_reset/synch_regs_q [3]),
    .sr(n1),
    .q(reset));  // ../RTL/core/reset.v(16)
  EG_PHY_GCLK \u_pll/bufg_feedback  (
    .clki(\u_pll/clk0_buf ),
    .clko(clk_84mhz_keep));  // al_ip/pll.v(34)
  EG_PHY_PLL #(
    .CLKC0_CPHASE(11),
    .CLKC0_DIV(12),
    .CLKC0_DIV2_ENABLE("DISABLE"),
    .CLKC0_ENABLE("ENABLE"),
    .CLKC0_FPHASE(0),
    .CLKC1_CPHASE(1),
    .CLKC1_DIV(1),
    .CLKC1_DIV2_ENABLE("DISABLE"),
    .CLKC1_ENABLE("DISABLE"),
    .CLKC1_FPHASE(0),
    .CLKC2_CPHASE(1),
    .CLKC2_DIV(1),
    .CLKC2_DIV2_ENABLE("DISABLE"),
    .CLKC2_ENABLE("DISABLE"),
    .CLKC2_FPHASE(0),
    .CLKC3_CPHASE(1),
    .CLKC3_DIV(1),
    .CLKC3_DIV2_ENABLE("DISABLE"),
    .CLKC3_ENABLE("DISABLE"),
    .CLKC3_FPHASE(0),
    .CLKC4_CPHASE(1),
    .CLKC4_DIV(1),
    .CLKC4_DIV2_ENABLE("DISABLE"),
    .CLKC4_ENABLE("DISABLE"),
    .CLKC4_FPHASE(0),
    .DERIVE_PLL_CLOCKS("DISABLE"),
    .DPHASE_SOURCE("DISABLE"),
    .DYNCFG("DISABLE"),
    .FBCLK_DIV(7),
    .FEEDBK_MODE("NORMAL"),
    .FEEDBK_PATH("CLKC0_EXT"),
    .FIN("24.000"),
    .FREQ_LOCK_ACCURACY(2),
    .GEN_BASIC_CLOCK("DISABLE"),
    .GMC_GAIN(0),
    .GMC_TEST(14),
    .ICP_CURRENT(9),
    .IF_ESCLKSTSW("DISABLE"),
    .INTFB_WAKE("DISABLE"),
    .KVCO(2),
    .LPF_CAPACITOR(2),
    .LPF_RESISTOR(8),
    .NORESET("DISABLE"),
    .ODIV_MUXC0("DIV"),
    .ODIV_MUXC1("DIV"),
    .ODIV_MUXC2("DIV"),
    .ODIV_MUXC3("DIV"),
    .ODIV_MUXC4("DIV"),
    .PLLC2RST_ENA("DISABLE"),
    .PLLC34RST_ENA("DISABLE"),
    .PLLMRST_ENA("DISABLE"),
    .PLLRST_ENA("ENABLE"),
    .PLL_LOCK_MODE(0),
    .PREDIV_MUXC0("VCO"),
    .PREDIV_MUXC1("VCO"),
    .PREDIV_MUXC2("VCO"),
    .PREDIV_MUXC3("VCO"),
    .PREDIV_MUXC4("VCO"),
    .REFCLK_DIV(2),
    .REFCLK_SEL("INTERNAL"),
    .STDBY_ENABLE("DISABLE"),
    .STDBY_VCO_ENA("DISABLE"),
    .SYNC_ENABLE("DISABLE"),
    .VCO_NORESET("DISABLE"))
    \u_pll/pll_inst  (
    .daddr(6'b000000),
    .dclk(1'b0),
    .dcs(1'b0),
    .di(8'b00000000),
    .dwe(1'b0),
    .fbclk(clk_84mhz),
    .load_reg(1'b0),
    .psclk(1'b0),
    .psclksel(3'b000),
    .psdown(1'b0),
    .psstep(1'b0),
    .refclk(i_clk_pad),
    .reset(n0),
    .stdby(1'b0),
    .clkc({open_n1233,open_n1234,open_n1235,open_n1236,\u_pll/clk0_buf }),
    .extlock(extlock));  // al_ip/pll.v(57)

endmodule 

module AL_BUFKEEP
  (
  i,
  o
  );

  input i;
  output o;

  parameter KEEP = "OUT";

  buf u1 (o, i);

endmodule 

module CORE_TOP  // ../RTL/soc_top/core_top.v(8)
  (
  i_clk,
  i_ribp_gnt,
  i_ribp_rdata,
  i_ribp_rsp,
  i_ribx_gnt,
  i_ribx_rdata,
  i_ribx_rsp,
  i_rstn,
  o_ribp_addr,
  o_ribp_mask,
  o_ribp_rdy,
  o_ribp_req,
  o_ribp_wdata,
  o_ribp_wrcs,
  o_ribx_addr,
  o_ribx_mask,
  o_ribx_rdy,
  o_ribx_req,
  o_ribx_wdata,
  o_ribx_wrcs
  );

  input i_clk;  // ../RTL/soc_top/core_top.v(9)
  input i_ribp_gnt;  // ../RTL/soc_top/core_top.v(31)
  input [31:0] i_ribp_rdata;  // ../RTL/soc_top/core_top.v(29)
  input i_ribp_rsp;  // ../RTL/soc_top/core_top.v(32)
  input i_ribx_gnt;  // ../RTL/soc_top/core_top.v(19)
  input [31:0] i_ribx_rdata;  // ../RTL/soc_top/core_top.v(17)
  input i_ribx_rsp;  // ../RTL/soc_top/core_top.v(20)
  input i_rstn;  // ../RTL/soc_top/core_top.v(10)
  output [31:0] o_ribp_addr;  // ../RTL/soc_top/core_top.v(25)
  output [3:0] o_ribp_mask;  // ../RTL/soc_top/core_top.v(27)
  output o_ribp_rdy;  // ../RTL/soc_top/core_top.v(33)
  output o_ribp_req;  // ../RTL/soc_top/core_top.v(30)
  output [31:0] o_ribp_wdata;  // ../RTL/soc_top/core_top.v(28)
  output o_ribp_wrcs;  // ../RTL/soc_top/core_top.v(26)
  output [31:0] o_ribx_addr;  // ../RTL/soc_top/core_top.v(13)
  output [3:0] o_ribx_mask;  // ../RTL/soc_top/core_top.v(15)
  output o_ribx_rdy;  // ../RTL/soc_top/core_top.v(21)
  output o_ribx_req;  // ../RTL/soc_top/core_top.v(18)
  output [31:0] o_ribx_wdata;  // ../RTL/soc_top/core_top.v(16)
  output o_ribx_wrcs;  // ../RTL/soc_top/core_top.v(14)

  wire [1:0] \RIB_ARB0/sel_tag ;  // ../RTL/core/rib.v(78)
  wire [7:0] \RIB_ARB0/sel_tag_id ;  // ../RTL/core/rib.v(113)
  wire [1:0] \RIB_ARB1/n7 ;
  wire [7:0] \RIB_ARB1/sel_tag_id ;  // ../RTL/core/rib.v(113)
  wire [1:0] \RIB_ARB2/sel_tag_id ;  // ../RTL/core/rib.v(252)
  wire [31:0] arb2_addr0;  // ../RTL/soc_top/core_top.v(241)
  wire [0:0] arb2_addr0_piped;
  wire [31:0] arb2_wdata0;  // ../RTL/soc_top/core_top.v(244)
  wire [31:0] rib_addr0;  // ../RTL/soc_top/core_top.v(37)
  wire [31:0] rib_addr1;  // ../RTL/soc_top/core_top.v(48)
  wire [0:1] rib_addr1_piped;
  wire [3:0] rib_mask1;  // ../RTL/soc_top/core_top.v(50)
  wire [31:0] rib_rdata0;  // ../RTL/soc_top/core_top.v(41)
  wire [31:0] rib_rdata1;  // ../RTL/soc_top/core_top.v(52)
  wire [31:0] rib_wdata1;  // ../RTL/soc_top/core_top.v(51)
  wire [3:0] \u_DTCM_CTRL/bram_wea ;  // ../RTL/periph/bram2rib.v(27)
  wire [3:0] \u_ITCM_CTRL/bram_wea ;  // ../RTL/periph/bram2rib.v(98)
  wire \RIB_ARB0/default_cs ;  // ../RTL/core/rib.v(112)
  wire \RIB_ARB0/handshake_rdy_last ;  // ../RTL/core/rib.v(117)
  wire \RIB_ARB0/mux3_b0_sel_is_0_o ;
  wire \RIB_ARB0/n3 ;
  wire \RIB_ARB0/n6 ;
  wire \RIB_ARB1/default_cs ;  // ../RTL/core/rib.v(112)
  wire \RIB_ARB1/handshake_rdy_last ;  // ../RTL/core/rib.v(117)
  wire \RIB_ARB1/n3 ;
  wire \RIB_ARB1/n6 ;
  wire \RIB_ARB2/handshake_rdy_last ;  // ../RTL/core/rib.v(256)
  wire _al_u186_o;
  wire _al_u187_o;
  wire _al_u188_o;
  wire _al_u189_o;
  wire _al_u191_o;
  wire _al_u192_o;
  wire _al_u193_o;
  wire _al_u195_o;
  wire _al_u196_o;
  wire _al_u197_o;
  wire _al_u199_o;
  wire _al_u200_o;
  wire _al_u201_o;
  wire _al_u203_o;
  wire _al_u204_o;
  wire _al_u205_o;
  wire _al_u207_o;
  wire _al_u208_o;
  wire _al_u209_o;
  wire _al_u211_o;
  wire _al_u212_o;
  wire _al_u213_o;
  wire _al_u215_o;
  wire _al_u216_o;
  wire _al_u217_o;
  wire _al_u219_o;
  wire _al_u220_o;
  wire _al_u221_o;
  wire _al_u223_o;
  wire _al_u224_o;
  wire _al_u225_o;
  wire _al_u227_o;
  wire _al_u228_o;
  wire _al_u229_o;
  wire _al_u231_o;
  wire _al_u232_o;
  wire _al_u233_o;
  wire _al_u235_o;
  wire _al_u236_o;
  wire _al_u237_o;
  wire _al_u239_o;
  wire _al_u240_o;
  wire _al_u241_o;
  wire _al_u243_o;
  wire _al_u244_o;
  wire _al_u245_o;
  wire _al_u247_o;
  wire _al_u248_o;
  wire _al_u249_o;
  wire _al_u251_o;
  wire _al_u252_o;
  wire _al_u253_o;
  wire _al_u255_o;
  wire _al_u256_o;
  wire _al_u257_o;
  wire _al_u259_o;
  wire _al_u260_o;
  wire _al_u261_o;
  wire _al_u263_o;
  wire _al_u264_o;
  wire _al_u265_o;
  wire _al_u267_o;
  wire _al_u268_o;
  wire _al_u269_o;
  wire _al_u271_o;
  wire _al_u272_o;
  wire _al_u273_o;
  wire _al_u275_o;
  wire _al_u276_o;
  wire _al_u277_o;
  wire _al_u279_o;
  wire _al_u280_o;
  wire _al_u281_o;
  wire _al_u283_o;
  wire _al_u284_o;
  wire _al_u285_o;
  wire _al_u287_o;
  wire _al_u288_o;
  wire _al_u289_o;
  wire _al_u291_o;
  wire _al_u292_o;
  wire _al_u293_o;
  wire _al_u295_o;
  wire _al_u296_o;
  wire _al_u297_o;
  wire _al_u299_o;
  wire _al_u300_o;
  wire _al_u301_o;
  wire _al_u303_o;
  wire _al_u304_o;
  wire _al_u305_o;
  wire _al_u307_o;
  wire _al_u308_o;
  wire _al_u309_o;
  wire _al_u311_o;
  wire _al_u312_o;
  wire _al_u313_o;
  wire _al_u315_o;
  wire _al_u316_o;
  wire _al_u319_o;
  wire _al_u320_o;
  wire _al_u321_o;
  wire \and_Nrib_addr1[14]_N_o ;
  wire \and_Nrib_addr1[14]_r_o ;
  wire \and_rib_addr1[14]_Nr_o ;
  wire \and_rib_addr1[14]_ri_o ;
  wire arb0_gnt0;  // ../RTL/soc_top/core_top.v(95)
  wire arb0_rsp0;  // ../RTL/soc_top/core_top.v(96)
  wire arb1_req0;  // ../RTL/soc_top/core_top.v(164)
  wire arb1_req1;  // ../RTL/soc_top/core_top.v(174)
  wire arb1_rsp1;  // ../RTL/soc_top/core_top.v(176)
  wire arb2_req0;  // ../RTL/soc_top/core_top.v(246)
  wire rib_gnt1;  // ../RTL/soc_top/core_top.v(54)
  wire rib_req0;  // ../RTL/soc_top/core_top.v(42)
  wire rib_req1;  // ../RTL/soc_top/core_top.v(53)
  wire rib_rsp1;  // ../RTL/soc_top/core_top.v(55)
  wire rib_wrcs1;  // ../RTL/soc_top/core_top.v(49)
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_000 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_001 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_002 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_003 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_004 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_005 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_006 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_007 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_008 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_009 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_010 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_011 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_012 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_013 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_014 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_015 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_016 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_017 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_018 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_019 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_020 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_021 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_022 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_023 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_024 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_025 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_026 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_027 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_028 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_029 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_030 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_031 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_000 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_001 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_002 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_003 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_004 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_005 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_006 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_007 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_008 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_009 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_010 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_011 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_012 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_013 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_014 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_015 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_016 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_017 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_018 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_019 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_020 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_021 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_022 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_023 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_024 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_025 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_026 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_027 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_028 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_029 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_030 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_031 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_000 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_001 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_002 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_003 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_004 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_005 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_006 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_007 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_008 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_009 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_010 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_011 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_012 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_013 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_014 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_015 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_016 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_017 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_018 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_019 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_020 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_021 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_022 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_023 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_024 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_025 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_026 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_027 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_028 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_029 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_030 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_031 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_000 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_001 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_002 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_003 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_004 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_005 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_006 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_007 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_008 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_009 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_010 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_011 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_012 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_013 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_014 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_015 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_016 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_017 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_018 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_019 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_020 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_021 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_022 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_023 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_024 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_025 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_026 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_027 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_028 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_029 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_030 ;
  wire \u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_031 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_000 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_001 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_002 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_003 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_004 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_005 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_006 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_007 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_008 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_009 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_010 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_011 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_012 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_013 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_014 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_015 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_016 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_017 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_018 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_019 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_020 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_021 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_022 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_023 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_024 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_025 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_026 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_027 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_028 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_029 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_030 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_031 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_000 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_001 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_002 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_003 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_004 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_005 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_006 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_007 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_008 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_009 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_010 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_011 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_012 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_013 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_014 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_015 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_016 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_017 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_018 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_019 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_020 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_021 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_022 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_023 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_024 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_025 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_026 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_027 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_028 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_029 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_030 ;
  wire \u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_031 ;

  assign o_ribp_addr[31] = rib_addr1[31];
  assign o_ribp_addr[30] = rib_addr1[30];
  assign o_ribp_addr[29] = rib_addr1[29];
  assign o_ribp_addr[28] = rib_addr1[28];
  assign o_ribp_addr[27] = rib_addr1[27];
  assign o_ribp_addr[26] = rib_addr1[26];
  assign o_ribp_addr[25] = rib_addr1[25];
  assign o_ribp_addr[24] = rib_addr1[24];
  assign o_ribp_addr[15] = rib_addr1[15];
  assign o_ribp_addr[14] = rib_addr1[14];
  assign o_ribp_addr[13] = rib_addr1[13];
  assign o_ribp_addr[12] = rib_addr1[12];
  assign o_ribp_addr[11] = rib_addr1[11];
  assign o_ribp_addr[10] = rib_addr1[10];
  assign o_ribp_addr[9] = rib_addr1[9];
  assign o_ribp_addr[8] = rib_addr1[8];
  assign o_ribp_addr[7] = rib_addr1[7];
  assign o_ribp_addr[6] = rib_addr1[6];
  assign o_ribp_addr[5] = rib_addr1[5];
  assign o_ribp_addr[4] = rib_addr1[4];
  assign o_ribp_addr[3] = rib_addr1[3];
  assign o_ribp_addr[2] = rib_addr1[2];
  assign o_ribp_addr[1] = 1'b0;
  assign o_ribp_addr[0] = 1'b0;
  assign o_ribp_mask[3] = rib_mask1[3];
  assign o_ribp_mask[2] = rib_mask1[2];
  assign o_ribp_mask[1] = rib_mask1[1];
  assign o_ribp_mask[0] = rib_mask1[0];
  assign o_ribp_wdata[31] = rib_wdata1[31];
  assign o_ribp_wdata[30] = rib_wdata1[30];
  assign o_ribp_wdata[29] = rib_wdata1[29];
  assign o_ribp_wdata[28] = rib_wdata1[28];
  assign o_ribp_wdata[27] = rib_wdata1[27];
  assign o_ribp_wdata[26] = rib_wdata1[26];
  assign o_ribp_wdata[25] = rib_wdata1[25];
  assign o_ribp_wdata[24] = rib_wdata1[24];
  assign o_ribp_wdata[23] = rib_wdata1[23];
  assign o_ribp_wdata[22] = rib_wdata1[22];
  assign o_ribp_wdata[21] = rib_wdata1[21];
  assign o_ribp_wdata[20] = rib_wdata1[20];
  assign o_ribp_wdata[19] = rib_wdata1[19];
  assign o_ribp_wdata[18] = rib_wdata1[18];
  assign o_ribp_wdata[17] = rib_wdata1[17];
  assign o_ribp_wdata[16] = rib_wdata1[16];
  assign o_ribp_wdata[15] = rib_wdata1[15];
  assign o_ribp_wdata[14] = rib_wdata1[14];
  assign o_ribp_wdata[13] = rib_wdata1[13];
  assign o_ribp_wdata[12] = rib_wdata1[12];
  assign o_ribp_wdata[11] = rib_wdata1[11];
  assign o_ribp_wdata[10] = rib_wdata1[10];
  assign o_ribp_wdata[9] = rib_wdata1[9];
  assign o_ribp_wdata[8] = rib_wdata1[8];
  assign o_ribp_wdata[7] = rib_wdata1[7];
  assign o_ribp_wdata[6] = rib_wdata1[6];
  assign o_ribp_wdata[5] = rib_wdata1[5];
  assign o_ribp_wdata[4] = rib_wdata1[4];
  assign o_ribp_wdata[3] = rib_wdata1[3];
  assign o_ribp_wdata[2] = rib_wdata1[2];
  assign o_ribp_wdata[1] = rib_wdata1[1];
  assign o_ribp_wdata[0] = rib_wdata1[0];
  assign o_ribp_wrcs = rib_wrcs1;
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("SET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \RIB_ARB0/default_cs_reg  (
    .ce(\RIB_ARB0/n6 ),
    .clk(i_clk),
    .d(\RIB_ARB0/n3 ),
    .sr(i_rstn),
    .q(\RIB_ARB0/default_cs ));  // ../RTL/core/rib.v(121)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \RIB_ARB0/handshake_rdy_last_reg  (
    .ce(\RIB_ARB0/n6 ),
    .clk(i_clk),
    .d(arb0_gnt0),
    .sr(i_rstn),
    .q(\RIB_ARB0/handshake_rdy_last ));  // ../RTL/core/rib.v(121)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \RIB_ARB0/reg0_b0  (
    .ce(\RIB_ARB0/n6 ),
    .clk(i_clk),
    .d(\RIB_ARB0/sel_tag [1]),
    .sr(i_rstn),
    .q(\RIB_ARB0/sel_tag_id [0]));  // ../RTL/core/rib.v(121)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("SET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \RIB_ARB1/default_cs_reg  (
    .ce(\RIB_ARB1/n6 ),
    .clk(i_clk),
    .d(\RIB_ARB1/n3 ),
    .sr(i_rstn),
    .q(\RIB_ARB1/default_cs ));  // ../RTL/core/rib.v(121)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \RIB_ARB1/handshake_rdy_last_reg  (
    .ce(\RIB_ARB1/n6 ),
    .clk(i_clk),
    .d(rib_gnt1),
    .sr(i_rstn),
    .q(\RIB_ARB1/handshake_rdy_last ));  // ../RTL/core/rib.v(121)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \RIB_ARB1/reg0_b0  (
    .ce(\RIB_ARB1/n6 ),
    .clk(i_clk),
    .d(\RIB_ARB1/n7 [0]),
    .sr(i_rstn),
    .q(\RIB_ARB1/sel_tag_id [0]));  // ../RTL/core/rib.v(121)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \RIB_ARB1/reg0_b1  (
    .ce(\RIB_ARB1/n6 ),
    .clk(i_clk),
    .d(\RIB_ARB1/n7 [1]),
    .sr(i_rstn),
    .q(\RIB_ARB1/sel_tag_id [1]));  // ../RTL/core/rib.v(121)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \RIB_ARB2/handshake_rdy_last_reg  (
    .clk(i_clk),
    .d(arb2_req0),
    .sr(i_rstn),
    .q(\RIB_ARB2/handshake_rdy_last ));  // ../RTL/core/rib.v(260)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \RIB_ARB2/reg0_b0  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(arb1_req0),
    .q(\RIB_ARB2/sel_tag_id [0]));  // ../RTL/core/rib.v(260)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u145 (
    .a(rib_addr1[15]),
    .b(rib_addr1[14]),
    .o(\and_rib_addr1[14]_ri_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u146 (
    .a(rib_addr1[15]),
    .b(rib_addr1[14]),
    .o(\and_rib_addr1[14]_Nr_o ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u147 (
    .a(rib_addr1[15]),
    .b(rib_addr1[14]),
    .o(\and_Nrib_addr1[14]_r_o ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u148 (
    .a(rib_addr1[15]),
    .b(rib_addr1[14]),
    .o(\and_Nrib_addr1[14]_N_o ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u149 (
    .a(\RIB_ARB2/handshake_rdy_last ),
    .b(\RIB_ARB2/sel_tag_id [0]),
    .o(arb0_rsp0));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u150 (
    .a(\RIB_ARB0/default_cs ),
    .b(\RIB_ARB0/sel_tag_id [0]),
    .o(\RIB_ARB0/mux3_b0_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u151 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_009 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_009 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[9]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u152 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_008 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_008 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[8]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u153 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_007 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_007 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[7]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u154 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_006 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_006 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[6]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u155 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_005 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_005 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[5]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u156 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_004 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_004 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[4]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u157 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_003 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_003 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[3]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u158 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_031 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_031 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[31]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u159 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_030 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_030 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[30]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u160 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_002 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_002 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[2]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u161 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_029 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_029 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[29]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u162 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_028 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_028 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[28]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u163 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_027 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_027 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[27]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u164 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_026 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_026 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[26]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u165 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_025 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_025 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[25]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u166 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_024 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_024 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[24]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u167 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_023 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_023 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[23]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u168 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_022 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_022 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[22]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u169 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_021 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_021 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[21]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u170 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_020 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_020 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[20]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u171 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_001 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_001 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[1]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u172 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_019 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_019 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[19]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u173 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_018 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_018 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[18]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u174 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_017 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_017 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[17]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u175 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_016 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_016 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[16]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u176 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_015 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_015 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[15]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u177 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_014 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_014 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[14]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u178 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_013 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_013 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[13]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u179 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_012 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_012 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[12]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u180 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_011 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_011 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[11]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u181 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_010 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_010 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[10]));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u182 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_000 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_000 ),
    .c(\RIB_ARB0/mux3_b0_sel_is_0_o ),
    .d(arb2_addr0_piped),
    .o(rib_rdata0[0]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~A*~(C*B))"),
    .INIT(16'hffea))
    _al_u183 (
    .a(i_ribp_rsp),
    .b(\RIB_ARB2/handshake_rdy_last ),
    .c(\RIB_ARB2/sel_tag_id [0]),
    .d(arb1_rsp1),
    .o(rib_rsp1));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u184 (
    .a(arb0_rsp0),
    .b(\RIB_ARB0/handshake_rdy_last ),
    .o(\RIB_ARB0/n6 ));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u185 (
    .a(rib_rsp1),
    .b(\RIB_ARB1/handshake_rdy_last ),
    .o(\RIB_ARB1/n6 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u186 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_007 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_007 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_007 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u186_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u187 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_007 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u187_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u188 (
    .a(\RIB_ARB1/default_cs ),
    .b(\RIB_ARB1/sel_tag_id [1]),
    .o(_al_u188_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u189 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_007 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_007 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u189_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u190 (
    .a(_al_u186_o),
    .b(_al_u187_o),
    .c(_al_u189_o),
    .d(i_ribp_rdata[7]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[7]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u191 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_006 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_006 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_006 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u191_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u192 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_006 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u192_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u193 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_006 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_006 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u193_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u194 (
    .a(_al_u191_o),
    .b(_al_u192_o),
    .c(_al_u193_o),
    .d(i_ribp_rdata[6]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[6]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u195 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_005 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_005 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_005 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u195_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u196 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_005 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u196_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u197 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_005 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_005 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u197_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u198 (
    .a(_al_u195_o),
    .b(_al_u196_o),
    .c(_al_u197_o),
    .d(i_ribp_rdata[5]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[5]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u199 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_004 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_004 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_004 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u199_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u200 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_004 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u200_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u201 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_004 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_004 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u201_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u202 (
    .a(_al_u199_o),
    .b(_al_u200_o),
    .c(_al_u201_o),
    .d(i_ribp_rdata[4]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[4]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u203 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_003 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_003 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_003 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u203_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u204 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_003 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u204_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u205 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_003 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_003 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u205_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u206 (
    .a(_al_u203_o),
    .b(_al_u204_o),
    .c(_al_u205_o),
    .d(i_ribp_rdata[3]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[3]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u207 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_002 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_002 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_002 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u207_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u208 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_002 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u208_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u209 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_002 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_002 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u209_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u210 (
    .a(_al_u207_o),
    .b(_al_u208_o),
    .c(_al_u209_o),
    .d(i_ribp_rdata[2]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[2]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u211 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_001 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_001 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_001 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u211_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u212 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_001 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u212_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u213 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_001 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_001 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u213_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u214 (
    .a(_al_u211_o),
    .b(_al_u212_o),
    .c(_al_u213_o),
    .d(i_ribp_rdata[1]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[1]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u215 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_000 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_000 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_000 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u215_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u216 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_000 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u216_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u217 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_000 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_000 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u217_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u218 (
    .a(_al_u215_o),
    .b(_al_u216_o),
    .c(_al_u217_o),
    .d(i_ribp_rdata[0]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[0]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u219 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_015 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_015 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_015 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u219_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u220 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_015 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u220_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u221 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_015 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_015 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u221_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u222 (
    .a(_al_u219_o),
    .b(_al_u220_o),
    .c(_al_u221_o),
    .d(i_ribp_rdata[15]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[15]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u223 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_014 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_014 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_014 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u223_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u224 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_014 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u224_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u225 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_014 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_014 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u225_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u226 (
    .a(_al_u223_o),
    .b(_al_u224_o),
    .c(_al_u225_o),
    .d(i_ribp_rdata[14]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[14]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u227 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_013 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_013 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_013 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u227_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u228 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_013 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u228_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u229 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_013 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_013 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u229_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u230 (
    .a(_al_u227_o),
    .b(_al_u228_o),
    .c(_al_u229_o),
    .d(i_ribp_rdata[13]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[13]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u231 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_012 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_012 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_012 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u231_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u232 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_012 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u232_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u233 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_012 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_012 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u233_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u234 (
    .a(_al_u231_o),
    .b(_al_u232_o),
    .c(_al_u233_o),
    .d(i_ribp_rdata[12]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[12]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u235 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_011 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_011 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_011 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u235_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u236 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_011 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u236_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u237 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_011 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_011 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u237_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u238 (
    .a(_al_u235_o),
    .b(_al_u236_o),
    .c(_al_u237_o),
    .d(i_ribp_rdata[11]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[11]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u239 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_010 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_010 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_010 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u239_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u240 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_010 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u240_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u241 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_010 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_010 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u241_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u242 (
    .a(_al_u239_o),
    .b(_al_u240_o),
    .c(_al_u241_o),
    .d(i_ribp_rdata[10]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[10]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u243 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_009 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_009 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_009 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u243_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u244 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_009 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u244_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u245 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_009 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_009 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u245_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u246 (
    .a(_al_u243_o),
    .b(_al_u244_o),
    .c(_al_u245_o),
    .d(i_ribp_rdata[9]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[9]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u247 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_008 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_008 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_008 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u247_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u248 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_008 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u248_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u249 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_008 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_008 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u249_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u250 (
    .a(_al_u247_o),
    .b(_al_u248_o),
    .c(_al_u249_o),
    .d(i_ribp_rdata[8]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[8]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u251 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_023 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_023 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_023 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u251_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u252 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_023 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u252_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u253 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_023 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_023 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u253_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u254 (
    .a(_al_u251_o),
    .b(_al_u252_o),
    .c(_al_u253_o),
    .d(i_ribp_rdata[23]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[23]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u255 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_022 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_022 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_022 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u255_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u256 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_022 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u256_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u257 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_022 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_022 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u257_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u258 (
    .a(_al_u255_o),
    .b(_al_u256_o),
    .c(_al_u257_o),
    .d(i_ribp_rdata[22]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[22]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u259 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_021 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_021 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_021 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u259_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u260 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_021 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u260_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u261 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_021 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_021 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u261_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u262 (
    .a(_al_u259_o),
    .b(_al_u260_o),
    .c(_al_u261_o),
    .d(i_ribp_rdata[21]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[21]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u263 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_020 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_020 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_020 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u263_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u264 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_020 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u264_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u265 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_020 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_020 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u265_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u266 (
    .a(_al_u263_o),
    .b(_al_u264_o),
    .c(_al_u265_o),
    .d(i_ribp_rdata[20]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[20]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u267 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_019 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_019 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_019 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u267_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u268 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_019 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u268_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u269 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_019 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_019 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u269_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u270 (
    .a(_al_u267_o),
    .b(_al_u268_o),
    .c(_al_u269_o),
    .d(i_ribp_rdata[19]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[19]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u271 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_018 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_018 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_018 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u271_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u272 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_018 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u272_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u273 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_018 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_018 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u273_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u274 (
    .a(_al_u271_o),
    .b(_al_u272_o),
    .c(_al_u273_o),
    .d(i_ribp_rdata[18]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[18]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u275 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_017 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_017 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_017 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u275_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u276 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_017 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u276_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u277 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_017 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_017 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u277_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u278 (
    .a(_al_u275_o),
    .b(_al_u276_o),
    .c(_al_u277_o),
    .d(i_ribp_rdata[17]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[17]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u279 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_016 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_016 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_016 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u279_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u280 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_016 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u280_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u281 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_016 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_016 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u281_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u282 (
    .a(_al_u279_o),
    .b(_al_u280_o),
    .c(_al_u281_o),
    .d(i_ribp_rdata[16]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[16]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u283 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_031 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_031 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_031 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u283_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u284 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_031 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u284_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u285 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_031 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_031 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u285_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u286 (
    .a(_al_u283_o),
    .b(_al_u284_o),
    .c(_al_u285_o),
    .d(i_ribp_rdata[31]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[31]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u287 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_030 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_030 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_030 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u287_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u288 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_030 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u288_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u289 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_030 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_030 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u289_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u290 (
    .a(_al_u287_o),
    .b(_al_u288_o),
    .c(_al_u289_o),
    .d(i_ribp_rdata[30]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[30]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u291 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_029 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_029 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_029 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u291_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u292 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_029 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u292_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u293 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_029 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_029 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u293_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u294 (
    .a(_al_u291_o),
    .b(_al_u292_o),
    .c(_al_u293_o),
    .d(i_ribp_rdata[29]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[29]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u295 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_028 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_028 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_028 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u295_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u296 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_028 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u296_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u297 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_028 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_028 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u297_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u298 (
    .a(_al_u295_o),
    .b(_al_u296_o),
    .c(_al_u297_o),
    .d(i_ribp_rdata[28]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[28]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u299 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_027 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_027 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_027 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u299_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u300 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_027 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u300_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u301 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_027 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_027 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u301_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u302 (
    .a(_al_u299_o),
    .b(_al_u300_o),
    .c(_al_u301_o),
    .d(i_ribp_rdata[27]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[27]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u303 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_026 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_026 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_026 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u303_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u304 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_026 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u304_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u305 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_026 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_026 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u305_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u306 (
    .a(_al_u303_o),
    .b(_al_u304_o),
    .c(_al_u305_o),
    .d(i_ribp_rdata[26]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[26]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u307 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_025 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_025 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_025 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u307_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u308 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_025 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u308_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u309 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_025 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_025 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u309_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u310 (
    .a(_al_u307_o),
    .b(_al_u308_o),
    .c(_al_u309_o),
    .d(i_ribp_rdata[25]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[25]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f3355ff))
    _al_u311 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_024 ),
    .b(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_024 ),
    .c(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_024 ),
    .d(rib_addr1_piped[0]),
    .e(rib_addr1_piped[1]),
    .o(_al_u311_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*A))"),
    .INIT(16'hccc4))
    _al_u312 (
    .a(\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_024 ),
    .b(\RIB_ARB1/sel_tag_id [0]),
    .c(rib_addr1_piped[0]),
    .d(rib_addr1_piped[1]),
    .o(_al_u312_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'hf0c0f0a0))
    _al_u313 (
    .a(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_024 ),
    .b(\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_024 ),
    .c(_al_u188_o),
    .d(\RIB_ARB1/sel_tag_id [0]),
    .e(arb2_addr0_piped),
    .o(_al_u313_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*D)*~(C*~(B*A)))"),
    .INIT(32'hff707070))
    _al_u314 (
    .a(_al_u311_o),
    .b(_al_u312_o),
    .c(_al_u313_o),
    .d(i_ribp_rdata[24]),
    .e(\RIB_ARB1/default_cs ),
    .o(rib_rdata1[24]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u315 (
    .a(rib_addr0[31]),
    .b(rib_addr0[30]),
    .o(_al_u315_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u316 (
    .a(rib_addr0[29]),
    .b(rib_addr0[28]),
    .c(rib_addr0[24]),
    .o(_al_u316_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*B*A)"),
    .INIT(16'hfff7))
    _al_u317 (
    .a(_al_u316_o),
    .b(_al_u315_o),
    .c(rib_addr0[27]),
    .d(rib_addr0[26]),
    .o(\RIB_ARB0/n3 ));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'h00080000))
    _al_u318 (
    .a(_al_u316_o),
    .b(_al_u315_o),
    .c(rib_addr0[27]),
    .d(rib_addr0[26]),
    .e(rib_addr0[25]),
    .o(\RIB_ARB0/sel_tag [1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u319 (
    .a(rib_addr1[31]),
    .b(rib_addr1[30]),
    .c(rib_addr1[29]),
    .d(rib_addr1[28]),
    .o(_al_u319_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u320 (
    .a(rib_addr1[27]),
    .b(rib_addr1[26]),
    .o(_al_u320_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u321 (
    .a(rib_addr1[27]),
    .b(rib_addr1[26]),
    .c(rib_addr1[25]),
    .o(_al_u321_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u322 (
    .a(_al_u319_o),
    .b(_al_u321_o),
    .c(rib_addr1[24]),
    .d(rib_req1),
    .o(arb1_req0));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u323 (
    .a(_al_u319_o),
    .b(_al_u320_o),
    .c(rib_addr1[25]),
    .d(rib_addr1[24]),
    .o(\RIB_ARB1/n7 [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u324 (
    .a(_al_u319_o),
    .b(_al_u321_o),
    .c(rib_addr1[24]),
    .o(\RIB_ARB1/n7 [0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u325 (
    .a(_al_u319_o),
    .b(_al_u321_o),
    .c(rib_addr1[24]),
    .d(rib_req1),
    .o(arb1_req1));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(~C*~B*A))"),
    .INIT(16'hff02))
    _al_u326 (
    .a(rib_req0),
    .b(\RIB_ARB0/n3 ),
    .c(rib_addr0[25]),
    .d(arb1_req0),
    .o(arb2_req0));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u327 (
    .a(arb1_req0),
    .b(rib_wdata1[9]),
    .o(arb2_wdata0[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u328 (
    .a(arb1_req0),
    .b(rib_wdata1[8]),
    .o(arb2_wdata0[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u329 (
    .a(arb1_req0),
    .b(rib_wdata1[7]),
    .o(arb2_wdata0[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u330 (
    .a(arb1_req0),
    .b(rib_wdata1[6]),
    .o(arb2_wdata0[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u331 (
    .a(arb1_req0),
    .b(rib_wdata1[5]),
    .o(arb2_wdata0[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u332 (
    .a(arb1_req0),
    .b(rib_wdata1[4]),
    .o(arb2_wdata0[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u333 (
    .a(arb1_req0),
    .b(rib_wdata1[31]),
    .o(arb2_wdata0[31]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u334 (
    .a(arb1_req0),
    .b(rib_wdata1[30]),
    .o(arb2_wdata0[30]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u335 (
    .a(arb1_req0),
    .b(rib_wdata1[3]),
    .o(arb2_wdata0[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u336 (
    .a(arb1_req0),
    .b(rib_wdata1[29]),
    .o(arb2_wdata0[29]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u337 (
    .a(arb1_req0),
    .b(rib_wdata1[28]),
    .o(arb2_wdata0[28]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u338 (
    .a(arb1_req0),
    .b(rib_wdata1[27]),
    .o(arb2_wdata0[27]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u339 (
    .a(arb1_req0),
    .b(rib_wdata1[26]),
    .o(arb2_wdata0[26]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u340 (
    .a(arb1_req0),
    .b(rib_wdata1[25]),
    .o(arb2_wdata0[25]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u341 (
    .a(arb1_req0),
    .b(rib_wdata1[24]),
    .o(arb2_wdata0[24]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u342 (
    .a(arb1_req0),
    .b(rib_wdata1[23]),
    .o(arb2_wdata0[23]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u343 (
    .a(arb1_req0),
    .b(rib_wdata1[22]),
    .o(arb2_wdata0[22]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u344 (
    .a(arb1_req0),
    .b(rib_wdata1[21]),
    .o(arb2_wdata0[21]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u345 (
    .a(arb1_req0),
    .b(rib_wdata1[20]),
    .o(arb2_wdata0[20]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u346 (
    .a(arb1_req0),
    .b(rib_wdata1[2]),
    .o(arb2_wdata0[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u347 (
    .a(arb1_req0),
    .b(rib_wdata1[19]),
    .o(arb2_wdata0[19]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u348 (
    .a(arb1_req0),
    .b(rib_wdata1[18]),
    .o(arb2_wdata0[18]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u349 (
    .a(arb1_req0),
    .b(rib_wdata1[17]),
    .o(arb2_wdata0[17]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u350 (
    .a(arb1_req0),
    .b(rib_wdata1[16]),
    .o(arb2_wdata0[16]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u351 (
    .a(arb1_req0),
    .b(rib_wdata1[15]),
    .o(arb2_wdata0[15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u352 (
    .a(arb1_req0),
    .b(rib_wdata1[14]),
    .o(arb2_wdata0[14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u353 (
    .a(arb1_req0),
    .b(rib_wdata1[13]),
    .o(arb2_wdata0[13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u354 (
    .a(arb1_req0),
    .b(rib_wdata1[12]),
    .o(arb2_wdata0[12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u355 (
    .a(arb1_req0),
    .b(rib_wdata1[11]),
    .o(arb2_wdata0[11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u356 (
    .a(arb1_req0),
    .b(rib_wdata1[10]),
    .o(arb2_wdata0[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u357 (
    .a(arb1_req0),
    .b(rib_wdata1[1]),
    .o(arb2_wdata0[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u358 (
    .a(arb1_req0),
    .b(rib_wdata1[0]),
    .o(arb2_wdata0[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u359 (
    .a(rib_addr0[9]),
    .b(arb1_req0),
    .c(rib_addr1[9]),
    .o(arb2_addr0[9]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u360 (
    .a(rib_addr0[8]),
    .b(arb1_req0),
    .c(rib_addr1[8]),
    .o(arb2_addr0[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u361 (
    .a(rib_addr0[7]),
    .b(arb1_req0),
    .c(rib_addr1[7]),
    .o(arb2_addr0[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u362 (
    .a(rib_addr0[6]),
    .b(arb1_req0),
    .c(rib_addr1[6]),
    .o(arb2_addr0[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u363 (
    .a(rib_addr0[5]),
    .b(arb1_req0),
    .c(rib_addr1[5]),
    .o(arb2_addr0[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u364 (
    .a(rib_addr0[4]),
    .b(arb1_req0),
    .c(rib_addr1[4]),
    .o(arb2_addr0[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u365 (
    .a(rib_addr0[3]),
    .b(arb1_req0),
    .c(rib_addr1[3]),
    .o(arb2_addr0[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u366 (
    .a(rib_addr0[2]),
    .b(arb1_req0),
    .c(rib_addr1[2]),
    .o(arb2_addr0[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u367 (
    .a(rib_addr0[15]),
    .b(arb1_req0),
    .c(rib_addr1[15]),
    .o(arb2_addr0[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u368 (
    .a(rib_addr0[14]),
    .b(arb1_req0),
    .c(rib_addr1[14]),
    .o(arb2_addr0[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u369 (
    .a(rib_addr0[13]),
    .b(arb1_req0),
    .c(rib_addr1[13]),
    .o(arb2_addr0[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u370 (
    .a(rib_addr0[12]),
    .b(arb1_req0),
    .c(rib_addr1[12]),
    .o(arb2_addr0[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u371 (
    .a(rib_addr0[11]),
    .b(arb1_req0),
    .c(rib_addr1[11]),
    .o(arb2_addr0[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u372 (
    .a(rib_addr0[10]),
    .b(arb1_req0),
    .c(rib_addr1[10]),
    .o(arb2_addr0[10]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u373 (
    .a(rib_req0),
    .b(\RIB_ARB0/n3 ),
    .c(rib_addr0[25]),
    .d(arb1_req0),
    .o(arb0_gnt0));
  AL_MAP_LUT4 #(
    .EQN("~(B*A*~(D*C))"),
    .INIT(16'hf777))
    _al_u374 (
    .a(_al_u319_o),
    .b(_al_u320_o),
    .c(rib_addr1[25]),
    .d(rib_addr1[24]),
    .o(\RIB_ARB1/n3 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u375 (
    .a(arb1_req1),
    .b(rib_mask1[3]),
    .c(rib_wrcs1),
    .o(\u_DTCM_CTRL/bram_wea [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u376 (
    .a(arb1_req1),
    .b(rib_mask1[2]),
    .c(rib_wrcs1),
    .o(\u_DTCM_CTRL/bram_wea [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u377 (
    .a(arb1_req1),
    .b(rib_mask1[1]),
    .c(rib_wrcs1),
    .o(\u_DTCM_CTRL/bram_wea [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u378 (
    .a(arb1_req1),
    .b(rib_mask1[0]),
    .c(rib_wrcs1),
    .o(\u_DTCM_CTRL/bram_wea [0]));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    _al_u379 (
    .a(i_ribp_gnt),
    .b(arb1_req0),
    .c(arb1_req1),
    .o(rib_gnt1));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u380 (
    .a(arb1_req0),
    .b(rib_mask1[3]),
    .c(rib_wrcs1),
    .o(\u_ITCM_CTRL/bram_wea [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u381 (
    .a(arb1_req0),
    .b(rib_mask1[2]),
    .c(rib_wrcs1),
    .o(\u_ITCM_CTRL/bram_wea [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u382 (
    .a(arb1_req0),
    .b(rib_mask1[1]),
    .c(rib_wrcs1),
    .o(\u_ITCM_CTRL/bram_wea [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u383 (
    .a(arb1_req0),
    .b(rib_mask1[0]),
    .c(rib_wrcs1),
    .o(\u_ITCM_CTRL/bram_wea [0]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(B*A*~(D*C)))"),
    .INIT(32'hf7770000))
    _al_u384 (
    .a(_al_u319_o),
    .b(_al_u320_o),
    .c(rib_addr1[25]),
    .d(rib_addr1[24]),
    .e(rib_req1),
    .o(o_ribp_req));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    arb2_addr0_pipe (
    .clk(i_clk),
    .d(arb2_addr0[15]),
    .q(arb2_addr0_piped));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    rib_addr1_pipe_b0 (
    .clk(i_clk),
    .d(rib_addr1[14]),
    .q(rib_addr1_piped[0]));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    rib_addr1_pipe_b1 (
    .clk(i_clk),
    .d(rib_addr1[15]),
    .q(rib_addr1_piped[1]));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DTCM_CTRL/handshake_rdy_reg  (
    .clk(i_clk),
    .d(arb1_req1),
    .sr(i_rstn),
    .q(arb1_rsp1));  // ../RTL/periph/bram2rib.v(37)
  // address_offset=0;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x0044"),
    //.WID("0x0044"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_000000_000  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_Nrib_addr1[14]_N_o ),
    .dia({open_n13,open_n14,open_n15,open_n16,open_n17,open_n18,open_n19,open_n20,rib_wdata1[7:0]}),
    .wea(\u_DTCM_CTRL/bram_wea [0]),
    .doa({open_n42,open_n43,open_n44,open_n45,open_n46,open_n47,open_n48,open_n49,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_007 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_006 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_005 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_004 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_003 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_002 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_001 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_000 }));
  // address_offset=0;data_offset=8;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x0048"),
    //.WID("0x0048"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_000000_008  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_Nrib_addr1[14]_N_o ),
    .dia({open_n70,open_n71,open_n72,open_n73,open_n74,open_n75,open_n76,open_n77,rib_wdata1[15:8]}),
    .wea(\u_DTCM_CTRL/bram_wea [1]),
    .doa({open_n99,open_n100,open_n101,open_n102,open_n103,open_n104,open_n105,open_n106,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_015 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_014 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_013 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_012 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_011 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_010 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_009 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_008 }));
  // address_offset=0;data_offset=16;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x004C"),
    //.WID("0x004C"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_000000_016  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_Nrib_addr1[14]_N_o ),
    .dia({open_n127,open_n128,open_n129,open_n130,open_n131,open_n132,open_n133,open_n134,rib_wdata1[23:16]}),
    .wea(\u_DTCM_CTRL/bram_wea [2]),
    .doa({open_n156,open_n157,open_n158,open_n159,open_n160,open_n161,open_n162,open_n163,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_023 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_022 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_021 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_020 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_019 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_018 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_017 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_016 }));
  // address_offset=0;data_offset=24;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x0050"),
    //.WID("0x0050"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_000000_024  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_Nrib_addr1[14]_N_o ),
    .dia({open_n184,open_n185,open_n186,open_n187,open_n188,open_n189,open_n190,open_n191,rib_wdata1[31:24]}),
    .wea(\u_DTCM_CTRL/bram_wea [3]),
    .doa({open_n213,open_n214,open_n215,open_n216,open_n217,open_n218,open_n219,open_n220,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_031 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_030 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_029 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_028 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_027 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_026 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_025 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i0_024 }));
  // address_offset=4096;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x0054"),
    //.WID("0x0054"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_004096_000  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_rib_addr1[14]_Nr_o ),
    .dia({open_n241,open_n242,open_n243,open_n244,open_n245,open_n246,open_n247,open_n248,rib_wdata1[7:0]}),
    .wea(\u_DTCM_CTRL/bram_wea [0]),
    .doa({open_n270,open_n271,open_n272,open_n273,open_n274,open_n275,open_n276,open_n277,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_007 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_006 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_005 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_004 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_003 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_002 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_001 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_000 }));
  // address_offset=4096;data_offset=8;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x0058"),
    //.WID("0x0058"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_004096_008  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_rib_addr1[14]_Nr_o ),
    .dia({open_n298,open_n299,open_n300,open_n301,open_n302,open_n303,open_n304,open_n305,rib_wdata1[15:8]}),
    .wea(\u_DTCM_CTRL/bram_wea [1]),
    .doa({open_n327,open_n328,open_n329,open_n330,open_n331,open_n332,open_n333,open_n334,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_015 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_014 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_013 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_012 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_011 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_010 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_009 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_008 }));
  // address_offset=4096;data_offset=16;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x005C"),
    //.WID("0x005C"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_004096_016  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_rib_addr1[14]_Nr_o ),
    .dia({open_n355,open_n356,open_n357,open_n358,open_n359,open_n360,open_n361,open_n362,rib_wdata1[23:16]}),
    .wea(\u_DTCM_CTRL/bram_wea [2]),
    .doa({open_n384,open_n385,open_n386,open_n387,open_n388,open_n389,open_n390,open_n391,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_023 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_022 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_021 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_020 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_019 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_018 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_017 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_016 }));
  // address_offset=4096;data_offset=24;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x0060"),
    //.WID("0x0060"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_004096_024  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_rib_addr1[14]_Nr_o ),
    .dia({open_n412,open_n413,open_n414,open_n415,open_n416,open_n417,open_n418,open_n419,rib_wdata1[31:24]}),
    .wea(\u_DTCM_CTRL/bram_wea [3]),
    .doa({open_n441,open_n442,open_n443,open_n444,open_n445,open_n446,open_n447,open_n448,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_031 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_030 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_029 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_028 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_027 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_026 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_025 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i1_024 }));
  // address_offset=8192;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x0064"),
    //.WID("0x0064"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_008192_000  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_Nrib_addr1[14]_r_o ),
    .dia({open_n469,open_n470,open_n471,open_n472,open_n473,open_n474,open_n475,open_n476,rib_wdata1[7:0]}),
    .wea(\u_DTCM_CTRL/bram_wea [0]),
    .doa({open_n498,open_n499,open_n500,open_n501,open_n502,open_n503,open_n504,open_n505,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_007 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_006 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_005 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_004 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_003 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_002 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_001 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_000 }));
  // address_offset=8192;data_offset=8;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x0068"),
    //.WID("0x0068"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_008192_008  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_Nrib_addr1[14]_r_o ),
    .dia({open_n526,open_n527,open_n528,open_n529,open_n530,open_n531,open_n532,open_n533,rib_wdata1[15:8]}),
    .wea(\u_DTCM_CTRL/bram_wea [1]),
    .doa({open_n555,open_n556,open_n557,open_n558,open_n559,open_n560,open_n561,open_n562,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_015 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_014 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_013 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_012 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_011 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_010 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_009 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_008 }));
  // address_offset=8192;data_offset=16;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x006C"),
    //.WID("0x006C"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_008192_016  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_Nrib_addr1[14]_r_o ),
    .dia({open_n583,open_n584,open_n585,open_n586,open_n587,open_n588,open_n589,open_n590,rib_wdata1[23:16]}),
    .wea(\u_DTCM_CTRL/bram_wea [2]),
    .doa({open_n612,open_n613,open_n614,open_n615,open_n616,open_n617,open_n618,open_n619,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_023 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_022 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_021 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_020 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_019 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_018 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_017 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_016 }));
  // address_offset=8192;data_offset=24;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x0070"),
    //.WID("0x0070"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_008192_024  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_Nrib_addr1[14]_r_o ),
    .dia({open_n640,open_n641,open_n642,open_n643,open_n644,open_n645,open_n646,open_n647,rib_wdata1[31:24]}),
    .wea(\u_DTCM_CTRL/bram_wea [3]),
    .doa({open_n669,open_n670,open_n671,open_n672,open_n673,open_n674,open_n675,open_n676,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_031 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_030 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_029 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_028 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_027 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_026 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_025 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i2_024 }));
  // address_offset=12288;data_offset=0;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x0074"),
    //.WID("0x0074"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_012288_000  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_rib_addr1[14]_ri_o ),
    .dia({open_n697,open_n698,open_n699,open_n700,open_n701,open_n702,open_n703,open_n704,rib_wdata1[7:0]}),
    .wea(\u_DTCM_CTRL/bram_wea [0]),
    .doa({open_n726,open_n727,open_n728,open_n729,open_n730,open_n731,open_n732,open_n733,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_007 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_006 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_005 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_004 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_003 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_002 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_001 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_000 }));
  // address_offset=12288;data_offset=8;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x0078"),
    //.WID("0x0078"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_012288_008  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_rib_addr1[14]_ri_o ),
    .dia({open_n754,open_n755,open_n756,open_n757,open_n758,open_n759,open_n760,open_n761,rib_wdata1[15:8]}),
    .wea(\u_DTCM_CTRL/bram_wea [1]),
    .doa({open_n783,open_n784,open_n785,open_n786,open_n787,open_n788,open_n789,open_n790,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_015 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_014 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_013 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_012 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_011 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_010 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_009 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_008 }));
  // address_offset=12288;data_offset=16;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x007C"),
    //.WID("0x007C"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_012288_016  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_rib_addr1[14]_ri_o ),
    .dia({open_n811,open_n812,open_n813,open_n814,open_n815,open_n816,open_n817,open_n818,rib_wdata1[23:16]}),
    .wea(\u_DTCM_CTRL/bram_wea [2]),
    .doa({open_n840,open_n841,open_n842,open_n843,open_n844,open_n845,open_n846,open_n847,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_023 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_022 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_021 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_020 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_019 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_018 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_017 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_016 }));
  // address_offset=12288;data_offset=24;depth=4096;width=8;num_section=1;width_per_section=8;section_size=32;working_depth=4096;working_width=8;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM32K #(
    //.RID("0x0080"),
    //.WID("0x0080"),
    .CLKBMUX("0"),
    .CSBMUX("0"),
    .DATA_WIDTH_A("8"),
    .DATA_WIDTH_B("8"),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP16K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .SRMODE("SYNC"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_DTCM_CTRL/u_BRAM_DTCM/inst_16384x32_sub_012288_024  (
    .addra(rib_addr1[13:3]),
    .addrb(11'b00000000000),
    .bytea(rib_addr1[2]),
    .byteb(1'b0),
    .clka(i_clk),
    .csa(\and_rib_addr1[14]_ri_o ),
    .dia({open_n868,open_n869,open_n870,open_n871,open_n872,open_n873,open_n874,open_n875,rib_wdata1[31:24]}),
    .wea(\u_DTCM_CTRL/bram_wea [3]),
    .doa({open_n897,open_n898,open_n899,open_n900,open_n901,open_n902,open_n903,open_n904,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_031 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_030 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_029 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_028 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_027 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_026 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_025 ,\u_DTCM_CTRL/u_BRAM_DTCM/inst_doa_i3_024 }));
  // address_offset=0;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0004"),
    //.WID("0x0004"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000000000FFFFFFFFFFF),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_000  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n937,open_n938,arb2_addr0[15]}),
    .dia({open_n942,open_n943,open_n944,open_n945,open_n946,open_n947,open_n948,arb2_wdata0[0],open_n949}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n964,open_n965,open_n966,open_n967,open_n968,open_n969,open_n970,open_n971,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_000 }));
  // address_offset=0;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0005"),
    //.WID("0x0005"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000000000FFFFFFFFFFF),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_001  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n997,open_n998,arb2_addr0[15]}),
    .dia({open_n1002,open_n1003,open_n1004,open_n1005,open_n1006,open_n1007,open_n1008,arb2_wdata0[1],open_n1009}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n1024,open_n1025,open_n1026,open_n1027,open_n1028,open_n1029,open_n1030,open_n1031,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_001 }));
  // address_offset=0;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0006"),
    //.WID("0x0006"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000000000000000000000000000000000000000000000008782C0A0155),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_002  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1057,open_n1058,arb2_addr0[15]}),
    .dia({open_n1062,open_n1063,open_n1064,open_n1065,open_n1066,open_n1067,open_n1068,arb2_wdata0[2],open_n1069}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n1084,open_n1085,open_n1086,open_n1087,open_n1088,open_n1089,open_n1090,open_n1091,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_002 }));
  // address_offset=0;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0007"),
    //.WID("0x0007"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000002020000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_003  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1117,open_n1118,arb2_addr0[15]}),
    .dia({open_n1122,open_n1123,open_n1124,open_n1125,open_n1126,open_n1127,open_n1128,arb2_wdata0[3],open_n1129}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n1144,open_n1145,open_n1146,open_n1147,open_n1148,open_n1149,open_n1150,open_n1151,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_003 }));
  // address_offset=0;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0008"),
    //.WID("0x0008"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000014E569EC3FF),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_004  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1177,open_n1178,arb2_addr0[15]}),
    .dia({open_n1182,open_n1183,open_n1184,open_n1185,open_n1186,open_n1187,open_n1188,arb2_wdata0[4],open_n1189}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n1204,open_n1205,open_n1206,open_n1207,open_n1208,open_n1209,open_n1210,open_n1211,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_004 }));
  // address_offset=0;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0009"),
    //.WID("0x0009"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000000000E71A9611400),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_005  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1237,open_n1238,arb2_addr0[15]}),
    .dia({open_n1242,open_n1243,open_n1244,open_n1245,open_n1246,open_n1247,open_n1248,arb2_wdata0[5],open_n1249}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n1264,open_n1265,open_n1266,open_n1267,open_n1268,open_n1269,open_n1270,open_n1271,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_005 }));
  // address_offset=0;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000A"),
    //.WID("0x000A"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000000000A3029210400),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_006  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1297,open_n1298,arb2_addr0[15]}),
    .dia({open_n1302,open_n1303,open_n1304,open_n1305,open_n1306,open_n1307,open_n1308,arb2_wdata0[6],open_n1309}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n1324,open_n1325,open_n1326,open_n1327,open_n1328,open_n1329,open_n1330,open_n1331,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_006 }));
  // address_offset=0;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000B"),
    //.WID("0x000B"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000000000000000000000000000000000000000000000003981F1988C3),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_007  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1357,open_n1358,arb2_addr0[15]}),
    .dia({open_n1362,open_n1363,open_n1364,open_n1365,open_n1366,open_n1367,open_n1368,arb2_wdata0[7],open_n1369}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n1384,open_n1385,open_n1386,open_n1387,open_n1388,open_n1389,open_n1390,open_n1391,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_007 }));
  // address_offset=0;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000C"),
    //.WID("0x000C"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000000000000000000000000000000000000000000000001C4529EE0FF),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_008  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1417,open_n1418,arb2_addr0[15]}),
    .dia({open_n1422,open_n1423,open_n1424,open_n1425,open_n1426,open_n1427,open_n1428,arb2_wdata0[8],open_n1429}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n1444,open_n1445,open_n1446,open_n1447,open_n1448,open_n1449,open_n1450,open_n1451,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_008 }));
  // address_offset=0;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000D"),
    //.WID("0x000D"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000000000000000000000000000000000000000000000005C092012F00),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_009  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1477,open_n1478,arb2_addr0[15]}),
    .dia({open_n1482,open_n1483,open_n1484,open_n1485,open_n1486,open_n1487,open_n1488,arb2_wdata0[9],open_n1489}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n1504,open_n1505,open_n1506,open_n1507,open_n1508,open_n1509,open_n1510,open_n1511,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_009 }));
  // address_offset=0;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000E"),
    //.WID("0x000E"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000000000000000000000000000000000000000000000003C7939FC7F0),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_010  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1537,open_n1538,arb2_addr0[15]}),
    .dia({open_n1542,open_n1543,open_n1544,open_n1545,open_n1546,open_n1547,open_n1548,arb2_wdata0[10],open_n1549}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n1564,open_n1565,open_n1566,open_n1567,open_n1568,open_n1569,open_n1570,open_n1571,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_010 }));
  // address_offset=0;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x000F"),
    //.WID("0x000F"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000020013200400),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_011  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1597,open_n1598,arb2_addr0[15]}),
    .dia({open_n1602,open_n1603,open_n1604,open_n1605,open_n1606,open_n1607,open_n1608,arb2_wdata0[11],open_n1609}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n1624,open_n1625,open_n1626,open_n1627,open_n1628,open_n1629,open_n1630,open_n1631,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_011 }));
  // address_offset=0;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0010"),
    //.WID("0x0010"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000010000200401),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_012  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1657,open_n1658,arb2_addr0[15]}),
    .dia({open_n1662,open_n1663,open_n1664,open_n1665,open_n1666,open_n1667,open_n1668,arb2_wdata0[12],open_n1669}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n1684,open_n1685,open_n1686,open_n1687,open_n1688,open_n1689,open_n1690,open_n1691,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_012 }));
  // address_offset=0;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0011"),
    //.WID("0x0011"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000058181613C00),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_013  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1717,open_n1718,arb2_addr0[15]}),
    .dia({open_n1722,open_n1723,open_n1724,open_n1725,open_n1726,open_n1727,open_n1728,arb2_wdata0[13],open_n1729}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n1744,open_n1745,open_n1746,open_n1747,open_n1748,open_n1749,open_n1750,open_n1751,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_013 }));
  // address_offset=0;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0012"),
    //.WID("0x0012"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000010001210400),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_014  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1777,open_n1778,arb2_addr0[15]}),
    .dia({open_n1782,open_n1783,open_n1784,open_n1785,open_n1786,open_n1787,open_n1788,arb2_wdata0[14],open_n1789}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n1804,open_n1805,open_n1806,open_n1807,open_n1808,open_n1809,open_n1810,open_n1811,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_014 }));
  // address_offset=0;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0013"),
    //.WID("0x0013"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000000000B100811B482),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_015  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1837,open_n1838,arb2_addr0[15]}),
    .dia({open_n1842,open_n1843,open_n1844,open_n1845,open_n1846,open_n1847,open_n1848,arb2_wdata0[15],open_n1849}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n1864,open_n1865,open_n1866,open_n1867,open_n1868,open_n1869,open_n1870,open_n1871,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_015 }));
  // address_offset=0;data_offset=16;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0014"),
    //.WID("0x0014"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000000000783C1F5FCAE),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_016  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1897,open_n1898,arb2_addr0[15]}),
    .dia({open_n1902,open_n1903,open_n1904,open_n1905,open_n1906,open_n1907,open_n1908,arb2_wdata0[16],open_n1909}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n1924,open_n1925,open_n1926,open_n1927,open_n1928,open_n1929,open_n1930,open_n1931,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_016 }));
  // address_offset=0;data_offset=17;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0015"),
    //.WID("0x0015"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000078000000200),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_017  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n1957,open_n1958,arb2_addr0[15]}),
    .dia({open_n1962,open_n1963,open_n1964,open_n1965,open_n1966,open_n1967,open_n1968,arb2_wdata0[17],open_n1969}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n1984,open_n1985,open_n1986,open_n1987,open_n1988,open_n1989,open_n1990,open_n1991,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_017 }));
  // address_offset=0;data_offset=18;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0016"),
    //.WID("0x0016"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000078001F5FEA0),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_018  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2017,open_n2018,arb2_addr0[15]}),
    .dia({open_n2022,open_n2023,open_n2024,open_n2025,open_n2026,open_n2027,open_n2028,arb2_wdata0[18],open_n2029}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n2044,open_n2045,open_n2046,open_n2047,open_n2048,open_n2049,open_n2050,open_n2051,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_018 }));
  // address_offset=0;data_offset=19;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0017"),
    //.WID("0x0017"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_019  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2077,open_n2078,arb2_addr0[15]}),
    .dia({open_n2082,open_n2083,open_n2084,open_n2085,open_n2086,open_n2087,open_n2088,arb2_wdata0[19],open_n2089}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n2104,open_n2105,open_n2106,open_n2107,open_n2108,open_n2109,open_n2110,open_n2111,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_019 }));
  // address_offset=0;data_offset=20;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0018"),
    //.WID("0x0018"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000010481201000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_020  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2137,open_n2138,arb2_addr0[15]}),
    .dia({open_n2142,open_n2143,open_n2144,open_n2145,open_n2146,open_n2147,open_n2148,arb2_wdata0[20],open_n2149}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n2164,open_n2165,open_n2166,open_n2167,open_n2168,open_n2169,open_n2170,open_n2171,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_020 }));
  // address_offset=0;data_offset=21;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0019"),
    //.WID("0x0019"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000040011200000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_021  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2197,open_n2198,arb2_addr0[15]}),
    .dia({open_n2202,open_n2203,open_n2204,open_n2205,open_n2206,open_n2207,open_n2208,arb2_wdata0[21],open_n2209}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n2224,open_n2225,open_n2226,open_n2227,open_n2228,open_n2229,open_n2230,open_n2231,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_021 }));
  // address_offset=0;data_offset=22;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x001A"),
    //.WID("0x001A"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000000000000000000000000000000000000000000000000100095D400),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_022  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2257,open_n2258,arb2_addr0[15]}),
    .dia({open_n2262,open_n2263,open_n2264,open_n2265,open_n2266,open_n2267,open_n2268,arb2_wdata0[22],open_n2269}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n2284,open_n2285,open_n2286,open_n2287,open_n2288,open_n2289,open_n2290,open_n2291,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_022 }));
  // address_offset=0;data_offset=23;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x001B"),
    //.WID("0x001B"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000041111250488),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_023  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2317,open_n2318,arb2_addr0[15]}),
    .dia({open_n2322,open_n2323,open_n2324,open_n2325,open_n2326,open_n2327,open_n2328,arb2_wdata0[23],open_n2329}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n2344,open_n2345,open_n2346,open_n2347,open_n2348,open_n2349,open_n2350,open_n2351,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_023 }));
  // address_offset=0;data_offset=24;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x001C"),
    //.WID("0x001C"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000000000042481E014D),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_024  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2377,open_n2378,arb2_addr0[15]}),
    .dia({open_n2382,open_n2383,open_n2384,open_n2385,open_n2386,open_n2387,open_n2388,arb2_wdata0[24],open_n2389}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n2404,open_n2405,open_n2406,open_n2407,open_n2408,open_n2409,open_n2410,open_n2411,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_024 }));
  // address_offset=0;data_offset=25;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x001D"),
    //.WID("0x001D"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000000000204531502A8),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_025  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2437,open_n2438,arb2_addr0[15]}),
    .dia({open_n2442,open_n2443,open_n2444,open_n2445,open_n2446,open_n2447,open_n2448,arb2_wdata0[25],open_n2449}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n2464,open_n2465,open_n2466,open_n2467,open_n2468,open_n2469,open_n2470,open_n2471,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_025 }));
  // address_offset=0;data_offset=26;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x001E"),
    //.WID("0x001E"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000020441010288),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_026  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2497,open_n2498,arb2_addr0[15]}),
    .dia({open_n2502,open_n2503,open_n2504,open_n2505,open_n2506,open_n2507,open_n2508,arb2_wdata0[26],open_n2509}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n2524,open_n2525,open_n2526,open_n2527,open_n2528,open_n2529,open_n2530,open_n2531,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_026 }));
  // address_offset=0;data_offset=27;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x001F"),
    //.WID("0x001F"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00000000000000000000000000000000000000000000000000000200531502A8),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_027  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2557,open_n2558,arb2_addr0[15]}),
    .dia({open_n2562,open_n2563,open_n2564,open_n2565,open_n2566,open_n2567,open_n2568,arb2_wdata0[27],open_n2569}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n2584,open_n2585,open_n2586,open_n2587,open_n2588,open_n2589,open_n2590,open_n2591,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_027 }));
  // address_offset=0;data_offset=28;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0020"),
    //.WID("0x0020"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000024041150288),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_028  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2617,open_n2618,arb2_addr0[15]}),
    .dia({open_n2622,open_n2623,open_n2624,open_n2625,open_n2626,open_n2627,open_n2628,arb2_wdata0[28],open_n2629}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n2644,open_n2645,open_n2646,open_n2647,open_n2648,open_n2649,open_n2650,open_n2651,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_028 }));
  // address_offset=0;data_offset=29;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0021"),
    //.WID("0x0021"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000024041150288),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_029  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2677,open_n2678,arb2_addr0[15]}),
    .dia({open_n2682,open_n2683,open_n2684,open_n2685,open_n2686,open_n2687,open_n2688,arb2_wdata0[29],open_n2689}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n2704,open_n2705,open_n2706,open_n2707,open_n2708,open_n2709,open_n2710,open_n2711,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_029 }));
  // address_offset=0;data_offset=30;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0022"),
    //.WID("0x0022"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000024041150288),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_030  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2737,open_n2738,arb2_addr0[15]}),
    .dia({open_n2742,open_n2743,open_n2744,open_n2745,open_n2746,open_n2747,open_n2748,arb2_wdata0[30],open_n2749}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n2764,open_n2765,open_n2766,open_n2767,open_n2768,open_n2769,open_n2770,open_n2771,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_030 }));
  // address_offset=0;data_offset=31;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0023"),
    //.WID("0x0023"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000000000000000000000000000000000000000000000002404115028A),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_000000_031  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2797,open_n2798,arb2_addr0[15]}),
    .dia({open_n2802,open_n2803,open_n2804,open_n2805,open_n2806,open_n2807,open_n2808,arb2_wdata0[31],open_n2809}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n2824,open_n2825,open_n2826,open_n2827,open_n2828,open_n2829,open_n2830,open_n2831,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i0_031 }));
  // address_offset=8192;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0024"),
    //.WID("0x0024"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_000  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2857,open_n2858,arb2_addr0[15]}),
    .dia({open_n2862,open_n2863,open_n2864,open_n2865,open_n2866,open_n2867,open_n2868,arb2_wdata0[0],open_n2869}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n2884,open_n2885,open_n2886,open_n2887,open_n2888,open_n2889,open_n2890,open_n2891,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_000 }));
  // address_offset=8192;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0025"),
    //.WID("0x0025"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_001  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2917,open_n2918,arb2_addr0[15]}),
    .dia({open_n2922,open_n2923,open_n2924,open_n2925,open_n2926,open_n2927,open_n2928,arb2_wdata0[1],open_n2929}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n2944,open_n2945,open_n2946,open_n2947,open_n2948,open_n2949,open_n2950,open_n2951,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_001 }));
  // address_offset=8192;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0026"),
    //.WID("0x0026"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_002  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n2977,open_n2978,arb2_addr0[15]}),
    .dia({open_n2982,open_n2983,open_n2984,open_n2985,open_n2986,open_n2987,open_n2988,arb2_wdata0[2],open_n2989}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n3004,open_n3005,open_n3006,open_n3007,open_n3008,open_n3009,open_n3010,open_n3011,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_002 }));
  // address_offset=8192;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0027"),
    //.WID("0x0027"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_003  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3037,open_n3038,arb2_addr0[15]}),
    .dia({open_n3042,open_n3043,open_n3044,open_n3045,open_n3046,open_n3047,open_n3048,arb2_wdata0[3],open_n3049}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n3064,open_n3065,open_n3066,open_n3067,open_n3068,open_n3069,open_n3070,open_n3071,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_003 }));
  // address_offset=8192;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0028"),
    //.WID("0x0028"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_004  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3097,open_n3098,arb2_addr0[15]}),
    .dia({open_n3102,open_n3103,open_n3104,open_n3105,open_n3106,open_n3107,open_n3108,arb2_wdata0[4],open_n3109}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n3124,open_n3125,open_n3126,open_n3127,open_n3128,open_n3129,open_n3130,open_n3131,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_004 }));
  // address_offset=8192;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0029"),
    //.WID("0x0029"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_005  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3157,open_n3158,arb2_addr0[15]}),
    .dia({open_n3162,open_n3163,open_n3164,open_n3165,open_n3166,open_n3167,open_n3168,arb2_wdata0[5],open_n3169}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n3184,open_n3185,open_n3186,open_n3187,open_n3188,open_n3189,open_n3190,open_n3191,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_005 }));
  // address_offset=8192;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x002A"),
    //.WID("0x002A"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_006  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3217,open_n3218,arb2_addr0[15]}),
    .dia({open_n3222,open_n3223,open_n3224,open_n3225,open_n3226,open_n3227,open_n3228,arb2_wdata0[6],open_n3229}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n3244,open_n3245,open_n3246,open_n3247,open_n3248,open_n3249,open_n3250,open_n3251,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_006 }));
  // address_offset=8192;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x002B"),
    //.WID("0x002B"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_007  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3277,open_n3278,arb2_addr0[15]}),
    .dia({open_n3282,open_n3283,open_n3284,open_n3285,open_n3286,open_n3287,open_n3288,arb2_wdata0[7],open_n3289}),
    .wea(\u_ITCM_CTRL/bram_wea [0]),
    .doa({open_n3304,open_n3305,open_n3306,open_n3307,open_n3308,open_n3309,open_n3310,open_n3311,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_007 }));
  // address_offset=8192;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x002C"),
    //.WID("0x002C"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_008  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3337,open_n3338,arb2_addr0[15]}),
    .dia({open_n3342,open_n3343,open_n3344,open_n3345,open_n3346,open_n3347,open_n3348,arb2_wdata0[8],open_n3349}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n3364,open_n3365,open_n3366,open_n3367,open_n3368,open_n3369,open_n3370,open_n3371,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_008 }));
  // address_offset=8192;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x002D"),
    //.WID("0x002D"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_009  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3397,open_n3398,arb2_addr0[15]}),
    .dia({open_n3402,open_n3403,open_n3404,open_n3405,open_n3406,open_n3407,open_n3408,arb2_wdata0[9],open_n3409}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n3424,open_n3425,open_n3426,open_n3427,open_n3428,open_n3429,open_n3430,open_n3431,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_009 }));
  // address_offset=8192;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x002E"),
    //.WID("0x002E"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_010  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3457,open_n3458,arb2_addr0[15]}),
    .dia({open_n3462,open_n3463,open_n3464,open_n3465,open_n3466,open_n3467,open_n3468,arb2_wdata0[10],open_n3469}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n3484,open_n3485,open_n3486,open_n3487,open_n3488,open_n3489,open_n3490,open_n3491,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_010 }));
  // address_offset=8192;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x002F"),
    //.WID("0x002F"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_011  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3517,open_n3518,arb2_addr0[15]}),
    .dia({open_n3522,open_n3523,open_n3524,open_n3525,open_n3526,open_n3527,open_n3528,arb2_wdata0[11],open_n3529}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n3544,open_n3545,open_n3546,open_n3547,open_n3548,open_n3549,open_n3550,open_n3551,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_011 }));
  // address_offset=8192;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0030"),
    //.WID("0x0030"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_012  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3577,open_n3578,arb2_addr0[15]}),
    .dia({open_n3582,open_n3583,open_n3584,open_n3585,open_n3586,open_n3587,open_n3588,arb2_wdata0[12],open_n3589}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n3604,open_n3605,open_n3606,open_n3607,open_n3608,open_n3609,open_n3610,open_n3611,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_012 }));
  // address_offset=8192;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0031"),
    //.WID("0x0031"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_013  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3637,open_n3638,arb2_addr0[15]}),
    .dia({open_n3642,open_n3643,open_n3644,open_n3645,open_n3646,open_n3647,open_n3648,arb2_wdata0[13],open_n3649}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n3664,open_n3665,open_n3666,open_n3667,open_n3668,open_n3669,open_n3670,open_n3671,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_013 }));
  // address_offset=8192;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0032"),
    //.WID("0x0032"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_014  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3697,open_n3698,arb2_addr0[15]}),
    .dia({open_n3702,open_n3703,open_n3704,open_n3705,open_n3706,open_n3707,open_n3708,arb2_wdata0[14],open_n3709}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n3724,open_n3725,open_n3726,open_n3727,open_n3728,open_n3729,open_n3730,open_n3731,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_014 }));
  // address_offset=8192;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0033"),
    //.WID("0x0033"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_015  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3757,open_n3758,arb2_addr0[15]}),
    .dia({open_n3762,open_n3763,open_n3764,open_n3765,open_n3766,open_n3767,open_n3768,arb2_wdata0[15],open_n3769}),
    .wea(\u_ITCM_CTRL/bram_wea [1]),
    .doa({open_n3784,open_n3785,open_n3786,open_n3787,open_n3788,open_n3789,open_n3790,open_n3791,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_015 }));
  // address_offset=8192;data_offset=16;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0034"),
    //.WID("0x0034"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_016  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3817,open_n3818,arb2_addr0[15]}),
    .dia({open_n3822,open_n3823,open_n3824,open_n3825,open_n3826,open_n3827,open_n3828,arb2_wdata0[16],open_n3829}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n3844,open_n3845,open_n3846,open_n3847,open_n3848,open_n3849,open_n3850,open_n3851,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_016 }));
  // address_offset=8192;data_offset=17;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0035"),
    //.WID("0x0035"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_017  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3877,open_n3878,arb2_addr0[15]}),
    .dia({open_n3882,open_n3883,open_n3884,open_n3885,open_n3886,open_n3887,open_n3888,arb2_wdata0[17],open_n3889}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n3904,open_n3905,open_n3906,open_n3907,open_n3908,open_n3909,open_n3910,open_n3911,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_017 }));
  // address_offset=8192;data_offset=18;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0036"),
    //.WID("0x0036"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_018  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3937,open_n3938,arb2_addr0[15]}),
    .dia({open_n3942,open_n3943,open_n3944,open_n3945,open_n3946,open_n3947,open_n3948,arb2_wdata0[18],open_n3949}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n3964,open_n3965,open_n3966,open_n3967,open_n3968,open_n3969,open_n3970,open_n3971,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_018 }));
  // address_offset=8192;data_offset=19;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0037"),
    //.WID("0x0037"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_019  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n3997,open_n3998,arb2_addr0[15]}),
    .dia({open_n4002,open_n4003,open_n4004,open_n4005,open_n4006,open_n4007,open_n4008,arb2_wdata0[19],open_n4009}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n4024,open_n4025,open_n4026,open_n4027,open_n4028,open_n4029,open_n4030,open_n4031,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_019 }));
  // address_offset=8192;data_offset=20;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0038"),
    //.WID("0x0038"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_020  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n4057,open_n4058,arb2_addr0[15]}),
    .dia({open_n4062,open_n4063,open_n4064,open_n4065,open_n4066,open_n4067,open_n4068,arb2_wdata0[20],open_n4069}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n4084,open_n4085,open_n4086,open_n4087,open_n4088,open_n4089,open_n4090,open_n4091,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_020 }));
  // address_offset=8192;data_offset=21;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0039"),
    //.WID("0x0039"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_021  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n4117,open_n4118,arb2_addr0[15]}),
    .dia({open_n4122,open_n4123,open_n4124,open_n4125,open_n4126,open_n4127,open_n4128,arb2_wdata0[21],open_n4129}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n4144,open_n4145,open_n4146,open_n4147,open_n4148,open_n4149,open_n4150,open_n4151,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_021 }));
  // address_offset=8192;data_offset=22;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x003A"),
    //.WID("0x003A"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_022  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n4177,open_n4178,arb2_addr0[15]}),
    .dia({open_n4182,open_n4183,open_n4184,open_n4185,open_n4186,open_n4187,open_n4188,arb2_wdata0[22],open_n4189}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n4204,open_n4205,open_n4206,open_n4207,open_n4208,open_n4209,open_n4210,open_n4211,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_022 }));
  // address_offset=8192;data_offset=23;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x003B"),
    //.WID("0x003B"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_023  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n4237,open_n4238,arb2_addr0[15]}),
    .dia({open_n4242,open_n4243,open_n4244,open_n4245,open_n4246,open_n4247,open_n4248,arb2_wdata0[23],open_n4249}),
    .wea(\u_ITCM_CTRL/bram_wea [2]),
    .doa({open_n4264,open_n4265,open_n4266,open_n4267,open_n4268,open_n4269,open_n4270,open_n4271,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_023 }));
  // address_offset=8192;data_offset=24;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x003C"),
    //.WID("0x003C"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_024  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n4297,open_n4298,arb2_addr0[15]}),
    .dia({open_n4302,open_n4303,open_n4304,open_n4305,open_n4306,open_n4307,open_n4308,arb2_wdata0[24],open_n4309}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n4324,open_n4325,open_n4326,open_n4327,open_n4328,open_n4329,open_n4330,open_n4331,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_024 }));
  // address_offset=8192;data_offset=25;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x003D"),
    //.WID("0x003D"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_025  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n4357,open_n4358,arb2_addr0[15]}),
    .dia({open_n4362,open_n4363,open_n4364,open_n4365,open_n4366,open_n4367,open_n4368,arb2_wdata0[25],open_n4369}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n4384,open_n4385,open_n4386,open_n4387,open_n4388,open_n4389,open_n4390,open_n4391,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_025 }));
  // address_offset=8192;data_offset=26;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x003E"),
    //.WID("0x003E"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_026  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n4417,open_n4418,arb2_addr0[15]}),
    .dia({open_n4422,open_n4423,open_n4424,open_n4425,open_n4426,open_n4427,open_n4428,arb2_wdata0[26],open_n4429}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n4444,open_n4445,open_n4446,open_n4447,open_n4448,open_n4449,open_n4450,open_n4451,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_026 }));
  // address_offset=8192;data_offset=27;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x003F"),
    //.WID("0x003F"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_027  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n4477,open_n4478,arb2_addr0[15]}),
    .dia({open_n4482,open_n4483,open_n4484,open_n4485,open_n4486,open_n4487,open_n4488,arb2_wdata0[27],open_n4489}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n4504,open_n4505,open_n4506,open_n4507,open_n4508,open_n4509,open_n4510,open_n4511,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_027 }));
  // address_offset=8192;data_offset=28;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0040"),
    //.WID("0x0040"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_028  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n4537,open_n4538,arb2_addr0[15]}),
    .dia({open_n4542,open_n4543,open_n4544,open_n4545,open_n4546,open_n4547,open_n4548,arb2_wdata0[28],open_n4549}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n4564,open_n4565,open_n4566,open_n4567,open_n4568,open_n4569,open_n4570,open_n4571,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_028 }));
  // address_offset=8192;data_offset=29;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0041"),
    //.WID("0x0041"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_029  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n4597,open_n4598,arb2_addr0[15]}),
    .dia({open_n4602,open_n4603,open_n4604,open_n4605,open_n4606,open_n4607,open_n4608,arb2_wdata0[29],open_n4609}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n4624,open_n4625,open_n4626,open_n4627,open_n4628,open_n4629,open_n4630,open_n4631,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_029 }));
  // address_offset=8192;data_offset=30;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0042"),
    //.WID("0x0042"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_030  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n4657,open_n4658,arb2_addr0[15]}),
    .dia({open_n4662,open_n4663,open_n4664,open_n4665,open_n4666,open_n4667,open_n4668,arb2_wdata0[30],open_n4669}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n4684,open_n4685,open_n4686,open_n4687,open_n4688,open_n4689,open_n4690,open_n4691,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_030 }));
  // address_offset=8192;data_offset=31;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    //.RID("0x0043"),
    //.WID("0x0043"),
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .READBACK("ON"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    \u_ITCM_CTRL/u_BRAM_ITCM/inst_16384x32_sub_008192_031  (
    .addra(arb2_addr0[14:2]),
    .clka(i_clk),
    .csa({open_n4717,open_n4718,arb2_addr0[15]}),
    .dia({open_n4722,open_n4723,open_n4724,open_n4725,open_n4726,open_n4727,open_n4728,arb2_wdata0[31],open_n4729}),
    .wea(\u_ITCM_CTRL/bram_wea [3]),
    .doa({open_n4744,open_n4745,open_n4746,open_n4747,open_n4748,open_n4749,open_n4750,open_n4751,\u_ITCM_CTRL/u_BRAM_ITCM/inst_doa_i1_031 }));
  RITTER_TOP u_RITTER_TOP (
    .i_clk(i_clk),
    .i_ribm_gnt0(arb0_gnt0),
    .i_ribm_gnt1(rib_gnt1),
    .i_ribm_rdata0(rib_rdata0),
    .i_ribm_rdata1(rib_rdata1),
    .i_ribm_rsp0(arb0_rsp0),
    .i_ribm_rsp1(rib_rsp1),
    .i_rstn(i_rstn),
    .o_ribm_addr0({rib_addr0[31:24],open_n4761,open_n4762,open_n4763,open_n4764,open_n4765,open_n4766,open_n4767,open_n4768,rib_addr0[15:2],open_n4769,open_n4770}),
    .o_ribm_addr1({rib_addr1[31:24],open_n4771,open_n4772,open_n4773,open_n4774,open_n4775,open_n4776,open_n4777,open_n4778,rib_addr1[15:2],open_n4779,open_n4780}),
    .o_ribm_mask1(rib_mask1),
    .o_ribm_req0(rib_req0),
    .o_ribm_req1(rib_req1),
    .o_ribm_wdata1(rib_wdata1),
    .o_ribm_wrcs1(rib_wrcs1));  // ../RTL/soc_top/core_top.v(59)

endmodule 

module RITTER_TOP  // ../RTL/core/ritter_top.v(6)
  (
  i_clk,
  i_ribm_gnt0,
  i_ribm_gnt1,
  i_ribm_rdata0,
  i_ribm_rdata1,
  i_ribm_rsp0,
  i_ribm_rsp1,
  i_rstn,
  o_ribm_addr0,
  o_ribm_addr1,
  o_ribm_mask0,
  o_ribm_mask1,
  o_ribm_rdy0,
  o_ribm_rdy1,
  o_ribm_req0,
  o_ribm_req1,
  o_ribm_wdata0,
  o_ribm_wdata1,
  o_ribm_wrcs0,
  o_ribm_wrcs1
  );

  input i_clk;  // ../RTL/core/ritter_top.v(7)
  input i_ribm_gnt0;  // ../RTL/core/ritter_top.v(17)
  input i_ribm_gnt1;  // ../RTL/core/ritter_top.v(27)
  input [31:0] i_ribm_rdata0;  // ../RTL/core/ritter_top.v(15)
  input [31:0] i_ribm_rdata1;  // ../RTL/core/ritter_top.v(25)
  input i_ribm_rsp0;  // ../RTL/core/ritter_top.v(18)
  input i_ribm_rsp1;  // ../RTL/core/ritter_top.v(28)
  input i_rstn;  // ../RTL/core/ritter_top.v(8)
  output [31:0] o_ribm_addr0;  // ../RTL/core/ritter_top.v(11)
  output [31:0] o_ribm_addr1;  // ../RTL/core/ritter_top.v(21)
  output [3:0] o_ribm_mask0;  // ../RTL/core/ritter_top.v(13)
  output [3:0] o_ribm_mask1;  // ../RTL/core/ritter_top.v(23)
  output o_ribm_rdy0;  // ../RTL/core/ritter_top.v(19)
  output o_ribm_rdy1;  // ../RTL/core/ritter_top.v(29)
  output o_ribm_req0;  // ../RTL/core/ritter_top.v(16)
  output o_ribm_req1;  // ../RTL/core/ritter_top.v(26)
  output [31:0] o_ribm_wdata0;  // ../RTL/core/ritter_top.v(14)
  output [31:0] o_ribm_wdata1;  // ../RTL/core/ritter_top.v(24)
  output o_ribm_wrcs0;  // ../RTL/core/ritter_top.v(12)
  output o_ribm_wrcs1;  // ../RTL/core/ritter_top.v(22)

  wire [31:0] bpu_csr_zimm;  // ../RTL/core/ritter_top.v(153)
  wire [11:0] bpu_csridx;  // ../RTL/core/ritter_top.v(151)
  wire [9:0] bpu_decinfo;  // ../RTL/core/ritter_top.v(155)
  wire [5:0] bpu_decinfo_grp;  // ../RTL/core/ritter_top.v(154)
  wire [31:0] bpu_exu_op1;  // ../RTL/core/ritter_top.v(143)
  wire [31:0] bpu_exu_op2;  // ../RTL/core/ritter_top.v(144)
  wire [31:0] bpu_iaddr;  // ../RTL/core/ritter_top.v(156)
  wire [31:0] bpu_imm;  // ../RTL/core/ritter_top.v(146)
  wire [31:0] bpu_jaddr;  // ../RTL/core/ritter_top.v(141)
  wire [31:0] bpu_jaddr_gen;  // ../RTL/core/ritter_top.v(79)
  wire [4:0] bpu_rdidx;  // ../RTL/core/ritter_top.v(148)
  wire [31:0] bpu_rs2rdata;  // ../RTL/core/ritter_top.v(145)
  wire [31:0] csr_rdata;  // ../RTL/core/ritter_top.v(200)
  wire [4:0] ctrl2bpu_rs1idx;  // ../RTL/core/ritter_top.v(34)
  wire [4:0] ctrl2bpu_rs2idx;  // ../RTL/core/ritter_top.v(36)
  wire [4:0] ctrl2exu_rdidx0;  // ../RTL/core/ritter_top.v(39)
  wire [4:0] ctrl2exu_rdidx1;  // ../RTL/core/ritter_top.v(42)
  wire [4:0] ctrl2exu_rdidx2;  // ../RTL/core/ritter_top.v(44)
  wire [31:0] dis_csr_rdata;  // ../RTL/core/ritter_top.v(230)
  wire [31:0] dis_csr_zimm;  // ../RTL/core/ritter_top.v(231)
  wire [11:0] dis_csridx;  // ../RTL/core/ritter_top.v(229)
  wire [9:0] dis_decinfo;  // ../RTL/core/ritter_top.v(234)
  wire [5:0] dis_decinfo_grp;  // ../RTL/core/ritter_top.v(233)
  wire [31:0] dis_exu_op1;  // ../RTL/core/ritter_top.v(222)
  wire [31:0] dis_exu_op2;  // ../RTL/core/ritter_top.v(223)
  wire [31:0] dis_iaddr;  // ../RTL/core/ritter_top.v(235)
  wire [31:0] dis_imm;  // ../RTL/core/ritter_top.v(225)
  wire [4:0] dis_rdidx;  // ../RTL/core/ritter_top.v(227)
  wire [31:0] dis_rs2rdata;  // ../RTL/core/ritter_top.v(224)
  wire [31:0] exu_jaddr;  // ../RTL/core/ritter_top.v(296)
  wire [31:0] exu_jaddr_gen;  // ../RTL/core/ritter_top.v(81)
  wire [4:0] exu_rdidx0;  // ../RTL/core/ritter_top.v(284)
  wire [4:0] exu_rdidx1;  // ../RTL/core/ritter_top.v(288)
  wire [4:0] exu_rdidx2;  // ../RTL/core/ritter_top.v(292)
  wire [31:0] exu_rdwdata0;  // ../RTL/core/ritter_top.v(285)
  wire [31:0] exu_rdwdata1;  // ../RTL/core/ritter_top.v(289)
  wire [31:0] exu_rdwdata2;  // ../RTL/core/ritter_top.v(293)
  wire [31:0] ifu2bpu_data;  // ../RTL/core/ritter_top.v(117)
  wire [31:0] ifu2bpu_iaddr;  // ../RTL/core/ritter_top.v(116)
  wire [31:0] ifu_iaddr;  // ../RTL/core/ritter_top.v(83)
  wire [5:0] \u_DISPATCH/n5 ;
  wire [31:0] \u_IFU/fetch_addr ;  // ../RTL/core/ifu.v(80)
  wire [0:0] \u_IFU/fifo_cnt ;  // ../RTL/core/ifu.v(130)
  wire [31:0] \u_IFU/jump_addr ;  // ../RTL/core/ifu.v(62)
  wire [31:0] \u_IFU/u_IFU_PC/n10 ;
  wire [29:0] \u_IFU/u_IFU_PC/n2 ;
  wire [29:0] \u_IFU/u_IFU_PC/n4 ;
  wire [31:0] \u_IFU/u_IFU_PC/n9 ;
  wire [31:0] \u_IFU/u_IFU_PC/pc ;  // ../RTL/core/ifu_pc.v(23)
  wire [8:0] \u_IFU2BPU/fifo_cnt ;  // ../RTL/core/ifu2bpu.v(37)
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_di ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_waddr ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/eptr ;  // ../RTL/core/fifos.v(36)
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/hptr ;  // ../RTL/core/fifos.v(36)
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n16 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n22 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n23 ;
  wire [3:0] \u_IFU2BPU/u_SYNC_FIFO/n24 ;
  wire [31:0] \u_PIPE_CTRL/n1 ;
  wire [31:0] \u_PIPE_CTRL/n11 ;
  wire [31:0] \u_PIPE_CTRL/n14 ;
  wire [31:0] \u_PIPE_CTRL/n3 ;
  wire [31:0] \u_PIPE_CTRL/n6 ;
  wire [31:0] \u_PIPE_CTRL/n9 ;
  wire [4:0] \u_WB/rdidx0 ;  // ../RTL/core/wb.v(48)
  wire [4:0] \u_WB/rdidx1 ;  // ../RTL/core/wb.v(49)
  wire [4:0] \u_WB/rdidx2 ;  // ../RTL/core/wb.v(50)
  wire [31:0] \u_WB/rdwdata0 ;  // ../RTL/core/wb.v(51)
  wire [31:0] \u_WB/rdwdata1 ;  // ../RTL/core/wb.v(52)
  wire [31:0] \u_WB/rdwdata2 ;  // ../RTL/core/wb.v(53)
  wire [31:0] wb_csr_wdata;  // ../RTL/core/ritter_top.v(204)
  wire [11:0] wb_csridx;  // ../RTL/core/ritter_top.v(203)
  wire [4:0] wb_rdidx;  // ../RTL/core/ritter_top.v(137)
  wire [31:0] wb_rdwdata;  // ../RTL/core/ritter_top.v(138)
  wire _al_u564_o;
  wire _al_u571_o;
  wire _al_u572_o;
  wire _al_u574_o;
  wire _al_u575_o;
  wire _al_u577_o;
  wire _al_u578_o;
  wire _al_u581_o;
  wire _al_u582_o;
  wire _al_u584_o;
  wire _al_u585_o;
  wire _al_u587_o;
  wire _al_u588_o;
  wire _al_u590_o;
  wire _al_u603_o;
  wire _al_u605_o;
  wire _al_u611_o;
  wire _al_u614_o;
  wire _al_u617_o;
  wire _al_u620_o;
  wire _al_u623_o;
  wire _al_u626_o;
  wire _al_u629_o;
  wire _al_u632_o;
  wire _al_u635_o;
  wire _al_u638_o;
  wire _al_u641_o;
  wire _al_u644_o;
  wire _al_u647_o;
  wire _al_u650_o;
  wire _al_u653_o;
  wire _al_u656_o;
  wire _al_u659_o;
  wire _al_u662_o;
  wire _al_u665_o;
  wire _al_u667_o;
  wire _al_u668_o;
  wire _al_u671_o;
  wire _al_u674_o;
  wire _al_u677_o;
  wire _al_u680_o;
  wire _al_u683_o;
  wire _al_u686_o;
  wire _al_u689_o;
  wire _al_u692_o;
  wire _al_u695_o;
  wire _al_u698_o;
  wire _al_u700_o;
  wire _al_u702_o;
  wire _al_u704_o;
  wire _al_u710_o;
  wire _al_u713_o;
  wire bpu_inst_vld;  // ../RTL/core/ritter_top.v(142)
  wire bpu_rdwen;  // ../RTL/core/ritter_top.v(147)
  wire bpu_taken;  // ../RTL/core/ritter_top.v(140)
  wire bpu_taken_gen;  // ../RTL/core/ritter_top.v(78)
  wire ctrl2bpu_rs1ren;  // ../RTL/core/ritter_top.v(33)
  wire ctrl2bpu_rs2ren;  // ../RTL/core/ritter_top.v(35)
  wire ctrl2bpu_wait;  // ../RTL/core/ritter_top.v(50)
  wire ctrl2exu_rdwen0;  // ../RTL/core/ritter_top.v(38)
  wire ctrl2exu_rdwen1;  // ../RTL/core/ritter_top.v(41)
  wire ctrl2exu_rdwen2;  // ../RTL/core/ritter_top.v(43)
  wire ctrl2exu_resource_match;  // ../RTL/core/ritter_top.v(46)
  wire dis_rdwen;  // ../RTL/core/ritter_top.v(226)
  wire exu_rdwen0;  // ../RTL/core/ritter_top.v(283)
  wire exu_rdwen1;  // ../RTL/core/ritter_top.v(287)
  wire exu_rdwen2;  // ../RTL/core/ritter_top.v(291)
  wire exu_taken;  // ../RTL/core/ritter_top.v(295)
  wire exu_taken_gen;  // ../RTL/core/ritter_top.v(80)
  wire ifu_data_vld;  // ../RTL/core/ritter_top.v(82)
  wire n3_lutinv;
  wire n5;
  wire \u_DISPATCH/mux12_b0_sel_is_2_o ;
  wire \u_DISPATCH/n1 ;
  wire \u_DISPATCH/n28 ;
  wire \u_DISPATCH/n4 ;
  wire \u_IFU/jump_flag ;  // ../RTL/core/ifu.v(61)
  wire \u_IFU/u_IFU_FETCH/handshake_rdy_last ;  // ../RTL/core/ifu_fetch.v(70)
  wire \u_IFU/u_IFU_FETCH/n7 ;
  wire \u_IFU/u_IFU_FIFO/n13 ;
  wire \u_IFU/u_IFU_FIFO/n9 ;
  wire \u_IFU/u_IFU_PC/add0/c11 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add0/c15 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add0/c19 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add0/c23 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add0/c27 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add0/c3 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add0/c7 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c1 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c11 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c13 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c15 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c17 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c19 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c21 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c23 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c25 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c27 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c29 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c3 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c5 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c7 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/add1/c9 ;  // ../RTL/core/ifu_pc.v(32)
  wire \u_IFU/u_IFU_PC/n7_lutinv ;
  wire \u_IFU/u_IFU_PC/n8 ;
  wire \u_IFU2BPU/fifo_full_lutinv ;  // ../RTL/core/ifu2bpu.v(34)
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_mode ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_wclk ;
  wire \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_we ;
  wire \u_IFU2BPU/u_SYNC_FIFO/eq3/or_or_xor_i0[0]_i1[0_o ;  // ../RTL/core/fifos.v(45)
  wire \u_IFU2BPU/u_SYNC_FIFO/n19 ;
  wire \u_PIPE_CTRL/rs2_match_lutinv ;  // ../RTL/core/pipe_ctrl.v(45)
  wire \u_WB/mux10_b0_sel_is_2_o ;
  wire \u_WB/n1 ;
  wire \u_WB/n15 ;
  wire \u_WB/n16 ;
  wire \u_WB/n2 ;
  wire \u_WB/n37 ;
  wire \u_WB/rdwen0 ;  // ../RTL/core/wb.v(45)
  wire \u_WB/rdwen1 ;  // ../RTL/core/wb.v(46)
  wire \u_WB/rdwen2 ;  // ../RTL/core/wb.v(47)
  wire wb_csr_wen;  // ../RTL/core/ritter_top.v(202)
  wire wb_rdwen;  // ../RTL/core/ritter_top.v(136)

  assign o_ribm_addr0[1] = 1'b0;
  assign o_ribm_addr0[0] = 1'b0;
  assign o_ribm_addr1[1] = 1'b0;
  assign o_ribm_addr1[0] = 1'b0;
  assign o_ribm_mask0[3] = 1'b1;
  assign o_ribm_mask0[2] = 1'b1;
  assign o_ribm_mask0[1] = 1'b1;
  assign o_ribm_mask0[0] = 1'b1;
  assign o_ribm_rdy0 = i_ribm_rsp0;
  assign o_ribm_wdata0[31] = 1'b0;
  assign o_ribm_wdata0[30] = 1'b0;
  assign o_ribm_wdata0[29] = 1'b0;
  assign o_ribm_wdata0[28] = 1'b0;
  assign o_ribm_wdata0[27] = 1'b0;
  assign o_ribm_wdata0[26] = 1'b0;
  assign o_ribm_wdata0[25] = 1'b0;
  assign o_ribm_wdata0[24] = 1'b0;
  assign o_ribm_wdata0[23] = 1'b0;
  assign o_ribm_wdata0[22] = 1'b0;
  assign o_ribm_wdata0[21] = 1'b0;
  assign o_ribm_wdata0[20] = 1'b0;
  assign o_ribm_wdata0[19] = 1'b0;
  assign o_ribm_wdata0[18] = 1'b0;
  assign o_ribm_wdata0[17] = 1'b0;
  assign o_ribm_wdata0[16] = 1'b0;
  assign o_ribm_wdata0[15] = 1'b0;
  assign o_ribm_wdata0[14] = 1'b0;
  assign o_ribm_wdata0[13] = 1'b0;
  assign o_ribm_wdata0[12] = 1'b0;
  assign o_ribm_wdata0[11] = 1'b0;
  assign o_ribm_wdata0[10] = 1'b0;
  assign o_ribm_wdata0[9] = 1'b0;
  assign o_ribm_wdata0[8] = 1'b0;
  assign o_ribm_wdata0[7] = 1'b0;
  assign o_ribm_wdata0[6] = 1'b0;
  assign o_ribm_wdata0[5] = 1'b0;
  assign o_ribm_wdata0[4] = 1'b0;
  assign o_ribm_wdata0[3] = 1'b0;
  assign o_ribm_wdata0[2] = 1'b0;
  assign o_ribm_wdata0[1] = 1'b0;
  assign o_ribm_wdata0[0] = 1'b0;
  assign o_ribm_wrcs0 = 1'b0;
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u456 (
    .a(i_ribm_gnt0),
    .b(i_ribm_rsp0),
    .o(\u_IFU/u_IFU_FIFO/n9 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u457 (
    .a(exu_rdwen0),
    .b(exu_taken_gen),
    .o(\u_WB/n2 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u458 (
    .a(exu_taken),
    .b(exu_taken_gen),
    .o(\u_WB/n37 ));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u459 (
    .a(bpu_taken_gen),
    .b(exu_taken_gen),
    .o(\u_IFU/jump_flag ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u460 (
    .a(bpu_jaddr_gen[10]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[10]),
    .o(\u_IFU/jump_addr [10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u461 (
    .a(bpu_jaddr_gen[11]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[11]),
    .o(\u_IFU/jump_addr [11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u462 (
    .a(bpu_jaddr_gen[12]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[12]),
    .o(\u_IFU/jump_addr [12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u463 (
    .a(bpu_jaddr_gen[13]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[13]),
    .o(\u_IFU/jump_addr [13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u464 (
    .a(bpu_jaddr_gen[14]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[14]),
    .o(\u_IFU/jump_addr [14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u465 (
    .a(bpu_jaddr_gen[15]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[15]),
    .o(\u_IFU/jump_addr [15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u466 (
    .a(bpu_jaddr_gen[16]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[16]),
    .o(\u_IFU/jump_addr [16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u467 (
    .a(bpu_jaddr_gen[17]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[17]),
    .o(\u_IFU/jump_addr [17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u468 (
    .a(bpu_jaddr_gen[18]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[18]),
    .o(\u_IFU/jump_addr [18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u469 (
    .a(bpu_jaddr_gen[19]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[19]),
    .o(\u_IFU/jump_addr [19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u470 (
    .a(bpu_jaddr_gen[2]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[2]),
    .o(\u_IFU/jump_addr [2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u471 (
    .a(bpu_jaddr_gen[20]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[20]),
    .o(\u_IFU/jump_addr [20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u472 (
    .a(bpu_jaddr_gen[21]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[21]),
    .o(\u_IFU/jump_addr [21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u473 (
    .a(bpu_jaddr_gen[22]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[22]),
    .o(\u_IFU/jump_addr [22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u474 (
    .a(bpu_jaddr_gen[23]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[23]),
    .o(\u_IFU/jump_addr [23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u475 (
    .a(bpu_jaddr_gen[24]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[24]),
    .o(\u_IFU/jump_addr [24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u476 (
    .a(bpu_jaddr_gen[25]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[25]),
    .o(\u_IFU/jump_addr [25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u477 (
    .a(bpu_jaddr_gen[26]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[26]),
    .o(\u_IFU/jump_addr [26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u478 (
    .a(bpu_jaddr_gen[27]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[27]),
    .o(\u_IFU/jump_addr [27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u479 (
    .a(bpu_jaddr_gen[28]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[28]),
    .o(\u_IFU/jump_addr [28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u480 (
    .a(bpu_jaddr_gen[29]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[29]),
    .o(\u_IFU/jump_addr [29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u481 (
    .a(bpu_jaddr_gen[3]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[3]),
    .o(\u_IFU/jump_addr [3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u482 (
    .a(bpu_jaddr_gen[30]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[30]),
    .o(\u_IFU/jump_addr [30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u483 (
    .a(bpu_jaddr_gen[31]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[31]),
    .o(\u_IFU/jump_addr [31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u484 (
    .a(bpu_jaddr_gen[4]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[4]),
    .o(\u_IFU/jump_addr [4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u485 (
    .a(bpu_jaddr_gen[5]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[5]),
    .o(\u_IFU/jump_addr [5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u486 (
    .a(bpu_jaddr_gen[6]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[6]),
    .o(\u_IFU/jump_addr [6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u487 (
    .a(bpu_jaddr_gen[7]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[7]),
    .o(\u_IFU/jump_addr [7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u488 (
    .a(bpu_jaddr_gen[8]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[8]),
    .o(\u_IFU/jump_addr [8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u489 (
    .a(bpu_jaddr_gen[9]),
    .b(exu_taken_gen),
    .c(exu_jaddr_gen[9]),
    .o(\u_IFU/jump_addr [9]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*~B*~A)"),
    .INIT(16'hfffe))
    _al_u490 (
    .a(\u_IFU2BPU/fifo_cnt [0]),
    .b(\u_IFU2BPU/fifo_cnt [1]),
    .c(\u_IFU2BPU/fifo_cnt [2]),
    .d(\u_IFU2BPU/fifo_cnt [3]),
    .o(\u_IFU2BPU/u_SYNC_FIFO/eq3/or_or_xor_i0[0]_i1[0_o ));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~B*~A)"),
    .INIT(8'hfe))
    _al_u491 (
    .a(\u_WB/rdwen0 ),
    .b(\u_WB/rdwen1 ),
    .c(\u_WB/rdwen2 ),
    .o(wb_rdwen));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u492 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdidx0 [0]),
    .d(\u_WB/rdidx1 [0]),
    .e(\u_WB/rdidx2 [0]),
    .o(wb_rdidx[0]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u493 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdidx0 [1]),
    .d(\u_WB/rdidx1 [1]),
    .e(\u_WB/rdidx2 [1]),
    .o(wb_rdidx[1]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u494 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdidx0 [2]),
    .d(\u_WB/rdidx1 [2]),
    .e(\u_WB/rdidx2 [2]),
    .o(wb_rdidx[2]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u495 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdidx0 [3]),
    .d(\u_WB/rdidx1 [3]),
    .e(\u_WB/rdidx2 [3]),
    .o(wb_rdidx[3]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u496 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdidx0 [4]),
    .d(\u_WB/rdidx1 [4]),
    .e(\u_WB/rdidx2 [4]),
    .o(wb_rdidx[4]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u497 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [0]),
    .d(\u_WB/rdwdata1 [0]),
    .e(\u_WB/rdwdata2 [0]),
    .o(wb_rdwdata[0]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u498 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [1]),
    .d(\u_WB/rdwdata1 [1]),
    .e(\u_WB/rdwdata2 [1]),
    .o(wb_rdwdata[1]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u499 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [10]),
    .d(\u_WB/rdwdata1 [10]),
    .e(\u_WB/rdwdata2 [10]),
    .o(wb_rdwdata[10]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u500 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [11]),
    .d(\u_WB/rdwdata1 [11]),
    .e(\u_WB/rdwdata2 [11]),
    .o(wb_rdwdata[11]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u501 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [12]),
    .d(\u_WB/rdwdata1 [12]),
    .e(\u_WB/rdwdata2 [12]),
    .o(wb_rdwdata[12]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u502 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [13]),
    .d(\u_WB/rdwdata1 [13]),
    .e(\u_WB/rdwdata2 [13]),
    .o(wb_rdwdata[13]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u503 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [14]),
    .d(\u_WB/rdwdata1 [14]),
    .e(\u_WB/rdwdata2 [14]),
    .o(wb_rdwdata[14]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u504 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [15]),
    .d(\u_WB/rdwdata1 [15]),
    .e(\u_WB/rdwdata2 [15]),
    .o(wb_rdwdata[15]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u505 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [16]),
    .d(\u_WB/rdwdata1 [16]),
    .e(\u_WB/rdwdata2 [16]),
    .o(wb_rdwdata[16]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u506 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [17]),
    .d(\u_WB/rdwdata1 [17]),
    .e(\u_WB/rdwdata2 [17]),
    .o(wb_rdwdata[17]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u507 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [18]),
    .d(\u_WB/rdwdata1 [18]),
    .e(\u_WB/rdwdata2 [18]),
    .o(wb_rdwdata[18]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u508 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [19]),
    .d(\u_WB/rdwdata1 [19]),
    .e(\u_WB/rdwdata2 [19]),
    .o(wb_rdwdata[19]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u509 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [2]),
    .d(\u_WB/rdwdata1 [2]),
    .e(\u_WB/rdwdata2 [2]),
    .o(wb_rdwdata[2]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u510 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [20]),
    .d(\u_WB/rdwdata1 [20]),
    .e(\u_WB/rdwdata2 [20]),
    .o(wb_rdwdata[20]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u511 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [21]),
    .d(\u_WB/rdwdata1 [21]),
    .e(\u_WB/rdwdata2 [21]),
    .o(wb_rdwdata[21]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u512 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [22]),
    .d(\u_WB/rdwdata1 [22]),
    .e(\u_WB/rdwdata2 [22]),
    .o(wb_rdwdata[22]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u513 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [23]),
    .d(\u_WB/rdwdata1 [23]),
    .e(\u_WB/rdwdata2 [23]),
    .o(wb_rdwdata[23]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u514 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [24]),
    .d(\u_WB/rdwdata1 [24]),
    .e(\u_WB/rdwdata2 [24]),
    .o(wb_rdwdata[24]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u515 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [25]),
    .d(\u_WB/rdwdata1 [25]),
    .e(\u_WB/rdwdata2 [25]),
    .o(wb_rdwdata[25]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u516 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [26]),
    .d(\u_WB/rdwdata1 [26]),
    .e(\u_WB/rdwdata2 [26]),
    .o(wb_rdwdata[26]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u517 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [27]),
    .d(\u_WB/rdwdata1 [27]),
    .e(\u_WB/rdwdata2 [27]),
    .o(wb_rdwdata[27]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u518 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [28]),
    .d(\u_WB/rdwdata1 [28]),
    .e(\u_WB/rdwdata2 [28]),
    .o(wb_rdwdata[28]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u519 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [29]),
    .d(\u_WB/rdwdata1 [29]),
    .e(\u_WB/rdwdata2 [29]),
    .o(wb_rdwdata[29]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u520 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [3]),
    .d(\u_WB/rdwdata1 [3]),
    .e(\u_WB/rdwdata2 [3]),
    .o(wb_rdwdata[3]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u521 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [30]),
    .d(\u_WB/rdwdata1 [30]),
    .e(\u_WB/rdwdata2 [30]),
    .o(wb_rdwdata[30]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u522 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [31]),
    .d(\u_WB/rdwdata1 [31]),
    .e(\u_WB/rdwdata2 [31]),
    .o(wb_rdwdata[31]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u523 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [4]),
    .d(\u_WB/rdwdata1 [4]),
    .e(\u_WB/rdwdata2 [4]),
    .o(wb_rdwdata[4]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u524 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [5]),
    .d(\u_WB/rdwdata1 [5]),
    .e(\u_WB/rdwdata2 [5]),
    .o(wb_rdwdata[5]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u525 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [6]),
    .d(\u_WB/rdwdata1 [6]),
    .e(\u_WB/rdwdata2 [6]),
    .o(wb_rdwdata[6]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u526 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [7]),
    .d(\u_WB/rdwdata1 [7]),
    .e(\u_WB/rdwdata2 [7]),
    .o(wb_rdwdata[7]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u527 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [8]),
    .d(\u_WB/rdwdata1 [8]),
    .e(\u_WB/rdwdata2 [8]),
    .o(wb_rdwdata[8]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*~(E)*~(B)+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*~(B)+~((C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))*E*B+(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A)*E*B)"),
    .INIT(32'hfedc3210))
    _al_u528 (
    .a(\u_WB/rdwen1 ),
    .b(\u_WB/rdwen2 ),
    .c(\u_WB/rdwdata0 [9]),
    .d(\u_WB/rdwdata1 [9]),
    .e(\u_WB/rdwdata2 [9]),
    .o(wb_rdwdata[9]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*~(E)*~(D)+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*~(D)+~((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))*E*D+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*D)"),
    .INIT(32'hffd800d8))
    _al_u529 (
    .a(bpu_taken_gen),
    .b(bpu_jaddr_gen[0]),
    .c(\u_IFU/u_IFU_PC/pc [0]),
    .d(exu_taken_gen),
    .e(exu_jaddr_gen[0]),
    .o(\u_IFU/fetch_addr [0]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*~(E)*~(D)+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*~(D)+~((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))*E*D+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*D)"),
    .INIT(32'hffd800d8))
    _al_u530 (
    .a(bpu_taken_gen),
    .b(bpu_jaddr_gen[1]),
    .c(\u_IFU/u_IFU_PC/pc [1]),
    .d(exu_taken_gen),
    .e(exu_jaddr_gen[1]),
    .o(\u_IFU/fetch_addr [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u531 (
    .a(\u_IFU/jump_addr [10]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [10]),
    .o(o_ribm_addr0[10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u532 (
    .a(\u_IFU/jump_addr [11]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [11]),
    .o(o_ribm_addr0[11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u533 (
    .a(\u_IFU/jump_addr [12]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [12]),
    .o(o_ribm_addr0[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u534 (
    .a(\u_IFU/jump_addr [13]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [13]),
    .o(o_ribm_addr0[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u535 (
    .a(\u_IFU/jump_addr [14]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [14]),
    .o(o_ribm_addr0[14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u536 (
    .a(\u_IFU/jump_addr [15]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [15]),
    .o(o_ribm_addr0[15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u537 (
    .a(\u_IFU/jump_addr [16]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [16]),
    .o(o_ribm_addr0[16]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u538 (
    .a(\u_IFU/jump_addr [17]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [17]),
    .o(o_ribm_addr0[17]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u539 (
    .a(\u_IFU/jump_addr [18]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [18]),
    .o(o_ribm_addr0[18]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u540 (
    .a(\u_IFU/jump_addr [19]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [19]),
    .o(o_ribm_addr0[19]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u541 (
    .a(\u_IFU/jump_addr [2]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [2]),
    .o(o_ribm_addr0[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u542 (
    .a(\u_IFU/jump_addr [20]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [20]),
    .o(o_ribm_addr0[20]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u543 (
    .a(\u_IFU/jump_addr [21]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [21]),
    .o(o_ribm_addr0[21]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u544 (
    .a(\u_IFU/jump_addr [22]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [22]),
    .o(o_ribm_addr0[22]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u545 (
    .a(\u_IFU/jump_addr [23]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [23]),
    .o(o_ribm_addr0[23]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*~(E)*~(D)+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*~(D)+~((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))*E*D+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*D)"),
    .INIT(32'hffd800d8))
    _al_u546 (
    .a(bpu_taken_gen),
    .b(bpu_jaddr_gen[24]),
    .c(\u_IFU/u_IFU_PC/pc [24]),
    .d(exu_taken_gen),
    .e(exu_jaddr_gen[24]),
    .o(o_ribm_addr0[24]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*~(E)*~(D)+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*~(D)+~((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))*E*D+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*D)"),
    .INIT(32'hffd800d8))
    _al_u547 (
    .a(bpu_taken_gen),
    .b(bpu_jaddr_gen[25]),
    .c(\u_IFU/u_IFU_PC/pc [25]),
    .d(exu_taken_gen),
    .e(exu_jaddr_gen[25]),
    .o(o_ribm_addr0[25]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*~(E)*~(D)+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*~(D)+~((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))*E*D+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*D)"),
    .INIT(32'hffd800d8))
    _al_u548 (
    .a(bpu_taken_gen),
    .b(bpu_jaddr_gen[26]),
    .c(\u_IFU/u_IFU_PC/pc [26]),
    .d(exu_taken_gen),
    .e(exu_jaddr_gen[26]),
    .o(o_ribm_addr0[26]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*~(E)*~(D)+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*~(D)+~((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))*E*D+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*D)"),
    .INIT(32'hffd800d8))
    _al_u549 (
    .a(bpu_taken_gen),
    .b(bpu_jaddr_gen[27]),
    .c(\u_IFU/u_IFU_PC/pc [27]),
    .d(exu_taken_gen),
    .e(exu_jaddr_gen[27]),
    .o(o_ribm_addr0[27]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*~(E)*~(D)+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*~(D)+~((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))*E*D+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*D)"),
    .INIT(32'hffd800d8))
    _al_u550 (
    .a(bpu_taken_gen),
    .b(bpu_jaddr_gen[28]),
    .c(\u_IFU/u_IFU_PC/pc [28]),
    .d(exu_taken_gen),
    .e(exu_jaddr_gen[28]),
    .o(o_ribm_addr0[28]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*~(E)*~(D)+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*~(D)+~((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))*E*D+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*D)"),
    .INIT(32'hffd800d8))
    _al_u551 (
    .a(bpu_taken_gen),
    .b(bpu_jaddr_gen[29]),
    .c(\u_IFU/u_IFU_PC/pc [29]),
    .d(exu_taken_gen),
    .e(exu_jaddr_gen[29]),
    .o(o_ribm_addr0[29]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u552 (
    .a(\u_IFU/jump_addr [3]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [3]),
    .o(o_ribm_addr0[3]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*~(E)*~(D)+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*~(D)+~((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))*E*D+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*D)"),
    .INIT(32'hffd800d8))
    _al_u553 (
    .a(bpu_taken_gen),
    .b(bpu_jaddr_gen[30]),
    .c(\u_IFU/u_IFU_PC/pc [30]),
    .d(exu_taken_gen),
    .e(exu_jaddr_gen[30]),
    .o(o_ribm_addr0[30]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*~(E)*~(D)+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*~(D)+~((C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))*E*D+(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)*E*D)"),
    .INIT(32'hffd800d8))
    _al_u554 (
    .a(bpu_taken_gen),
    .b(bpu_jaddr_gen[31]),
    .c(\u_IFU/u_IFU_PC/pc [31]),
    .d(exu_taken_gen),
    .e(exu_jaddr_gen[31]),
    .o(o_ribm_addr0[31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u555 (
    .a(\u_IFU/jump_addr [4]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [4]),
    .o(o_ribm_addr0[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u556 (
    .a(\u_IFU/jump_addr [5]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [5]),
    .o(o_ribm_addr0[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u557 (
    .a(\u_IFU/jump_addr [6]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [6]),
    .o(o_ribm_addr0[6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u558 (
    .a(\u_IFU/jump_addr [7]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [7]),
    .o(o_ribm_addr0[7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u559 (
    .a(\u_IFU/jump_addr [8]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [8]),
    .o(o_ribm_addr0[8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u560 (
    .a(\u_IFU/jump_addr [9]),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU/u_IFU_PC/pc [9]),
    .o(o_ribm_addr0[9]));
  AL_MAP_LUT3 #(
    .EQN("~(C@(~B*~A))"),
    .INIT(8'h1e))
    _al_u561 (
    .a(i_ribm_gnt0),
    .b(i_ribm_rsp0),
    .c(\u_IFU/fifo_cnt ),
    .o(\u_IFU/u_IFU_FIFO/n13 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    _al_u562 (
    .a(bpu_inst_vld),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU2BPU/u_SYNC_FIFO/eptr [0]),
    .d(\u_IFU2BPU/u_SYNC_FIFO/eptr [1]),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n23 [1]));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    _al_u563 (
    .a(bpu_inst_vld),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU2BPU/u_SYNC_FIFO/eptr [0]),
    .d(\u_IFU2BPU/u_SYNC_FIFO/eptr [1]),
    .e(\u_IFU2BPU/u_SYNC_FIFO/eptr [2]),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n23 [2]));
  AL_MAP_LUT3 #(
    .EQN("(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'he8))
    _al_u564 (
    .a(\u_WB/rdwen0 ),
    .b(\u_WB/rdwen1 ),
    .c(\u_WB/rdwen2 ),
    .o(_al_u564_o));
  AL_MAP_LUT2 #(
    .EQN("~(~B*A)"),
    .INIT(4'hd))
    _al_u565 (
    .a(_al_u564_o),
    .b(exu_taken_gen),
    .o(\u_WB/n1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u566 (
    .a(\u_WB/n1 ),
    .b(i_rstn),
    .o(\u_WB/mux10_b0_sel_is_2_o ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hbb8a8aaa))
    _al_u567 (
    .a(exu_rdwen1),
    .b(exu_taken_gen),
    .c(\u_WB/rdwen0 ),
    .d(\u_WB/rdwen1 ),
    .e(\u_WB/rdwen2 ),
    .o(\u_WB/n15 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u568 (
    .a(exu_rdwen2),
    .b(\u_WB/n1 ),
    .o(\u_WB/n16 ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u569 (
    .a(ctrl2exu_resource_match),
    .b(_al_u564_o),
    .c(exu_taken_gen),
    .o(n5));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    _al_u570 (
    .a(bpu_inst_vld),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU2BPU/u_SYNC_FIFO/eptr [0]),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n23 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u571 (
    .a(ctrl2exu_rdidx0[4]),
    .b(ctrl2exu_rdidx0[3]),
    .c(ctrl2bpu_rs2idx[4]),
    .d(ctrl2bpu_rs2idx[3]),
    .o(_al_u571_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u572 (
    .a(ctrl2exu_rdidx0[1]),
    .b(ctrl2exu_rdidx0[0]),
    .c(ctrl2bpu_rs2idx[1]),
    .d(ctrl2bpu_rs2idx[0]),
    .o(_al_u572_o));
  AL_MAP_LUT5 #(
    .EQN("(D*B*A*~(E@C))"),
    .INIT(32'h80000800))
    _al_u573 (
    .a(_al_u571_o),
    .b(_al_u572_o),
    .c(ctrl2exu_rdidx0[2]),
    .d(ctrl2exu_rdwen0),
    .e(ctrl2bpu_rs2idx[2]),
    .o(\u_PIPE_CTRL/n9 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u574 (
    .a(ctrl2exu_rdidx2[4]),
    .b(ctrl2exu_rdidx2[3]),
    .c(ctrl2bpu_rs2idx[4]),
    .d(ctrl2bpu_rs2idx[3]),
    .o(_al_u574_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u575 (
    .a(ctrl2exu_rdidx2[1]),
    .b(ctrl2exu_rdidx2[0]),
    .c(ctrl2bpu_rs2idx[1]),
    .d(ctrl2bpu_rs2idx[0]),
    .o(_al_u575_o));
  AL_MAP_LUT5 #(
    .EQN("(D*B*A*~(E@C))"),
    .INIT(32'h80000800))
    _al_u576 (
    .a(_al_u574_o),
    .b(_al_u575_o),
    .c(ctrl2exu_rdidx2[2]),
    .d(ctrl2exu_rdwen2),
    .e(ctrl2bpu_rs2idx[2]),
    .o(\u_PIPE_CTRL/n14 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u577 (
    .a(ctrl2exu_rdidx1[4]),
    .b(ctrl2exu_rdidx1[3]),
    .c(ctrl2bpu_rs2idx[4]),
    .d(ctrl2bpu_rs2idx[3]),
    .o(_al_u577_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u578 (
    .a(ctrl2exu_rdidx1[1]),
    .b(ctrl2exu_rdidx1[0]),
    .c(ctrl2bpu_rs2idx[1]),
    .d(ctrl2bpu_rs2idx[0]),
    .o(_al_u578_o));
  AL_MAP_LUT5 #(
    .EQN("(D*B*A*~(E@C))"),
    .INIT(32'h80000800))
    _al_u579 (
    .a(_al_u577_o),
    .b(_al_u578_o),
    .c(ctrl2exu_rdidx1[2]),
    .d(ctrl2exu_rdwen1),
    .e(ctrl2bpu_rs2idx[2]),
    .o(\u_PIPE_CTRL/n11 [0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u580 (
    .a(\u_PIPE_CTRL/n9 [0]),
    .b(\u_PIPE_CTRL/n14 [0]),
    .c(\u_PIPE_CTRL/n11 [0]),
    .d(ctrl2bpu_rs2ren),
    .o(\u_PIPE_CTRL/rs2_match_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u581 (
    .a(ctrl2exu_rdidx0[4]),
    .b(ctrl2exu_rdidx0[3]),
    .c(ctrl2bpu_rs1idx[4]),
    .d(ctrl2bpu_rs1idx[3]),
    .o(_al_u581_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u582 (
    .a(ctrl2exu_rdidx0[1]),
    .b(ctrl2exu_rdidx0[0]),
    .c(ctrl2bpu_rs1idx[1]),
    .d(ctrl2bpu_rs1idx[0]),
    .o(_al_u582_o));
  AL_MAP_LUT5 #(
    .EQN("(D*B*A*~(E@C))"),
    .INIT(32'h80000800))
    _al_u583 (
    .a(_al_u581_o),
    .b(_al_u582_o),
    .c(ctrl2exu_rdidx0[2]),
    .d(ctrl2exu_rdwen0),
    .e(ctrl2bpu_rs1idx[2]),
    .o(\u_PIPE_CTRL/n1 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u584 (
    .a(ctrl2exu_rdidx2[4]),
    .b(ctrl2exu_rdidx2[3]),
    .c(ctrl2bpu_rs1idx[4]),
    .d(ctrl2bpu_rs1idx[3]),
    .o(_al_u584_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u585 (
    .a(ctrl2exu_rdidx2[1]),
    .b(ctrl2exu_rdidx2[0]),
    .c(ctrl2bpu_rs1idx[1]),
    .d(ctrl2bpu_rs1idx[0]),
    .o(_al_u585_o));
  AL_MAP_LUT5 #(
    .EQN("(D*B*A*~(E@C))"),
    .INIT(32'h80000800))
    _al_u586 (
    .a(_al_u584_o),
    .b(_al_u585_o),
    .c(ctrl2exu_rdidx2[2]),
    .d(ctrl2exu_rdwen2),
    .e(ctrl2bpu_rs1idx[2]),
    .o(\u_PIPE_CTRL/n6 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u587 (
    .a(ctrl2exu_rdidx1[4]),
    .b(ctrl2exu_rdidx1[3]),
    .c(ctrl2bpu_rs1idx[4]),
    .d(ctrl2bpu_rs1idx[3]),
    .o(_al_u587_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u588 (
    .a(ctrl2exu_rdidx1[1]),
    .b(ctrl2exu_rdidx1[0]),
    .c(ctrl2bpu_rs1idx[1]),
    .d(ctrl2bpu_rs1idx[0]),
    .o(_al_u588_o));
  AL_MAP_LUT5 #(
    .EQN("(D*B*A*~(E@C))"),
    .INIT(32'h80000800))
    _al_u589 (
    .a(_al_u587_o),
    .b(_al_u588_o),
    .c(ctrl2exu_rdidx1[2]),
    .d(ctrl2exu_rdwen1),
    .e(ctrl2bpu_rs1idx[2]),
    .o(\u_PIPE_CTRL/n3 [0]));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*~(~D*~C*~B)))"),
    .INIT(32'h00015555))
    _al_u590 (
    .a(\u_PIPE_CTRL/rs2_match_lutinv ),
    .b(\u_PIPE_CTRL/n1 [0]),
    .c(\u_PIPE_CTRL/n6 [0]),
    .d(\u_PIPE_CTRL/n3 [0]),
    .e(ctrl2bpu_rs1ren),
    .o(_al_u590_o));
  AL_MAP_LUT3 #(
    .EQN("~(~C*B*~A)"),
    .INIT(8'hfb))
    _al_u591 (
    .a(ctrl2exu_resource_match),
    .b(_al_u590_o),
    .c(_al_u564_o),
    .o(ctrl2bpu_wait));
  AL_MAP_LUT3 #(
    .EQN("~(~C*~(~B*~A))"),
    .INIT(8'hf1))
    _al_u592 (
    .a(ctrl2exu_resource_match),
    .b(_al_u564_o),
    .c(\u_IFU/jump_flag ),
    .o(\u_DISPATCH/n1 ));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u593 (
    .a(\u_DISPATCH/n1 ),
    .b(_al_u590_o),
    .c(\u_IFU/jump_flag ),
    .o(n3_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u594 (
    .a(bpu_inst_vld),
    .b(n3_lutinv),
    .c(bpu_taken),
    .o(\u_DISPATCH/n28 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u595 (
    .a(bpu_inst_vld),
    .b(n3_lutinv),
    .c(bpu_rdwen),
    .o(\u_DISPATCH/n4 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u596 (
    .a(bpu_inst_vld),
    .b(n3_lutinv),
    .c(bpu_decinfo_grp[5]),
    .o(\u_DISPATCH/n5 [5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u597 (
    .a(bpu_inst_vld),
    .b(n3_lutinv),
    .c(bpu_decinfo_grp[4]),
    .o(\u_DISPATCH/n5 [4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u598 (
    .a(bpu_inst_vld),
    .b(n3_lutinv),
    .c(bpu_decinfo_grp[3]),
    .o(\u_DISPATCH/n5 [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u599 (
    .a(bpu_inst_vld),
    .b(n3_lutinv),
    .c(bpu_decinfo_grp[2]),
    .o(\u_DISPATCH/n5 [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u600 (
    .a(bpu_inst_vld),
    .b(n3_lutinv),
    .c(bpu_decinfo_grp[1]),
    .o(\u_DISPATCH/n5 [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u601 (
    .a(bpu_inst_vld),
    .b(n3_lutinv),
    .c(bpu_decinfo_grp[0]),
    .o(\u_DISPATCH/n5 [0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~(~B*~A)))"),
    .INIT(16'hf100))
    _al_u602 (
    .a(ctrl2exu_resource_match),
    .b(_al_u564_o),
    .c(\u_IFU/jump_flag ),
    .d(i_rstn),
    .o(\u_DISPATCH/mux12_b0_sel_is_2_o ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u603 (
    .a(\u_IFU2BPU/fifo_cnt [0]),
    .b(\u_IFU2BPU/fifo_cnt [1]),
    .c(\u_IFU2BPU/fifo_cnt [2]),
    .o(_al_u603_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u604 (
    .a(_al_u603_o),
    .b(\u_IFU2BPU/fifo_cnt [3]),
    .o(\u_IFU2BPU/fifo_full_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u605 (
    .a(\u_IFU2BPU/fifo_full_lutinv ),
    .b(\u_IFU/jump_flag ),
    .o(_al_u605_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(C*~(~D*B*~A)))"),
    .INIT(32'h0f4f0000))
    _al_u606 (
    .a(ctrl2exu_resource_match),
    .b(_al_u590_o),
    .c(_al_u605_o),
    .d(_al_u564_o),
    .e(i_rstn),
    .o(o_ribm_req0));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u607 (
    .a(ctrl2bpu_wait),
    .b(_al_u605_o),
    .o(\u_IFU/u_IFU_PC/n7_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(~A*~(E*~D*~C)))"),
    .INIT(32'h22232222))
    _al_u608 (
    .a(i_ribm_gnt0),
    .b(\u_IFU/u_IFU_PC/n7_lutinv ),
    .c(i_ribm_rsp0),
    .d(\u_IFU/jump_flag ),
    .e(\u_IFU/u_IFU_FETCH/handshake_rdy_last ),
    .o(\u_IFU/u_IFU_FETCH/n7 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u609 (
    .a(\u_IFU/u_IFU_PC/n7_lutinv ),
    .b(\u_IFU/fifo_cnt ),
    .o(\u_IFU/u_IFU_PC/n8 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u610 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[9]),
    .c(\u_IFU/u_IFU_PC/pc [9]),
    .o(\u_IFU/u_IFU_PC/n9 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u611 (
    .a(\u_IFU/u_IFU_PC/n2 [7]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [9]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u611_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u612 (
    .a(\u_IFU/u_IFU_PC/n9 [9]),
    .b(\u_IFU/u_IFU_PC/n4 [7]),
    .c(_al_u611_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [9]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u613 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[8]),
    .c(\u_IFU/u_IFU_PC/pc [8]),
    .o(\u_IFU/u_IFU_PC/n9 [8]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u614 (
    .a(\u_IFU/u_IFU_PC/n2 [6]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [8]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u614_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u615 (
    .a(\u_IFU/u_IFU_PC/n9 [8]),
    .b(\u_IFU/u_IFU_PC/n4 [6]),
    .c(_al_u614_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u616 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[7]),
    .c(\u_IFU/u_IFU_PC/pc [7]),
    .o(\u_IFU/u_IFU_PC/n9 [7]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u617 (
    .a(\u_IFU/u_IFU_PC/n2 [5]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [7]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u617_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u618 (
    .a(\u_IFU/u_IFU_PC/n9 [7]),
    .b(\u_IFU/u_IFU_PC/n4 [5]),
    .c(_al_u617_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u619 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[6]),
    .c(\u_IFU/u_IFU_PC/pc [6]),
    .o(\u_IFU/u_IFU_PC/n9 [6]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u620 (
    .a(\u_IFU/u_IFU_PC/n2 [4]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [6]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u620_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u621 (
    .a(\u_IFU/u_IFU_PC/n9 [6]),
    .b(\u_IFU/u_IFU_PC/n4 [4]),
    .c(_al_u620_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u622 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[5]),
    .c(\u_IFU/u_IFU_PC/pc [5]),
    .o(\u_IFU/u_IFU_PC/n9 [5]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u623 (
    .a(\u_IFU/u_IFU_PC/n2 [3]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [5]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u623_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u624 (
    .a(\u_IFU/u_IFU_PC/n9 [5]),
    .b(\u_IFU/u_IFU_PC/n4 [3]),
    .c(_al_u623_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u625 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[4]),
    .c(\u_IFU/u_IFU_PC/pc [4]),
    .o(\u_IFU/u_IFU_PC/n9 [4]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u626 (
    .a(\u_IFU/u_IFU_PC/n2 [2]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [4]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u626_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u627 (
    .a(\u_IFU/u_IFU_PC/n9 [4]),
    .b(\u_IFU/u_IFU_PC/n4 [2]),
    .c(_al_u626_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u628 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[31]),
    .c(\u_IFU/u_IFU_PC/pc [31]),
    .o(\u_IFU/u_IFU_PC/n9 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u629 (
    .a(\u_IFU/u_IFU_PC/n2 [29]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [31]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u629_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u630 (
    .a(\u_IFU/u_IFU_PC/n9 [31]),
    .b(\u_IFU/u_IFU_PC/n4 [29]),
    .c(_al_u629_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [31]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u631 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[30]),
    .c(\u_IFU/u_IFU_PC/pc [30]),
    .o(\u_IFU/u_IFU_PC/n9 [30]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u632 (
    .a(\u_IFU/u_IFU_PC/n2 [28]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [30]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u632_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u633 (
    .a(\u_IFU/u_IFU_PC/n9 [30]),
    .b(\u_IFU/u_IFU_PC/n4 [28]),
    .c(_al_u632_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [30]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u634 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[3]),
    .c(\u_IFU/u_IFU_PC/pc [3]),
    .o(\u_IFU/u_IFU_PC/n9 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u635 (
    .a(\u_IFU/u_IFU_PC/n2 [1]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [3]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u635_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u636 (
    .a(\u_IFU/u_IFU_PC/n9 [3]),
    .b(\u_IFU/u_IFU_PC/n4 [1]),
    .c(_al_u635_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u637 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[29]),
    .c(\u_IFU/u_IFU_PC/pc [29]),
    .o(\u_IFU/u_IFU_PC/n9 [29]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u638 (
    .a(\u_IFU/u_IFU_PC/n2 [27]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [29]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u638_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u639 (
    .a(\u_IFU/u_IFU_PC/n9 [29]),
    .b(\u_IFU/u_IFU_PC/n4 [27]),
    .c(_al_u638_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [29]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u640 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[28]),
    .c(\u_IFU/u_IFU_PC/pc [28]),
    .o(\u_IFU/u_IFU_PC/n9 [28]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u641 (
    .a(\u_IFU/u_IFU_PC/n2 [26]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [28]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u641_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u642 (
    .a(\u_IFU/u_IFU_PC/n9 [28]),
    .b(\u_IFU/u_IFU_PC/n4 [26]),
    .c(_al_u641_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [28]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u643 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[27]),
    .c(\u_IFU/u_IFU_PC/pc [27]),
    .o(\u_IFU/u_IFU_PC/n9 [27]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u644 (
    .a(\u_IFU/u_IFU_PC/n2 [25]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [27]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u644_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u645 (
    .a(\u_IFU/u_IFU_PC/n9 [27]),
    .b(\u_IFU/u_IFU_PC/n4 [25]),
    .c(_al_u644_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [27]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u646 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[26]),
    .c(\u_IFU/u_IFU_PC/pc [26]),
    .o(\u_IFU/u_IFU_PC/n9 [26]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u647 (
    .a(\u_IFU/u_IFU_PC/n2 [24]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [26]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u647_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u648 (
    .a(\u_IFU/u_IFU_PC/n9 [26]),
    .b(\u_IFU/u_IFU_PC/n4 [24]),
    .c(_al_u647_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [26]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u649 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[25]),
    .c(\u_IFU/u_IFU_PC/pc [25]),
    .o(\u_IFU/u_IFU_PC/n9 [25]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u650 (
    .a(\u_IFU/u_IFU_PC/n2 [23]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [25]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u650_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u651 (
    .a(\u_IFU/u_IFU_PC/n9 [25]),
    .b(\u_IFU/u_IFU_PC/n4 [23]),
    .c(_al_u650_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [25]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u652 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[24]),
    .c(\u_IFU/u_IFU_PC/pc [24]),
    .o(\u_IFU/u_IFU_PC/n9 [24]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u653 (
    .a(\u_IFU/u_IFU_PC/n2 [22]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [24]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u653_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u654 (
    .a(\u_IFU/u_IFU_PC/n9 [24]),
    .b(\u_IFU/u_IFU_PC/n4 [22]),
    .c(_al_u653_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [24]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u655 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[23]),
    .c(\u_IFU/u_IFU_PC/pc [23]),
    .o(\u_IFU/u_IFU_PC/n9 [23]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u656 (
    .a(\u_IFU/u_IFU_PC/n2 [21]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [23]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u656_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u657 (
    .a(\u_IFU/u_IFU_PC/n9 [23]),
    .b(\u_IFU/u_IFU_PC/n4 [21]),
    .c(_al_u656_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [23]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u658 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[22]),
    .c(\u_IFU/u_IFU_PC/pc [22]),
    .o(\u_IFU/u_IFU_PC/n9 [22]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u659 (
    .a(\u_IFU/u_IFU_PC/n2 [20]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [22]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u659_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u660 (
    .a(\u_IFU/u_IFU_PC/n9 [22]),
    .b(\u_IFU/u_IFU_PC/n4 [20]),
    .c(_al_u659_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [22]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u661 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[21]),
    .c(\u_IFU/u_IFU_PC/pc [21]),
    .o(\u_IFU/u_IFU_PC/n9 [21]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u662 (
    .a(\u_IFU/u_IFU_PC/n2 [19]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [21]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u662_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u663 (
    .a(\u_IFU/u_IFU_PC/n9 [21]),
    .b(\u_IFU/u_IFU_PC/n4 [19]),
    .c(_al_u662_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [21]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u664 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[20]),
    .c(\u_IFU/u_IFU_PC/pc [20]),
    .o(\u_IFU/u_IFU_PC/n9 [20]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u665 (
    .a(\u_IFU/u_IFU_PC/n2 [18]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [20]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u665_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u666 (
    .a(\u_IFU/u_IFU_PC/n9 [20]),
    .b(\u_IFU/u_IFU_PC/n4 [18]),
    .c(_al_u665_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [20]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u667 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[2]),
    .c(\u_IFU/u_IFU_PC/pc [2]),
    .o(_al_u667_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hac0f))
    _al_u668 (
    .a(\u_IFU/u_IFU_PC/n2 [0]),
    .b(\u_IFU/u_IFU_PC/n4 [0]),
    .c(\u_IFU/jump_flag ),
    .d(i_ribm_gnt0),
    .o(_al_u668_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf05c))
    _al_u669 (
    .a(_al_u667_o),
    .b(\u_IFU/jump_addr [2]),
    .c(_al_u668_o),
    .d(i_ribm_gnt0),
    .o(\u_IFU/u_IFU_PC/n10 [2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u670 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[19]),
    .c(\u_IFU/u_IFU_PC/pc [19]),
    .o(\u_IFU/u_IFU_PC/n9 [19]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u671 (
    .a(\u_IFU/u_IFU_PC/n2 [17]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [19]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u671_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u672 (
    .a(\u_IFU/u_IFU_PC/n9 [19]),
    .b(\u_IFU/u_IFU_PC/n4 [17]),
    .c(_al_u671_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [19]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u673 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[18]),
    .c(\u_IFU/u_IFU_PC/pc [18]),
    .o(\u_IFU/u_IFU_PC/n9 [18]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u674 (
    .a(\u_IFU/u_IFU_PC/n2 [16]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [18]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u674_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u675 (
    .a(\u_IFU/u_IFU_PC/n9 [18]),
    .b(\u_IFU/u_IFU_PC/n4 [16]),
    .c(_al_u674_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [18]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u676 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[17]),
    .c(\u_IFU/u_IFU_PC/pc [17]),
    .o(\u_IFU/u_IFU_PC/n9 [17]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u677 (
    .a(\u_IFU/u_IFU_PC/n2 [15]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [17]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u677_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u678 (
    .a(\u_IFU/u_IFU_PC/n9 [17]),
    .b(\u_IFU/u_IFU_PC/n4 [15]),
    .c(_al_u677_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [17]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u679 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[16]),
    .c(\u_IFU/u_IFU_PC/pc [16]),
    .o(\u_IFU/u_IFU_PC/n9 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u680 (
    .a(\u_IFU/u_IFU_PC/n2 [14]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [16]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u680_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u681 (
    .a(\u_IFU/u_IFU_PC/n9 [16]),
    .b(\u_IFU/u_IFU_PC/n4 [14]),
    .c(_al_u680_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [16]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u682 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[15]),
    .c(\u_IFU/u_IFU_PC/pc [15]),
    .o(\u_IFU/u_IFU_PC/n9 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u683 (
    .a(\u_IFU/u_IFU_PC/n2 [13]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [15]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u683_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u684 (
    .a(\u_IFU/u_IFU_PC/n9 [15]),
    .b(\u_IFU/u_IFU_PC/n4 [13]),
    .c(_al_u683_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [15]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u685 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[14]),
    .c(\u_IFU/u_IFU_PC/pc [14]),
    .o(\u_IFU/u_IFU_PC/n9 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u686 (
    .a(\u_IFU/u_IFU_PC/n2 [12]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [14]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u686_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u687 (
    .a(\u_IFU/u_IFU_PC/n9 [14]),
    .b(\u_IFU/u_IFU_PC/n4 [12]),
    .c(_al_u686_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [14]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u688 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[13]),
    .c(\u_IFU/u_IFU_PC/pc [13]),
    .o(\u_IFU/u_IFU_PC/n9 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u689 (
    .a(\u_IFU/u_IFU_PC/n2 [11]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [13]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u689_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u690 (
    .a(\u_IFU/u_IFU_PC/n9 [13]),
    .b(\u_IFU/u_IFU_PC/n4 [11]),
    .c(_al_u689_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [13]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u691 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[12]),
    .c(\u_IFU/u_IFU_PC/pc [12]),
    .o(\u_IFU/u_IFU_PC/n9 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u692 (
    .a(\u_IFU/u_IFU_PC/n2 [10]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [12]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u692_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u693 (
    .a(\u_IFU/u_IFU_PC/n9 [12]),
    .b(\u_IFU/u_IFU_PC/n4 [10]),
    .c(_al_u692_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u694 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[11]),
    .c(\u_IFU/u_IFU_PC/pc [11]),
    .o(\u_IFU/u_IFU_PC/n9 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u695 (
    .a(\u_IFU/u_IFU_PC/n2 [9]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [11]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u695_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u696 (
    .a(\u_IFU/u_IFU_PC/n9 [11]),
    .b(\u_IFU/u_IFU_PC/n4 [9]),
    .c(_al_u695_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [11]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u697 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[10]),
    .c(\u_IFU/u_IFU_PC/pc [10]),
    .o(\u_IFU/u_IFU_PC/n9 [10]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb8cc))
    _al_u698 (
    .a(\u_IFU/u_IFU_PC/n2 [8]),
    .b(i_ribm_gnt0),
    .c(\u_IFU/jump_addr [10]),
    .d(\u_IFU/jump_flag ),
    .o(_al_u698_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u699 (
    .a(\u_IFU/u_IFU_PC/n9 [10]),
    .b(\u_IFU/u_IFU_PC/n4 [8]),
    .c(_al_u698_o),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [10]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u700 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[1]),
    .c(\u_IFU/u_IFU_PC/pc [1]),
    .o(_al_u700_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(B)*~((~D*~A))+~C*B*~((~D*~A))+~(~C)*B*(~D*~A)+~C*B*(~D*~A))"),
    .INIT(16'hf0b1))
    _al_u701 (
    .a(i_ribm_gnt0),
    .b(_al_u700_o),
    .c(\u_IFU/fetch_addr [1]),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u702 (
    .a(\u_IFU/u_IFU_PC/n8 ),
    .b(ifu_iaddr[0]),
    .c(\u_IFU/u_IFU_PC/pc [0]),
    .o(_al_u702_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(B)*~((~D*~A))+~C*B*~((~D*~A))+~(~C)*B*(~D*~A)+~C*B*(~D*~A))"),
    .INIT(16'hf0b1))
    _al_u703 (
    .a(i_ribm_gnt0),
    .b(_al_u702_o),
    .c(\u_IFU/fetch_addr [0]),
    .d(\u_IFU/jump_flag ),
    .o(\u_IFU/u_IFU_PC/n10 [0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u704 (
    .a(i_ribm_rsp0),
    .b(\u_IFU/u_IFU_FETCH/handshake_rdy_last ),
    .c(\u_IFU/fifo_cnt ),
    .o(_al_u704_o));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C*~(~E*B*~A)))"),
    .INIT(32'h0f004f00))
    _al_u705 (
    .a(ctrl2exu_resource_match),
    .b(_al_u590_o),
    .c(_al_u605_o),
    .d(_al_u704_o),
    .e(_al_u564_o),
    .o(ifu_data_vld));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u706 (
    .a(ifu_data_vld),
    .b(\u_IFU/jump_flag ),
    .c(i_rstn),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n19 ));
  AL_MAP_LUT5 #(
    .EQN("(~B*(E@(D*C*A)))"),
    .INIT(32'h13332000))
    _al_u707 (
    .a(ifu_data_vld),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU2BPU/u_SYNC_FIFO/hptr [0]),
    .d(\u_IFU2BPU/u_SYNC_FIFO/hptr [1]),
    .e(\u_IFU2BPU/u_SYNC_FIFO/hptr [2]),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n22 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D@(C*A)))"),
    .INIT(16'h1320))
    _al_u708 (
    .a(ifu_data_vld),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU2BPU/u_SYNC_FIFO/hptr [0]),
    .d(\u_IFU2BPU/u_SYNC_FIFO/hptr [1]),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n22 [1]));
  AL_MAP_LUT3 #(
    .EQN("(~B*(C@A))"),
    .INIT(8'h12))
    _al_u709 (
    .a(ifu_data_vld),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU2BPU/u_SYNC_FIFO/hptr [0]),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n22 [0]));
  AL_MAP_LUT5 #(
    .EQN("(A*(B*C*D*~(E)+B*~(C)*~(D)*E+~(B)*C*~(D)*E+B*C*~(D)*E+~(B)*~(C)*D*E+B*~(C)*D*E+~(B)*C*D*E))"),
    .INIT(32'h2aa88000))
    _al_u710 (
    .a(_al_u704_o),
    .b(\u_IFU2BPU/fifo_cnt [0]),
    .c(\u_IFU2BPU/fifo_cnt [1]),
    .d(\u_IFU2BPU/fifo_cnt [2]),
    .e(\u_IFU2BPU/fifo_cnt [3]),
    .o(_al_u710_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hddfb7270))
    _al_u711 (
    .a(bpu_inst_vld),
    .b(ifu_data_vld),
    .c(_al_u710_o),
    .d(_al_u603_o),
    .e(\u_IFU2BPU/fifo_cnt [3]),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n16 [3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u712 (
    .a(\u_IFU2BPU/u_SYNC_FIFO/n16 [3]),
    .b(\u_IFU/jump_flag ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n24 [3]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hbffd))
    _al_u713 (
    .a(bpu_inst_vld),
    .b(ifu_data_vld),
    .c(\u_IFU2BPU/fifo_cnt [0]),
    .d(\u_IFU2BPU/fifo_cnt [1]),
    .o(_al_u713_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    _al_u714 (
    .a(_al_u713_o),
    .b(\u_IFU/jump_flag ),
    .c(\u_IFU2BPU/fifo_cnt [2]),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n24 [2]));
  AL_MAP_LUT5 #(
    .EQN("(~C*(E@(A*~(B)*~(D)+~(A)*B*D)))"),
    .INIT(32'h0b0d0402))
    _al_u715 (
    .a(bpu_inst_vld),
    .b(ifu_data_vld),
    .c(\u_IFU/jump_flag ),
    .d(\u_IFU2BPU/fifo_cnt [0]),
    .e(\u_IFU2BPU/fifo_cnt [1]),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n24 [1]));
  AL_MAP_LUT5 #(
    .EQN("(~C*(A*~(B)*~(D)*~(E)+~(A)*B*~(D)*~(E)+~(A)*~(B)*D*~(E)+A*B*D*~(E)+A*~(B)*~(D)*E+~(A)*~(B)*D*E+A*B*D*E))"),
    .INIT(32'h09020906))
    _al_u716 (
    .a(bpu_inst_vld),
    .b(ifu_data_vld),
    .c(\u_IFU/jump_flag ),
    .d(\u_IFU2BPU/fifo_cnt [0]),
    .e(\u_IFU2BPU/fifo_full_lutinv ),
    .o(\u_IFU2BPU/u_SYNC_FIFO/n24 [0]));
  BPU u_BPU (
    .i_clk(i_clk),
    .i_data(ifu2bpu_data),
    .i_data_vld(\u_IFU2BPU/u_SYNC_FIFO/eq3/or_or_xor_i0[0]_i1[0_o ),
    .i_flush(\u_IFU/jump_flag ),
    .i_iaddr(ifu2bpu_iaddr),
    .i_rd_wdata(wb_rdwdata),
    .i_rdidx(wb_rdidx),
    .i_rdwen(wb_rdwen),
    .i_rstn(i_rstn),
    .i_stop(ctrl2bpu_wait),
    .o_bpu_jaddr(bpu_jaddr),
    .o_bpu_rs1idx(ctrl2bpu_rs1idx),
    .o_bpu_rs1ren(ctrl2bpu_rs1ren),
    .o_bpu_rs2idx(ctrl2bpu_rs2idx),
    .o_bpu_rs2ren(ctrl2bpu_rs2ren),
    .o_bpu_taken(bpu_taken),
    .o_csr_zimm({open_n1,open_n2,open_n3,open_n4,open_n5,open_n6,open_n7,open_n8,open_n9,open_n10,open_n11,open_n12,open_n13,open_n14,open_n15,open_n16,open_n17,open_n18,open_n19,open_n20,open_n21,open_n22,open_n23,open_n24,open_n25,open_n26,open_n27,bpu_csr_zimm[4:0]}),
    .o_csridx(bpu_csridx),
    .o_decinfo({bpu_decinfo[9:1],open_n28}),
    .o_decinfo_grp(bpu_decinfo_grp),
    .o_exu_op1(bpu_exu_op1),
    .o_exu_op2(bpu_exu_op2),
    .o_iaddr(bpu_iaddr),
    .o_imm(bpu_imm),
    .o_inst_vld(bpu_inst_vld),
    .o_rdidx(bpu_rdidx),
    .o_rdwen(bpu_rdwen),
    .o_rs2rdata(bpu_rs2rdata));  // ../RTL/core/ritter_top.v(157)
  CSR_REGFILE u_CSR_REGFILE (
    .i_clk(i_clk),
    .i_csr_ridx(bpu_csridx),
    .i_csr_wdata(wb_csr_wdata),
    .i_csr_wen(wb_csr_wen),
    .i_csr_widx(wb_csridx),
    .i_rstn(i_rstn),
    .o_csr_rdata(csr_rdata));  // ../RTL/core/ritter_top.v(206)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DISPATCH/o_bpu_taken_reg  (
    .ce(\u_DISPATCH/n1 ),
    .clk(i_clk),
    .d(\u_DISPATCH/n28 ),
    .sr(i_rstn),
    .q(bpu_taken_gen));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DISPATCH/o_rdwen_reg  (
    .ce(\u_DISPATCH/n1 ),
    .clk(i_clk),
    .d(\u_DISPATCH/n4 ),
    .sr(i_rstn),
    .q(dis_rdwen));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DISPATCH/reg0_b0  (
    .ce(\u_DISPATCH/n1 ),
    .clk(i_clk),
    .d(\u_DISPATCH/n5 [0]),
    .sr(i_rstn),
    .q(dis_decinfo_grp[0]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DISPATCH/reg0_b1  (
    .ce(\u_DISPATCH/n1 ),
    .clk(i_clk),
    .d(\u_DISPATCH/n5 [1]),
    .sr(i_rstn),
    .q(dis_decinfo_grp[1]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DISPATCH/reg0_b2  (
    .ce(\u_DISPATCH/n1 ),
    .clk(i_clk),
    .d(\u_DISPATCH/n5 [2]),
    .sr(i_rstn),
    .q(dis_decinfo_grp[2]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DISPATCH/reg0_b3  (
    .ce(\u_DISPATCH/n1 ),
    .clk(i_clk),
    .d(\u_DISPATCH/n5 [3]),
    .sr(i_rstn),
    .q(dis_decinfo_grp[3]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DISPATCH/reg0_b4  (
    .ce(\u_DISPATCH/n1 ),
    .clk(i_clk),
    .d(\u_DISPATCH/n5 [4]),
    .sr(i_rstn),
    .q(dis_decinfo_grp[4]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DISPATCH/reg0_b5  (
    .ce(\u_DISPATCH/n1 ),
    .clk(i_clk),
    .d(\u_DISPATCH/n5 [5]),
    .sr(i_rstn),
    .q(dis_decinfo_grp[5]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b0  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[0]),
    .q(dis_iaddr[0]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b1  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[1]),
    .q(dis_iaddr[1]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b10  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[10]),
    .q(dis_iaddr[10]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b11  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[11]),
    .q(dis_iaddr[11]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b12  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[12]),
    .q(dis_iaddr[12]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b13  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[13]),
    .q(dis_iaddr[13]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b14  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[14]),
    .q(dis_iaddr[14]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b15  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[15]),
    .q(dis_iaddr[15]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b16  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[16]),
    .q(dis_iaddr[16]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b17  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[17]),
    .q(dis_iaddr[17]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b18  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[18]),
    .q(dis_iaddr[18]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b19  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[19]),
    .q(dis_iaddr[19]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b2  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[2]),
    .q(dis_iaddr[2]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b20  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[20]),
    .q(dis_iaddr[20]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b21  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[21]),
    .q(dis_iaddr[21]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b22  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[22]),
    .q(dis_iaddr[22]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b23  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[23]),
    .q(dis_iaddr[23]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b24  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[24]),
    .q(dis_iaddr[24]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b25  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[25]),
    .q(dis_iaddr[25]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b26  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[26]),
    .q(dis_iaddr[26]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b27  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[27]),
    .q(dis_iaddr[27]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b28  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[28]),
    .q(dis_iaddr[28]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b29  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[29]),
    .q(dis_iaddr[29]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b3  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[3]),
    .q(dis_iaddr[3]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b30  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[30]),
    .q(dis_iaddr[30]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b31  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[31]),
    .q(dis_iaddr[31]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b4  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[4]),
    .q(dis_iaddr[4]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b5  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[5]),
    .q(dis_iaddr[5]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b6  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[6]),
    .q(dis_iaddr[6]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b7  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[7]),
    .q(dis_iaddr[7]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b8  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[8]),
    .q(dis_iaddr[8]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg10_b9  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_iaddr[9]),
    .q(dis_iaddr[9]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b0  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[0]),
    .q(bpu_jaddr_gen[0]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b1  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[1]),
    .q(bpu_jaddr_gen[1]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b10  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[10]),
    .q(bpu_jaddr_gen[10]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b11  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[11]),
    .q(bpu_jaddr_gen[11]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b12  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[12]),
    .q(bpu_jaddr_gen[12]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b13  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[13]),
    .q(bpu_jaddr_gen[13]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b14  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[14]),
    .q(bpu_jaddr_gen[14]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b15  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[15]),
    .q(bpu_jaddr_gen[15]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b16  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[16]),
    .q(bpu_jaddr_gen[16]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b17  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[17]),
    .q(bpu_jaddr_gen[17]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b18  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[18]),
    .q(bpu_jaddr_gen[18]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b19  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[19]),
    .q(bpu_jaddr_gen[19]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b2  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[2]),
    .q(bpu_jaddr_gen[2]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b20  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[20]),
    .q(bpu_jaddr_gen[20]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b21  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[21]),
    .q(bpu_jaddr_gen[21]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b22  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[22]),
    .q(bpu_jaddr_gen[22]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b23  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[23]),
    .q(bpu_jaddr_gen[23]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b24  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[24]),
    .q(bpu_jaddr_gen[24]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b25  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[25]),
    .q(bpu_jaddr_gen[25]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b26  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[26]),
    .q(bpu_jaddr_gen[26]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b27  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[27]),
    .q(bpu_jaddr_gen[27]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b28  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[28]),
    .q(bpu_jaddr_gen[28]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b29  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[29]),
    .q(bpu_jaddr_gen[29]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b3  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[3]),
    .q(bpu_jaddr_gen[3]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b30  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[30]),
    .q(bpu_jaddr_gen[30]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b31  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[31]),
    .q(bpu_jaddr_gen[31]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b4  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[4]),
    .q(bpu_jaddr_gen[4]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b5  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[5]),
    .q(bpu_jaddr_gen[5]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b6  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[6]),
    .q(bpu_jaddr_gen[6]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b7  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[7]),
    .q(bpu_jaddr_gen[7]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b8  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[8]),
    .q(bpu_jaddr_gen[8]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg11_b9  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_jaddr[9]),
    .q(bpu_jaddr_gen[9]));  // ../RTL/core/dispatch.v(113)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b0  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[0]),
    .q(dis_exu_op1[0]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b1  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[1]),
    .q(dis_exu_op1[1]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b10  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[10]),
    .q(dis_exu_op1[10]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b11  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[11]),
    .q(dis_exu_op1[11]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b12  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[12]),
    .q(dis_exu_op1[12]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b13  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[13]),
    .q(dis_exu_op1[13]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b14  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[14]),
    .q(dis_exu_op1[14]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b15  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[15]),
    .q(dis_exu_op1[15]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b16  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[16]),
    .q(dis_exu_op1[16]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b17  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[17]),
    .q(dis_exu_op1[17]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b18  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[18]),
    .q(dis_exu_op1[18]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b19  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[19]),
    .q(dis_exu_op1[19]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b2  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[2]),
    .q(dis_exu_op1[2]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b20  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[20]),
    .q(dis_exu_op1[20]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b21  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[21]),
    .q(dis_exu_op1[21]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b22  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[22]),
    .q(dis_exu_op1[22]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b23  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[23]),
    .q(dis_exu_op1[23]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b24  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[24]),
    .q(dis_exu_op1[24]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b25  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[25]),
    .q(dis_exu_op1[25]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b26  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[26]),
    .q(dis_exu_op1[26]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b27  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[27]),
    .q(dis_exu_op1[27]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b28  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[28]),
    .q(dis_exu_op1[28]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b29  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[29]),
    .q(dis_exu_op1[29]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b3  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[3]),
    .q(dis_exu_op1[3]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b30  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[30]),
    .q(dis_exu_op1[30]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b31  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[31]),
    .q(dis_exu_op1[31]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b4  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[4]),
    .q(dis_exu_op1[4]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b5  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[5]),
    .q(dis_exu_op1[5]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b6  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[6]),
    .q(dis_exu_op1[6]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b7  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[7]),
    .q(dis_exu_op1[7]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b8  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[8]),
    .q(dis_exu_op1[8]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg1_b9  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op1[9]),
    .q(dis_exu_op1[9]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b0  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[0]),
    .q(dis_exu_op2[0]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b1  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[1]),
    .q(dis_exu_op2[1]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b10  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[10]),
    .q(dis_exu_op2[10]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b11  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[11]),
    .q(dis_exu_op2[11]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b12  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[12]),
    .q(dis_exu_op2[12]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b13  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[13]),
    .q(dis_exu_op2[13]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b14  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[14]),
    .q(dis_exu_op2[14]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b15  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[15]),
    .q(dis_exu_op2[15]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b16  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[16]),
    .q(dis_exu_op2[16]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b17  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[17]),
    .q(dis_exu_op2[17]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b18  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[18]),
    .q(dis_exu_op2[18]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b19  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[19]),
    .q(dis_exu_op2[19]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b2  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[2]),
    .q(dis_exu_op2[2]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b20  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[20]),
    .q(dis_exu_op2[20]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b21  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[21]),
    .q(dis_exu_op2[21]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b22  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[22]),
    .q(dis_exu_op2[22]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b23  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[23]),
    .q(dis_exu_op2[23]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b24  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[24]),
    .q(dis_exu_op2[24]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b25  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[25]),
    .q(dis_exu_op2[25]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b26  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[26]),
    .q(dis_exu_op2[26]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b27  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[27]),
    .q(dis_exu_op2[27]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b28  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[28]),
    .q(dis_exu_op2[28]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b29  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[29]),
    .q(dis_exu_op2[29]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b3  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[3]),
    .q(dis_exu_op2[3]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b30  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[30]),
    .q(dis_exu_op2[30]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b31  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[31]),
    .q(dis_exu_op2[31]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b4  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[4]),
    .q(dis_exu_op2[4]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b5  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[5]),
    .q(dis_exu_op2[5]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b6  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[6]),
    .q(dis_exu_op2[6]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b7  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[7]),
    .q(dis_exu_op2[7]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b8  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[8]),
    .q(dis_exu_op2[8]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg2_b9  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_exu_op2[9]),
    .q(dis_exu_op2[9]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b0  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[0]),
    .q(dis_rs2rdata[0]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b1  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[1]),
    .q(dis_rs2rdata[1]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b10  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[10]),
    .q(dis_rs2rdata[10]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b11  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[11]),
    .q(dis_rs2rdata[11]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b12  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[12]),
    .q(dis_rs2rdata[12]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b13  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[13]),
    .q(dis_rs2rdata[13]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b14  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[14]),
    .q(dis_rs2rdata[14]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b15  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[15]),
    .q(dis_rs2rdata[15]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b16  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[16]),
    .q(dis_rs2rdata[16]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b17  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[17]),
    .q(dis_rs2rdata[17]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b18  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[18]),
    .q(dis_rs2rdata[18]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b19  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[19]),
    .q(dis_rs2rdata[19]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b2  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[2]),
    .q(dis_rs2rdata[2]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b20  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[20]),
    .q(dis_rs2rdata[20]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b21  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[21]),
    .q(dis_rs2rdata[21]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b22  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[22]),
    .q(dis_rs2rdata[22]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b23  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[23]),
    .q(dis_rs2rdata[23]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b24  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[24]),
    .q(dis_rs2rdata[24]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b25  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[25]),
    .q(dis_rs2rdata[25]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b26  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[26]),
    .q(dis_rs2rdata[26]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b27  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[27]),
    .q(dis_rs2rdata[27]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b28  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[28]),
    .q(dis_rs2rdata[28]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b29  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[29]),
    .q(dis_rs2rdata[29]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b3  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[3]),
    .q(dis_rs2rdata[3]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b30  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[30]),
    .q(dis_rs2rdata[30]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b31  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[31]),
    .q(dis_rs2rdata[31]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b4  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[4]),
    .q(dis_rs2rdata[4]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b5  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[5]),
    .q(dis_rs2rdata[5]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b6  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[6]),
    .q(dis_rs2rdata[6]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b7  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[7]),
    .q(dis_rs2rdata[7]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b8  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[8]),
    .q(dis_rs2rdata[8]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg3_b9  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rs2rdata[9]),
    .q(dis_rs2rdata[9]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b0  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[0]),
    .q(dis_imm[0]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b1  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[1]),
    .q(dis_imm[1]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b10  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[10]),
    .q(dis_imm[10]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b11  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[11]),
    .q(dis_imm[11]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b12  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[12]),
    .q(dis_imm[12]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b13  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[13]),
    .q(dis_imm[13]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b14  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[14]),
    .q(dis_imm[14]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b15  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[15]),
    .q(dis_imm[15]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b16  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[16]),
    .q(dis_imm[16]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b17  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[17]),
    .q(dis_imm[17]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b18  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[18]),
    .q(dis_imm[18]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b19  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[19]),
    .q(dis_imm[19]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b2  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[2]),
    .q(dis_imm[2]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b20  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[20]),
    .q(dis_imm[20]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b21  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[21]),
    .q(dis_imm[21]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b22  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[22]),
    .q(dis_imm[22]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b23  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[23]),
    .q(dis_imm[23]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b24  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[24]),
    .q(dis_imm[24]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b25  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[25]),
    .q(dis_imm[25]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b26  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[26]),
    .q(dis_imm[26]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b27  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[27]),
    .q(dis_imm[27]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b28  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[28]),
    .q(dis_imm[28]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b29  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[29]),
    .q(dis_imm[29]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b3  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[3]),
    .q(dis_imm[3]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b30  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[30]),
    .q(dis_imm[30]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b31  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[31]),
    .q(dis_imm[31]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b4  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[4]),
    .q(dis_imm[4]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b5  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[5]),
    .q(dis_imm[5]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b6  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[6]),
    .q(dis_imm[6]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b7  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[7]),
    .q(dis_imm[7]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b8  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[8]),
    .q(dis_imm[8]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg4_b9  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_imm[9]),
    .q(dis_imm[9]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg5_b0  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rdidx[0]),
    .q(dis_rdidx[0]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg5_b1  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rdidx[1]),
    .q(dis_rdidx[1]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg5_b2  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rdidx[2]),
    .q(dis_rdidx[2]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg5_b3  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rdidx[3]),
    .q(dis_rdidx[3]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg5_b4  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_rdidx[4]),
    .q(dis_rdidx[4]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg6_b0  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csridx[0]),
    .q(dis_csridx[0]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg6_b1  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csridx[1]),
    .q(dis_csridx[1]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg6_b10  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csridx[10]),
    .q(dis_csridx[10]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg6_b11  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csridx[11]),
    .q(dis_csridx[11]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg6_b2  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csridx[2]),
    .q(dis_csridx[2]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg6_b3  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csridx[3]),
    .q(dis_csridx[3]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg6_b4  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csridx[4]),
    .q(dis_csridx[4]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg6_b5  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csridx[5]),
    .q(dis_csridx[5]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg6_b6  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csridx[6]),
    .q(dis_csridx[6]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg6_b7  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csridx[7]),
    .q(dis_csridx[7]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg6_b8  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csridx[8]),
    .q(dis_csridx[8]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg6_b9  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csridx[9]),
    .q(dis_csridx[9]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b0  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[0]),
    .q(dis_csr_rdata[0]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b1  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[1]),
    .q(dis_csr_rdata[1]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b10  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[10]),
    .q(dis_csr_rdata[10]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b11  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[11]),
    .q(dis_csr_rdata[11]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b12  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[12]),
    .q(dis_csr_rdata[12]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b13  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[13]),
    .q(dis_csr_rdata[13]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b14  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[14]),
    .q(dis_csr_rdata[14]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b15  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[15]),
    .q(dis_csr_rdata[15]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b16  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[16]),
    .q(dis_csr_rdata[16]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b17  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[17]),
    .q(dis_csr_rdata[17]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b18  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[18]),
    .q(dis_csr_rdata[18]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b19  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[19]),
    .q(dis_csr_rdata[19]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b2  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[2]),
    .q(dis_csr_rdata[2]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b20  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[20]),
    .q(dis_csr_rdata[20]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b21  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[21]),
    .q(dis_csr_rdata[21]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b22  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[22]),
    .q(dis_csr_rdata[22]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b23  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[23]),
    .q(dis_csr_rdata[23]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b24  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[24]),
    .q(dis_csr_rdata[24]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b25  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[25]),
    .q(dis_csr_rdata[25]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b26  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[26]),
    .q(dis_csr_rdata[26]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b27  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[27]),
    .q(dis_csr_rdata[27]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b28  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[28]),
    .q(dis_csr_rdata[28]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b29  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[29]),
    .q(dis_csr_rdata[29]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b3  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[3]),
    .q(dis_csr_rdata[3]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b30  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[30]),
    .q(dis_csr_rdata[30]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b31  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[31]),
    .q(dis_csr_rdata[31]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b4  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[4]),
    .q(dis_csr_rdata[4]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b5  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[5]),
    .q(dis_csr_rdata[5]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b6  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[6]),
    .q(dis_csr_rdata[6]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b7  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[7]),
    .q(dis_csr_rdata[7]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b8  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[8]),
    .q(dis_csr_rdata[8]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg7_b9  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(csr_rdata[9]),
    .q(dis_csr_rdata[9]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg8_b0  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csr_zimm[0]),
    .q(dis_csr_zimm[0]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg8_b1  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csr_zimm[1]),
    .q(dis_csr_zimm[1]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg8_b2  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csr_zimm[2]),
    .q(dis_csr_zimm[2]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg8_b3  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csr_zimm[3]),
    .q(dis_csr_zimm[3]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg8_b4  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_csr_zimm[4]),
    .q(dis_csr_zimm[4]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg9_b1  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_decinfo[1]),
    .q(dis_decinfo[1]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg9_b2  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_decinfo[2]),
    .q(dis_decinfo[2]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg9_b3  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_decinfo[3]),
    .q(dis_decinfo[3]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg9_b4  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_decinfo[4]),
    .q(dis_decinfo[4]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg9_b5  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_decinfo[5]),
    .q(dis_decinfo[5]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg9_b6  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_decinfo[6]),
    .q(dis_decinfo[6]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg9_b7  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_decinfo[7]),
    .q(dis_decinfo[7]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg9_b8  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_decinfo[8]),
    .q(dis_decinfo[8]));  // ../RTL/core/dispatch.v(90)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DISPATCH/reg9_b9  (
    .ce(\u_DISPATCH/mux12_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(bpu_decinfo[9]),
    .q(dis_decinfo[9]));  // ../RTL/core/dispatch.v(90)
  EXU u_EXU (
    .i_clk(i_clk),
    .i_csr_rdata(dis_csr_rdata),
    .i_csr_zimm({27'b000000000000000000000000000,dis_csr_zimm[4:0]}),
    .i_csridx(dis_csridx),
    .i_decinfo({dis_decinfo[9:1],1'b0}),
    .i_decinfo_grp(dis_decinfo_grp),
    .i_exu_op1(dis_exu_op1),
    .i_exu_op2(dis_exu_op2),
    .i_iaddr(dis_iaddr),
    .i_imm(dis_imm),
    .i_rdidx(dis_rdidx),
    .i_rdwen(dis_rdwen),
    .i_ribm_gnt(i_ribm_gnt1),
    .i_ribm_rdata(i_ribm_rdata1),
    .i_ribm_rsp(i_ribm_rsp1),
    .i_rs2rdata(dis_rs2rdata),
    .i_rstn(i_rstn),
    .i_vld(n5),
    .o_csr_wdata(wb_csr_wdata),
    .o_csr_wen(wb_csr_wen),
    .o_csridx(wb_csridx),
    .o_exu_jaddr(exu_jaddr),
    .o_exu_rdidx0(ctrl2exu_rdidx0),
    .o_exu_rdidx1(ctrl2exu_rdidx1),
    .o_exu_rdidx2(ctrl2exu_rdidx2),
    .o_exu_rdwen0(ctrl2exu_rdwen0),
    .o_exu_rdwen1(ctrl2exu_rdwen1),
    .o_exu_rdwen2(ctrl2exu_rdwen2),
    .o_exu_resource_match(ctrl2exu_resource_match),
    .o_exu_taken(exu_taken),
    .o_rdidx0(exu_rdidx0),
    .o_rdidx1(exu_rdidx1),
    .o_rdidx2(exu_rdidx2),
    .o_rdwdata0(exu_rdwdata0),
    .o_rdwdata1(exu_rdwdata1),
    .o_rdwdata2(exu_rdwdata2),
    .o_rdwen0(exu_rdwen0),
    .o_rdwen1(exu_rdwen1),
    .o_rdwen2(exu_rdwen2),
    .o_ribm_addr({o_ribm_addr1[31:24],open_n287,open_n288,open_n289,open_n290,open_n291,open_n292,open_n293,open_n294,o_ribm_addr1[15:2],open_n295,open_n296}),
    .o_ribm_mask(o_ribm_mask1),
    .o_ribm_req(o_ribm_req1),
    .o_ribm_wdata(o_ribm_wdata1),
    .o_ribm_wrcs(o_ribm_wrcs1));  // ../RTL/core/ritter_top.v(297)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_FETCH/handshake_rdy_last_reg  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_FETCH/n7 ),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_FETCH/handshake_rdy_last ));  // ../RTL/core/ifu_fetch.v(75)
  AL_MAP_SEQ #(
    .CEMUX("INV"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_FIFO/o_fifo_cnt_reg[0]  (
    .ce(\u_IFU/u_IFU_FIFO/n9 ),
    .clk(i_clk),
    .d(\u_IFU/u_IFU_FIFO/n13 ),
    .sr(i_rstn),
    .q(\u_IFU/fifo_cnt ));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b0  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(\u_IFU/fetch_addr [0]),
    .q(ifu_iaddr[0]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b1  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(\u_IFU/fetch_addr [1]),
    .q(ifu_iaddr[1]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b10  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[10]),
    .q(ifu_iaddr[10]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b11  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[11]),
    .q(ifu_iaddr[11]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b12  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[12]),
    .q(ifu_iaddr[12]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b13  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[13]),
    .q(ifu_iaddr[13]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b14  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[14]),
    .q(ifu_iaddr[14]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b15  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[15]),
    .q(ifu_iaddr[15]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b16  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[16]),
    .q(ifu_iaddr[16]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b17  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[17]),
    .q(ifu_iaddr[17]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b18  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[18]),
    .q(ifu_iaddr[18]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b19  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[19]),
    .q(ifu_iaddr[19]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b2  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[2]),
    .q(ifu_iaddr[2]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b20  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[20]),
    .q(ifu_iaddr[20]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b21  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[21]),
    .q(ifu_iaddr[21]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b22  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[22]),
    .q(ifu_iaddr[22]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b23  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[23]),
    .q(ifu_iaddr[23]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b24  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[24]),
    .q(ifu_iaddr[24]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b25  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[25]),
    .q(ifu_iaddr[25]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b26  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[26]),
    .q(ifu_iaddr[26]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b27  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[27]),
    .q(ifu_iaddr[27]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b28  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[28]),
    .q(ifu_iaddr[28]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b29  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[29]),
    .q(ifu_iaddr[29]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b3  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[3]),
    .q(ifu_iaddr[3]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b30  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[30]),
    .q(ifu_iaddr[30]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b31  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[31]),
    .q(ifu_iaddr[31]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b4  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[4]),
    .q(ifu_iaddr[4]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b5  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[5]),
    .q(ifu_iaddr[5]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b6  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[6]),
    .q(ifu_iaddr[6]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b7  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[7]),
    .q(ifu_iaddr[7]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b8  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[8]),
    .q(ifu_iaddr[8]));  // ../RTL/core/fifos.v(131)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_IFU/u_IFU_FIFO/reg0_b9  (
    .ce(i_ribm_gnt0),
    .clk(i_clk),
    .d(o_ribm_addr0[9]),
    .q(ifu_iaddr[9]));  // ../RTL/core/fifos.v(131)
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add0/ucin_al_u717"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add0/u11_al_u720  (
    .a({\u_IFU/jump_addr [15],\u_IFU/jump_addr [13]}),
    .b({\u_IFU/jump_addr [16],\u_IFU/jump_addr [14]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_IFU/u_IFU_PC/add0/c11 ),
    .f({\u_IFU/u_IFU_PC/n2 [13],\u_IFU/u_IFU_PC/n2 [11]}),
    .fco(\u_IFU/u_IFU_PC/add0/c15 ),
    .fx({\u_IFU/u_IFU_PC/n2 [14],\u_IFU/u_IFU_PC/n2 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add0/ucin_al_u717"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add0/u15_al_u721  (
    .a({\u_IFU/jump_addr [19],\u_IFU/jump_addr [17]}),
    .b({\u_IFU/jump_addr [20],\u_IFU/jump_addr [18]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_IFU/u_IFU_PC/add0/c15 ),
    .f({\u_IFU/u_IFU_PC/n2 [17],\u_IFU/u_IFU_PC/n2 [15]}),
    .fco(\u_IFU/u_IFU_PC/add0/c19 ),
    .fx({\u_IFU/u_IFU_PC/n2 [18],\u_IFU/u_IFU_PC/n2 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add0/ucin_al_u717"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add0/u19_al_u722  (
    .a({\u_IFU/jump_addr [23],\u_IFU/jump_addr [21]}),
    .b({\u_IFU/jump_addr [24],\u_IFU/jump_addr [22]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_IFU/u_IFU_PC/add0/c19 ),
    .f({\u_IFU/u_IFU_PC/n2 [21],\u_IFU/u_IFU_PC/n2 [19]}),
    .fco(\u_IFU/u_IFU_PC/add0/c23 ),
    .fx({\u_IFU/u_IFU_PC/n2 [22],\u_IFU/u_IFU_PC/n2 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add0/ucin_al_u717"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add0/u23_al_u723  (
    .a({\u_IFU/jump_addr [27],\u_IFU/jump_addr [25]}),
    .b({\u_IFU/jump_addr [28],\u_IFU/jump_addr [26]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_IFU/u_IFU_PC/add0/c23 ),
    .f({\u_IFU/u_IFU_PC/n2 [25],\u_IFU/u_IFU_PC/n2 [23]}),
    .fco(\u_IFU/u_IFU_PC/add0/c27 ),
    .fx({\u_IFU/u_IFU_PC/n2 [26],\u_IFU/u_IFU_PC/n2 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add0/ucin_al_u717"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add0/u27_al_u724  (
    .a({\u_IFU/jump_addr [31],\u_IFU/jump_addr [29]}),
    .b({open_n403,\u_IFU/jump_addr [30]}),
    .c(2'b00),
    .d(2'b00),
    .e({open_n406,1'b0}),
    .fci(\u_IFU/u_IFU_PC/add0/c27 ),
    .f({\u_IFU/u_IFU_PC/n2 [29],\u_IFU/u_IFU_PC/n2 [27]}),
    .fx({open_n422,\u_IFU/u_IFU_PC/n2 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add0/ucin_al_u717"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add0/u3_al_u718  (
    .a({\u_IFU/jump_addr [7],\u_IFU/jump_addr [5]}),
    .b({\u_IFU/jump_addr [8],\u_IFU/jump_addr [6]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_IFU/u_IFU_PC/add0/c3 ),
    .f({\u_IFU/u_IFU_PC/n2 [5],\u_IFU/u_IFU_PC/n2 [3]}),
    .fco(\u_IFU/u_IFU_PC/add0/c7 ),
    .fx({\u_IFU/u_IFU_PC/n2 [6],\u_IFU/u_IFU_PC/n2 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add0/ucin_al_u717"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add0/u7_al_u719  (
    .a({\u_IFU/jump_addr [11],\u_IFU/jump_addr [9]}),
    .b({\u_IFU/jump_addr [12],\u_IFU/jump_addr [10]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_IFU/u_IFU_PC/add0/c7 ),
    .f({\u_IFU/u_IFU_PC/n2 [9],\u_IFU/u_IFU_PC/n2 [7]}),
    .fco(\u_IFU/u_IFU_PC/add0/c11 ),
    .fx({\u_IFU/u_IFU_PC/n2 [10],\u_IFU/u_IFU_PC/n2 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add0/ucin_al_u717"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add0/ucin_al_u717  (
    .a({\u_IFU/jump_addr [3],1'b0}),
    .b({\u_IFU/jump_addr [4],\u_IFU/jump_addr [2]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({\u_IFU/u_IFU_PC/n2 [1],open_n478}),
    .fco(\u_IFU/u_IFU_PC/add0/c3 ),
    .fx({\u_IFU/u_IFU_PC/n2 [2],\u_IFU/u_IFU_PC/n2 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin  (
    .a({\u_IFU/u_IFU_PC/pc [2],1'b0}),
    .b({1'b1,open_n481}),
    .f({\u_IFU/u_IFU_PC/n4 [0],open_n501}),
    .fco(\u_IFU/u_IFU_PC/add1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u10|u_IFU/u_IFU_PC/add1/u9  (
    .a(\u_IFU/u_IFU_PC/pc [12:11]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c9 ),
    .f(\u_IFU/u_IFU_PC/n4 [10:9]),
    .fco(\u_IFU/u_IFU_PC/add1/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u12|u_IFU/u_IFU_PC/add1/u11  (
    .a(\u_IFU/u_IFU_PC/pc [14:13]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c11 ),
    .f(\u_IFU/u_IFU_PC/n4 [12:11]),
    .fco(\u_IFU/u_IFU_PC/add1/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u14|u_IFU/u_IFU_PC/add1/u13  (
    .a(\u_IFU/u_IFU_PC/pc [16:15]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c13 ),
    .f(\u_IFU/u_IFU_PC/n4 [14:13]),
    .fco(\u_IFU/u_IFU_PC/add1/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u16|u_IFU/u_IFU_PC/add1/u15  (
    .a(\u_IFU/u_IFU_PC/pc [18:17]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c15 ),
    .f(\u_IFU/u_IFU_PC/n4 [16:15]),
    .fco(\u_IFU/u_IFU_PC/add1/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u18|u_IFU/u_IFU_PC/add1/u17  (
    .a(\u_IFU/u_IFU_PC/pc [20:19]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c17 ),
    .f(\u_IFU/u_IFU_PC/n4 [18:17]),
    .fco(\u_IFU/u_IFU_PC/add1/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u20|u_IFU/u_IFU_PC/add1/u19  (
    .a(\u_IFU/u_IFU_PC/pc [22:21]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c19 ),
    .f(\u_IFU/u_IFU_PC/n4 [20:19]),
    .fco(\u_IFU/u_IFU_PC/add1/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u22|u_IFU/u_IFU_PC/add1/u21  (
    .a(\u_IFU/u_IFU_PC/pc [24:23]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c21 ),
    .f(\u_IFU/u_IFU_PC/n4 [22:21]),
    .fco(\u_IFU/u_IFU_PC/add1/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u24|u_IFU/u_IFU_PC/add1/u23  (
    .a(\u_IFU/u_IFU_PC/pc [26:25]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c23 ),
    .f(\u_IFU/u_IFU_PC/n4 [24:23]),
    .fco(\u_IFU/u_IFU_PC/add1/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u26|u_IFU/u_IFU_PC/add1/u25  (
    .a(\u_IFU/u_IFU_PC/pc [28:27]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c25 ),
    .f(\u_IFU/u_IFU_PC/n4 [26:25]),
    .fco(\u_IFU/u_IFU_PC/add1/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u28|u_IFU/u_IFU_PC/add1/u27  (
    .a(\u_IFU/u_IFU_PC/pc [30:29]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c27 ),
    .f(\u_IFU/u_IFU_PC/n4 [28:27]),
    .fco(\u_IFU/u_IFU_PC/add1/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u29_al_u725  (
    .a({open_n726,\u_IFU/u_IFU_PC/pc [31]}),
    .b({open_n727,1'b0}),
    .fci(\u_IFU/u_IFU_PC/add1/c29 ),
    .f({open_n746,\u_IFU/u_IFU_PC/n4 [29]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u2|u_IFU/u_IFU_PC/add1/u1  (
    .a(\u_IFU/u_IFU_PC/pc [4:3]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c1 ),
    .f(\u_IFU/u_IFU_PC/n4 [2:1]),
    .fco(\u_IFU/u_IFU_PC/add1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u4|u_IFU/u_IFU_PC/add1/u3  (
    .a(\u_IFU/u_IFU_PC/pc [6:5]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c3 ),
    .f(\u_IFU/u_IFU_PC/n4 [4:3]),
    .fco(\u_IFU/u_IFU_PC/add1/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u6|u_IFU/u_IFU_PC/add1/u5  (
    .a(\u_IFU/u_IFU_PC/pc [8:7]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c5 ),
    .f(\u_IFU/u_IFU_PC/n4 [6:5]),
    .fco(\u_IFU/u_IFU_PC/add1/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU/u_IFU_PC/add1/u0|u_IFU/u_IFU_PC/add1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_IFU/u_IFU_PC/add1/u8|u_IFU/u_IFU_PC/add1/u7  (
    .a(\u_IFU/u_IFU_PC/pc [10:9]),
    .b(2'b00),
    .fci(\u_IFU/u_IFU_PC/add1/c7 ),
    .f(\u_IFU/u_IFU_PC/n4 [8:7]),
    .fco(\u_IFU/u_IFU_PC/add1/c9 ));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b0  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [0]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [0]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b1  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [1]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [1]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b10  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [10]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [10]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b11  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [11]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [11]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b12  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [12]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [12]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b13  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [13]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [13]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b14  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [14]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [14]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b15  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [15]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [15]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b16  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [16]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [16]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b17  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [17]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [17]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b18  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [18]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [18]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b19  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [19]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [19]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b2  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [2]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [2]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b20  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [20]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [20]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b21  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [21]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [21]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b22  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [22]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [22]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b23  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [23]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [23]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b24  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [24]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [24]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b25  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [25]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [25]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b26  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [26]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [26]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b27  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [27]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [27]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b28  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [28]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [28]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b29  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [29]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [29]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b3  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [3]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [3]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b30  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [30]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [30]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b31  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [31]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [31]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b4  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [4]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [4]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b5  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [5]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [5]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b6  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [6]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [6]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b7  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [7]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [7]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b8  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [8]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [8]));  // ../RTL/core/ifu_pc.v(26)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU/u_IFU_PC/reg0_b9  (
    .clk(i_clk),
    .d(\u_IFU/u_IFU_PC/n10 [9]),
    .sr(i_rstn),
    .q(\u_IFU/u_IFU_PC/pc [9]));  // ../RTL/core/ifu_pc.v(26)
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_l  (
    .a({ifu_iaddr[0],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({ifu_iaddr[1],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({ifu_iaddr[2],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({ifu_iaddr[3],1'b0}),
    .e({open_n873,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_we ),
    .f(ifu2bpu_iaddr[1:0]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c0_we ),
    .f(ifu2bpu_iaddr[3:2]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_l  (
    .a({i_ribm_rdata0[8],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({i_ribm_rdata0[9],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({i_ribm_rdata0[10],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({i_ribm_rdata0[11],1'b0}),
    .e({open_n908,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_we ),
    .f(ifu2bpu_data[9:8]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c10_we ),
    .f(ifu2bpu_data[11:10]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_l  (
    .a({i_ribm_rdata0[12],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({i_ribm_rdata0[13],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({i_ribm_rdata0[14],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({i_ribm_rdata0[15],1'b0}),
    .e({open_n943,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_we ),
    .f(ifu2bpu_data[13:12]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c11_we ),
    .f(ifu2bpu_data[15:14]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_l  (
    .a({i_ribm_rdata0[16],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({i_ribm_rdata0[17],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({i_ribm_rdata0[18],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({i_ribm_rdata0[19],1'b0}),
    .e({open_n978,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_we ),
    .f(ifu2bpu_data[17:16]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c12_we ),
    .f(ifu2bpu_data[19:18]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_l  (
    .a({i_ribm_rdata0[20],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({i_ribm_rdata0[21],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({i_ribm_rdata0[22],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({i_ribm_rdata0[23],1'b0}),
    .e({open_n1013,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_we ),
    .f(ifu2bpu_data[21:20]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c13_we ),
    .f(ifu2bpu_data[23:22]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_l  (
    .a({i_ribm_rdata0[24],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({i_ribm_rdata0[25],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({i_ribm_rdata0[26],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({i_ribm_rdata0[27],1'b0}),
    .e({open_n1048,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_we ),
    .f(ifu2bpu_data[25:24]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c14_we ),
    .f(ifu2bpu_data[27:26]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_l  (
    .a({i_ribm_rdata0[28],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({i_ribm_rdata0[29],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({i_ribm_rdata0[30],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({i_ribm_rdata0[31],1'b0}),
    .e({open_n1083,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_we ),
    .f(ifu2bpu_data[29:28]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c15_we ),
    .f(ifu2bpu_data[31:30]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_l  (
    .a({ifu_iaddr[4],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({ifu_iaddr[5],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({ifu_iaddr[6],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({ifu_iaddr[7],1'b0}),
    .e({open_n1118,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_we ),
    .f(ifu2bpu_iaddr[5:4]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c1_we ),
    .f(ifu2bpu_iaddr[7:6]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_l  (
    .a({ifu_iaddr[8],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({ifu_iaddr[9],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({ifu_iaddr[10],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({ifu_iaddr[11],1'b0}),
    .e({open_n1153,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_we ),
    .f(ifu2bpu_iaddr[9:8]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c2_we ),
    .f(ifu2bpu_iaddr[11:10]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_l  (
    .a({ifu_iaddr[12],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({ifu_iaddr[13],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({ifu_iaddr[14],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({ifu_iaddr[15],1'b0}),
    .e({open_n1188,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_we ),
    .f(ifu2bpu_iaddr[13:12]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c3_we ),
    .f(ifu2bpu_iaddr[15:14]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_l  (
    .a({ifu_iaddr[16],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({ifu_iaddr[17],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({ifu_iaddr[18],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({ifu_iaddr[19],1'b0}),
    .e({open_n1223,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_we ),
    .f(ifu2bpu_iaddr[17:16]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c4_we ),
    .f(ifu2bpu_iaddr[19:18]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_l  (
    .a({ifu_iaddr[20],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({ifu_iaddr[21],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({ifu_iaddr[22],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({ifu_iaddr[23],1'b0}),
    .e({open_n1258,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_we ),
    .f(ifu2bpu_iaddr[21:20]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c5_we ),
    .f(ifu2bpu_iaddr[23:22]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_l  (
    .a({ifu_iaddr[24],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({ifu_iaddr[25],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({ifu_iaddr[26],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({ifu_iaddr[27],1'b0}),
    .e({open_n1293,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_we ),
    .f(ifu2bpu_iaddr[25:24]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c6_we ),
    .f(ifu2bpu_iaddr[27:26]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_l  (
    .a({ifu_iaddr[28],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({ifu_iaddr[29],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({ifu_iaddr[30],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({ifu_iaddr[31],1'b0}),
    .e({open_n1328,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_we ),
    .f(ifu2bpu_iaddr[29:28]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c7_we ),
    .f(ifu2bpu_iaddr[31:30]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_l  (
    .a({i_ribm_rdata0[0],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({i_ribm_rdata0[1],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({i_ribm_rdata0[2],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({i_ribm_rdata0[3],1'b0}),
    .e({open_n1363,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_we ),
    .f(ifu2bpu_data[1:0]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c8_we ),
    .f(ifu2bpu_data[3:2]));
  EG_PHY_LSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_m0"),
    //.R_POSITION("X0Y0Z2"),
    .MODE("RAMW"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_l  (
    .a({i_ribm_rdata0[4],\u_IFU2BPU/u_SYNC_FIFO/hptr [0]}),
    .b({i_ribm_rdata0[5],\u_IFU2BPU/u_SYNC_FIFO/hptr [1]}),
    .c({i_ribm_rdata0[6],\u_IFU2BPU/u_SYNC_FIFO/hptr [2]}),
    .clk(i_clk),
    .d({i_ribm_rdata0[7],1'b0}),
    .e({open_n1398,\u_IFU2BPU/u_SYNC_FIFO/n19 }),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_di ),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_we ));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_m0"),
    //.R_POSITION("X0Y0Z0"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_m0  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_di [1:0]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_we ),
    .f(ifu2bpu_data[5:4]));
  EG_PHY_MSLICE #(
    //.MACRO("u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_m0"),
    //.R_POSITION("X0Y0Z1"),
    .MODE("DPRAM"))
    \u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_m1  (
    .a({\u_IFU2BPU/u_SYNC_FIFO/eptr [0],\u_IFU2BPU/u_SYNC_FIFO/eptr [0]}),
    .b({\u_IFU2BPU/u_SYNC_FIFO/eptr [1],\u_IFU2BPU/u_SYNC_FIFO/eptr [1]}),
    .c({\u_IFU2BPU/u_SYNC_FIFO/eptr [2],\u_IFU2BPU/u_SYNC_FIFO/eptr [2]}),
    .d(2'b00),
    .dpram_di(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_di [3:2]),
    .dpram_mode(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_mode ),
    .dpram_waddr(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_waddr ),
    .dpram_wclk(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_wclk ),
    .dpram_we(\u_IFU2BPU/u_SYNC_FIFO/al_ram_fifo_units_c9_we ),
    .f(ifu2bpu_data[7:6]));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU2BPU/u_SYNC_FIFO/reg0_b0  (
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n23 [0]),
    .sr(i_rstn),
    .q(\u_IFU2BPU/u_SYNC_FIFO/eptr [0]));  // ../RTL/core/fifos.v(48)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU2BPU/u_SYNC_FIFO/reg0_b1  (
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n23 [1]),
    .sr(i_rstn),
    .q(\u_IFU2BPU/u_SYNC_FIFO/eptr [1]));  // ../RTL/core/fifos.v(48)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU2BPU/u_SYNC_FIFO/reg0_b2  (
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n23 [2]),
    .sr(i_rstn),
    .q(\u_IFU2BPU/u_SYNC_FIFO/eptr [2]));  // ../RTL/core/fifos.v(48)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU2BPU/u_SYNC_FIFO/reg1_b0  (
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n24 [0]),
    .sr(i_rstn),
    .q(\u_IFU2BPU/fifo_cnt [0]));  // ../RTL/core/fifos.v(48)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU2BPU/u_SYNC_FIFO/reg1_b1  (
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n24 [1]),
    .sr(i_rstn),
    .q(\u_IFU2BPU/fifo_cnt [1]));  // ../RTL/core/fifos.v(48)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU2BPU/u_SYNC_FIFO/reg1_b2  (
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n24 [2]),
    .sr(i_rstn),
    .q(\u_IFU2BPU/fifo_cnt [2]));  // ../RTL/core/fifos.v(48)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU2BPU/u_SYNC_FIFO/reg1_b3  (
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n24 [3]),
    .sr(i_rstn),
    .q(\u_IFU2BPU/fifo_cnt [3]));  // ../RTL/core/fifos.v(48)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU2BPU/u_SYNC_FIFO/reg2_b0  (
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n22 [0]),
    .sr(i_rstn),
    .q(\u_IFU2BPU/u_SYNC_FIFO/hptr [0]));  // ../RTL/core/fifos.v(48)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU2BPU/u_SYNC_FIFO/reg2_b1  (
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n22 [1]),
    .sr(i_rstn),
    .q(\u_IFU2BPU/u_SYNC_FIFO/hptr [1]));  // ../RTL/core/fifos.v(48)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_IFU2BPU/u_SYNC_FIFO/reg2_b2  (
    .clk(i_clk),
    .d(\u_IFU2BPU/u_SYNC_FIFO/n22 [2]),
    .sr(i_rstn),
    .q(\u_IFU2BPU/u_SYNC_FIFO/hptr [2]));  // ../RTL/core/fifos.v(48)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/o_exu_taken_reg  (
    .clk(i_clk),
    .d(\u_WB/n37 ),
    .sr(i_rstn),
    .q(exu_taken_gen));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/rdwen0_reg  (
    .ce(\u_WB/n1 ),
    .clk(i_clk),
    .d(\u_WB/n2 ),
    .sr(i_rstn),
    .q(\u_WB/rdwen0 ));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/rdwen1_reg  (
    .clk(i_clk),
    .d(\u_WB/n15 ),
    .sr(i_rstn),
    .q(\u_WB/rdwen1 ));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/rdwen2_reg  (
    .clk(i_clk),
    .d(\u_WB/n16 ),
    .sr(i_rstn),
    .q(\u_WB/rdwen2 ));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg0_b0  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx0[0]),
    .q(\u_WB/rdidx0 [0]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg0_b1  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx0[1]),
    .q(\u_WB/rdidx0 [1]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg0_b2  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx0[2]),
    .q(\u_WB/rdidx0 [2]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg0_b3  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx0[3]),
    .q(\u_WB/rdidx0 [3]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg0_b4  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx0[4]),
    .q(\u_WB/rdidx0 [4]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg1_b0  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx1[0]),
    .q(\u_WB/rdidx1 [0]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg1_b1  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx1[1]),
    .q(\u_WB/rdidx1 [1]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg1_b2  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx1[2]),
    .q(\u_WB/rdidx1 [2]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg1_b3  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx1[3]),
    .q(\u_WB/rdidx1 [3]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg1_b4  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx1[4]),
    .q(\u_WB/rdidx1 [4]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg2_b0  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx2[0]),
    .q(\u_WB/rdidx2 [0]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg2_b1  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx2[1]),
    .q(\u_WB/rdidx2 [1]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg2_b2  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx2[2]),
    .q(\u_WB/rdidx2 [2]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg2_b3  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx2[3]),
    .q(\u_WB/rdidx2 [3]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg2_b4  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdidx2[4]),
    .q(\u_WB/rdidx2 [4]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b0  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[0]),
    .q(\u_WB/rdwdata0 [0]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b1  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[1]),
    .q(\u_WB/rdwdata0 [1]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b10  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[10]),
    .q(\u_WB/rdwdata0 [10]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b11  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[11]),
    .q(\u_WB/rdwdata0 [11]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b12  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[12]),
    .q(\u_WB/rdwdata0 [12]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b13  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[13]),
    .q(\u_WB/rdwdata0 [13]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b14  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[14]),
    .q(\u_WB/rdwdata0 [14]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b15  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[15]),
    .q(\u_WB/rdwdata0 [15]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b16  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[16]),
    .q(\u_WB/rdwdata0 [16]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b17  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[17]),
    .q(\u_WB/rdwdata0 [17]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b18  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[18]),
    .q(\u_WB/rdwdata0 [18]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b19  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[19]),
    .q(\u_WB/rdwdata0 [19]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b2  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[2]),
    .q(\u_WB/rdwdata0 [2]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b20  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[20]),
    .q(\u_WB/rdwdata0 [20]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b21  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[21]),
    .q(\u_WB/rdwdata0 [21]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b22  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[22]),
    .q(\u_WB/rdwdata0 [22]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b23  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[23]),
    .q(\u_WB/rdwdata0 [23]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b24  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[24]),
    .q(\u_WB/rdwdata0 [24]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b25  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[25]),
    .q(\u_WB/rdwdata0 [25]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b26  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[26]),
    .q(\u_WB/rdwdata0 [26]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b27  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[27]),
    .q(\u_WB/rdwdata0 [27]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b28  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[28]),
    .q(\u_WB/rdwdata0 [28]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b29  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[29]),
    .q(\u_WB/rdwdata0 [29]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b3  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[3]),
    .q(\u_WB/rdwdata0 [3]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b30  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[30]),
    .q(\u_WB/rdwdata0 [30]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b31  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[31]),
    .q(\u_WB/rdwdata0 [31]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b4  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[4]),
    .q(\u_WB/rdwdata0 [4]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b5  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[5]),
    .q(\u_WB/rdwdata0 [5]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b6  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[6]),
    .q(\u_WB/rdwdata0 [6]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b7  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[7]),
    .q(\u_WB/rdwdata0 [7]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b8  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[8]),
    .q(\u_WB/rdwdata0 [8]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg3_b9  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata0[9]),
    .q(\u_WB/rdwdata0 [9]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b0  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[0]),
    .q(\u_WB/rdwdata1 [0]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b1  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[1]),
    .q(\u_WB/rdwdata1 [1]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b10  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[10]),
    .q(\u_WB/rdwdata1 [10]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b11  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[11]),
    .q(\u_WB/rdwdata1 [11]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b12  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[12]),
    .q(\u_WB/rdwdata1 [12]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b13  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[13]),
    .q(\u_WB/rdwdata1 [13]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b14  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[14]),
    .q(\u_WB/rdwdata1 [14]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b15  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[15]),
    .q(\u_WB/rdwdata1 [15]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b16  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[16]),
    .q(\u_WB/rdwdata1 [16]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b17  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[17]),
    .q(\u_WB/rdwdata1 [17]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b18  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[18]),
    .q(\u_WB/rdwdata1 [18]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b19  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[19]),
    .q(\u_WB/rdwdata1 [19]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b2  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[2]),
    .q(\u_WB/rdwdata1 [2]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b20  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[20]),
    .q(\u_WB/rdwdata1 [20]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b21  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[21]),
    .q(\u_WB/rdwdata1 [21]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b22  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[22]),
    .q(\u_WB/rdwdata1 [22]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b23  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[23]),
    .q(\u_WB/rdwdata1 [23]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b24  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[24]),
    .q(\u_WB/rdwdata1 [24]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b25  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[25]),
    .q(\u_WB/rdwdata1 [25]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b26  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[26]),
    .q(\u_WB/rdwdata1 [26]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b27  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[27]),
    .q(\u_WB/rdwdata1 [27]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b28  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[28]),
    .q(\u_WB/rdwdata1 [28]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b29  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[29]),
    .q(\u_WB/rdwdata1 [29]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b3  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[3]),
    .q(\u_WB/rdwdata1 [3]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b30  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[30]),
    .q(\u_WB/rdwdata1 [30]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b31  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[31]),
    .q(\u_WB/rdwdata1 [31]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b4  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[4]),
    .q(\u_WB/rdwdata1 [4]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b5  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[5]),
    .q(\u_WB/rdwdata1 [5]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b6  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[6]),
    .q(\u_WB/rdwdata1 [6]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b7  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[7]),
    .q(\u_WB/rdwdata1 [7]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b8  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[8]),
    .q(\u_WB/rdwdata1 [8]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg4_b9  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata1[9]),
    .q(\u_WB/rdwdata1 [9]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b0  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[0]),
    .q(\u_WB/rdwdata2 [0]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b1  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[1]),
    .q(\u_WB/rdwdata2 [1]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b10  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[10]),
    .q(\u_WB/rdwdata2 [10]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b11  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[11]),
    .q(\u_WB/rdwdata2 [11]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b12  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[12]),
    .q(\u_WB/rdwdata2 [12]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b13  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[13]),
    .q(\u_WB/rdwdata2 [13]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b14  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[14]),
    .q(\u_WB/rdwdata2 [14]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b15  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[15]),
    .q(\u_WB/rdwdata2 [15]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b16  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[16]),
    .q(\u_WB/rdwdata2 [16]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b17  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[17]),
    .q(\u_WB/rdwdata2 [17]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b18  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[18]),
    .q(\u_WB/rdwdata2 [18]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b19  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[19]),
    .q(\u_WB/rdwdata2 [19]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b2  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[2]),
    .q(\u_WB/rdwdata2 [2]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b20  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[20]),
    .q(\u_WB/rdwdata2 [20]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b21  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[21]),
    .q(\u_WB/rdwdata2 [21]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b22  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[22]),
    .q(\u_WB/rdwdata2 [22]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b23  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[23]),
    .q(\u_WB/rdwdata2 [23]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b24  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[24]),
    .q(\u_WB/rdwdata2 [24]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b25  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[25]),
    .q(\u_WB/rdwdata2 [25]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b26  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[26]),
    .q(\u_WB/rdwdata2 [26]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b27  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[27]),
    .q(\u_WB/rdwdata2 [27]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b28  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[28]),
    .q(\u_WB/rdwdata2 [28]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b29  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[29]),
    .q(\u_WB/rdwdata2 [29]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b3  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[3]),
    .q(\u_WB/rdwdata2 [3]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b30  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[30]),
    .q(\u_WB/rdwdata2 [30]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b31  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[31]),
    .q(\u_WB/rdwdata2 [31]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b4  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[4]),
    .q(\u_WB/rdwdata2 [4]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b5  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[5]),
    .q(\u_WB/rdwdata2 [5]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b6  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[6]),
    .q(\u_WB/rdwdata2 [6]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b7  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[7]),
    .q(\u_WB/rdwdata2 [7]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b8  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[8]),
    .q(\u_WB/rdwdata2 [8]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_WB/reg5_b9  (
    .ce(\u_WB/mux10_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(exu_rdwdata2[9]),
    .q(\u_WB/rdwdata2 [9]));  // ../RTL/core/wb.v(57)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b0  (
    .clk(i_clk),
    .d(exu_jaddr[0]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[0]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b1  (
    .clk(i_clk),
    .d(exu_jaddr[1]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[1]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b10  (
    .clk(i_clk),
    .d(exu_jaddr[10]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[10]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b11  (
    .clk(i_clk),
    .d(exu_jaddr[11]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[11]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b12  (
    .clk(i_clk),
    .d(exu_jaddr[12]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[12]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b13  (
    .clk(i_clk),
    .d(exu_jaddr[13]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[13]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b14  (
    .clk(i_clk),
    .d(exu_jaddr[14]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[14]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b15  (
    .clk(i_clk),
    .d(exu_jaddr[15]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[15]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b16  (
    .clk(i_clk),
    .d(exu_jaddr[16]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[16]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b17  (
    .clk(i_clk),
    .d(exu_jaddr[17]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[17]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b18  (
    .clk(i_clk),
    .d(exu_jaddr[18]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[18]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b19  (
    .clk(i_clk),
    .d(exu_jaddr[19]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[19]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b2  (
    .clk(i_clk),
    .d(exu_jaddr[2]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[2]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b20  (
    .clk(i_clk),
    .d(exu_jaddr[20]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[20]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b21  (
    .clk(i_clk),
    .d(exu_jaddr[21]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[21]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b22  (
    .clk(i_clk),
    .d(exu_jaddr[22]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[22]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b23  (
    .clk(i_clk),
    .d(exu_jaddr[23]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[23]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b24  (
    .clk(i_clk),
    .d(exu_jaddr[24]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[24]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b25  (
    .clk(i_clk),
    .d(exu_jaddr[25]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[25]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b26  (
    .clk(i_clk),
    .d(exu_jaddr[26]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[26]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b27  (
    .clk(i_clk),
    .d(exu_jaddr[27]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[27]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b28  (
    .clk(i_clk),
    .d(exu_jaddr[28]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[28]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b29  (
    .clk(i_clk),
    .d(exu_jaddr[29]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[29]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b3  (
    .clk(i_clk),
    .d(exu_jaddr[3]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[3]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b30  (
    .clk(i_clk),
    .d(exu_jaddr[30]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[30]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b31  (
    .clk(i_clk),
    .d(exu_jaddr[31]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[31]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b4  (
    .clk(i_clk),
    .d(exu_jaddr[4]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[4]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b5  (
    .clk(i_clk),
    .d(exu_jaddr[5]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[5]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b6  (
    .clk(i_clk),
    .d(exu_jaddr[6]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[6]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b7  (
    .clk(i_clk),
    .d(exu_jaddr[7]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[7]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b8  (
    .clk(i_clk),
    .d(exu_jaddr[8]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[8]));  // ../RTL/core/wb.v(94)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_WB/reg6_b9  (
    .clk(i_clk),
    .d(exu_jaddr[9]),
    .sr(i_rstn),
    .q(exu_jaddr_gen[9]));  // ../RTL/core/wb.v(94)

endmodule 

module BPU  // ../RTL/core/bpu.v(14)
  (
  i_clk,
  i_data,
  i_data_vld,
  i_flush,
  i_iaddr,
  i_rd_wdata,
  i_rdidx,
  i_rdwen,
  i_rstn,
  i_stop,
  o_bpu_jaddr,
  o_bpu_rs1idx,
  o_bpu_rs1ren,
  o_bpu_rs2idx,
  o_bpu_rs2ren,
  o_bpu_taken,
  o_csr_ren,
  o_csr_zimm,
  o_csridx,
  o_decinfo,
  o_decinfo_grp,
  o_exu_op1,
  o_exu_op2,
  o_iaddr,
  o_imm,
  o_inst_vld,
  o_rdidx,
  o_rdwen,
  o_rs2rdata
  );

  input i_clk;  // ../RTL/core/bpu.v(15)
  input [31:0] i_data;  // ../RTL/core/bpu.v(24)
  input i_data_vld;  // ../RTL/core/bpu.v(22)
  input i_flush;  // ../RTL/core/bpu.v(19)
  input [31:0] i_iaddr;  // ../RTL/core/bpu.v(23)
  input [31:0] i_rd_wdata;  // ../RTL/core/bpu.v(35)
  input [4:0] i_rdidx;  // ../RTL/core/bpu.v(34)
  input i_rdwen;  // ../RTL/core/bpu.v(33)
  input i_rstn;  // ../RTL/core/bpu.v(16)
  input i_stop;  // ../RTL/core/bpu.v(18)
  output [31:0] o_bpu_jaddr;  // ../RTL/core/bpu.v(39)
  output [4:0] o_bpu_rs1idx;  // ../RTL/core/bpu.v(28)
  output o_bpu_rs1ren;  // ../RTL/core/bpu.v(27)
  output [4:0] o_bpu_rs2idx;  // ../RTL/core/bpu.v(30)
  output o_bpu_rs2ren;  // ../RTL/core/bpu.v(29)
  output o_bpu_taken;  // ../RTL/core/bpu.v(38)
  output o_csr_ren;  // ../RTL/core/bpu.v(50)
  output [31:0] o_csr_zimm;  // ../RTL/core/bpu.v(52)
  output [11:0] o_csridx;  // ../RTL/core/bpu.v(51)
  output [9:0] o_decinfo;  // ../RTL/core/bpu.v(55)
  output [5:0] o_decinfo_grp;  // ../RTL/core/bpu.v(54)
  output [31:0] o_exu_op1;  // ../RTL/core/bpu.v(43)
  output [31:0] o_exu_op2;  // ../RTL/core/bpu.v(44)
  output [31:0] o_iaddr;  // ../RTL/core/bpu.v(56)
  output [31:0] o_imm;  // ../RTL/core/bpu.v(46)
  output o_inst_vld;  // ../RTL/core/bpu.v(42)
  output [4:0] o_rdidx;  // ../RTL/core/bpu.v(48)
  output o_rdwen;  // ../RTL/core/bpu.v(47)
  output [31:0] o_rs2rdata;  // ../RTL/core/bpu.v(45)

  wire [31:0] bp_imm;  // ../RTL/core/bpu.v(105)
  wire [31:0] rs1_rdata;  // ../RTL/core/bpu.v(109)
  wire [31:0] \u_BPU_BP/n2 ;
  wire [31:0] \u_BPU_BP/n4 ;
  wire [9:0] \u_DECODE/aluinfo ;  // ../RTL/core/decode.v(261)
  wire [9:0] \u_DECODE/bjuinfo ;  // ../RTL/core/decode.v(287)
  wire [9:0] \u_DECODE/lsuinfo ;  // ../RTL/core/decode.v(278)
  wire [31:0] \u_DECODE/n23 ;
  wire [31:0] \u_DECODE/n4 ;
  wire [31:0] \u_DECODE/n5 ;
  wire [31:0] \u_DECODE/n57 ;
  wire [9:0] \u_DECODE/n67 ;
  wire [31:0] \u_DECODE/n7 ;
  wire [9:0] \u_DECODE/n71 ;
  wire _al_u103_o;
  wire _al_u109_o;
  wire _al_u112_o;
  wire _al_u124_o;
  wire _al_u129_o;
  wire _al_u156_o;
  wire _al_u158_o;
  wire _al_u172_o;
  wire _al_u193_o;
  wire _al_u195_o;
  wire _al_u197_o;
  wire _al_u199_o;
  wire _al_u200_o;
  wire _al_u201_o;
  wire _al_u216_o;
  wire _al_u236_o;
  wire _al_u237_o;
  wire _al_u260_o;
  wire _al_u262_o;
  wire _al_u264_o;
  wire _al_u265_o;
  wire _al_u266_o;
  wire _al_u268_o;
  wire _al_u26_o;
  wire _al_u271_o;
  wire _al_u276_o;
  wire _al_u277_o;
  wire _al_u279_o;
  wire _al_u27_o;
  wire _al_u63_o;
  wire _al_u65_o;
  wire _al_u66_o;
  wire _al_u95_o;
  wire _al_u99_o;
  wire inst_jalr_lutinv;  // ../RTL/core/bpu.v(102)
  wire jalr_rs1ren;  // ../RTL/core/bpu.v(162)
  wire rs1ren;  // ../RTL/core/bpu.v(107)
  wire rs1topc_lutinv;  // ../RTL/core/bpu.v(114)
  wire rs2ren;  // ../RTL/core/bpu.v(110)
  wire \u_BPU_BP/add0/c11 ;  // ../RTL/core/bpu_bp.v(44)
  wire \u_BPU_BP/add0/c15 ;  // ../RTL/core/bpu_bp.v(44)
  wire \u_BPU_BP/add0/c19 ;  // ../RTL/core/bpu_bp.v(44)
  wire \u_BPU_BP/add0/c23 ;  // ../RTL/core/bpu_bp.v(44)
  wire \u_BPU_BP/add0/c27 ;  // ../RTL/core/bpu_bp.v(44)
  wire \u_BPU_BP/add0/c3 ;  // ../RTL/core/bpu_bp.v(44)
  wire \u_BPU_BP/add0/c31 ;  // ../RTL/core/bpu_bp.v(44)
  wire \u_BPU_BP/add0/c7 ;  // ../RTL/core/bpu_bp.v(44)
  wire \u_BPU_BP/add1/c1 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c11 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c13 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c15 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c17 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c19 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c21 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c23 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c25 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c27 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c29 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c3 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c31 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c5 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c7 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_BPU_BP/add1/c9 ;  // ../RTL/core/bpu_bp.v(45)
  wire \u_DECODE/func7_0000000_lutinv ;  // ../RTL/core/decode.v(107)
  wire \u_DECODE/func7_0000001_lutinv ;  // ../RTL/core/decode.v(109)
  wire \u_DECODE/func7_0100000_lutinv ;  // ../RTL/core/decode.v(108)
  wire \u_DECODE/func_000_lutinv ;  // ../RTL/core/decode.v(97)
  wire \u_DECODE/func_001_lutinv ;  // ../RTL/core/decode.v(98)
  wire \u_DECODE/func_010_lutinv ;  // ../RTL/core/decode.v(99)
  wire \u_DECODE/func_011_lutinv ;  // ../RTL/core/decode.v(100)
  wire \u_DECODE/func_111_lutinv ;  // ../RTL/core/decode.v(104)
  wire \u_DECODE/inst_ebreak ;  // ../RTL/core/decode.v(165)
  wire \u_DECODE/n1_lutinv ;
  wire \u_DECODE/n21_lutinv ;
  wire \u_DECODE/n38_lutinv ;
  wire \u_DECODE/n3_lutinv ;
  wire \u_DECODE/n42_lutinv ;
  wire \u_DECODE/n47_lutinv ;
  wire \u_DECODE/n48_lutinv ;
  wire \u_DECODE/opc_op_lutinv ;  // ../RTL/core/decode.v(92)
  wire \u_DECODE/opc_opimm_lutinv ;  // ../RTL/core/decode.v(91)
  wire \u_DECODE/opc_rv32 ;  // ../RTL/core/decode.v(67)

  assign o_iaddr[31] = i_iaddr[31];
  assign o_iaddr[30] = i_iaddr[30];
  assign o_iaddr[29] = i_iaddr[29];
  assign o_iaddr[28] = i_iaddr[28];
  assign o_iaddr[27] = i_iaddr[27];
  assign o_iaddr[26] = i_iaddr[26];
  assign o_iaddr[25] = i_iaddr[25];
  assign o_iaddr[24] = i_iaddr[24];
  assign o_iaddr[23] = i_iaddr[23];
  assign o_iaddr[22] = i_iaddr[22];
  assign o_iaddr[21] = i_iaddr[21];
  assign o_iaddr[20] = i_iaddr[20];
  assign o_iaddr[19] = i_iaddr[19];
  assign o_iaddr[18] = i_iaddr[18];
  assign o_iaddr[17] = i_iaddr[17];
  assign o_iaddr[16] = i_iaddr[16];
  assign o_iaddr[15] = i_iaddr[15];
  assign o_iaddr[14] = i_iaddr[14];
  assign o_iaddr[13] = i_iaddr[13];
  assign o_iaddr[12] = i_iaddr[12];
  assign o_iaddr[11] = i_iaddr[11];
  assign o_iaddr[10] = i_iaddr[10];
  assign o_iaddr[9] = i_iaddr[9];
  assign o_iaddr[8] = i_iaddr[8];
  assign o_iaddr[7] = i_iaddr[7];
  assign o_iaddr[6] = i_iaddr[6];
  assign o_iaddr[5] = i_iaddr[5];
  assign o_iaddr[4] = i_iaddr[4];
  assign o_iaddr[3] = i_iaddr[3];
  assign o_iaddr[2] = i_iaddr[2];
  assign o_iaddr[1] = i_iaddr[1];
  assign o_iaddr[0] = i_iaddr[0];
  assign o_bpu_rs1idx[4] = i_data[19];
  assign o_bpu_rs1idx[3] = i_data[18];
  assign o_bpu_rs1idx[2] = i_data[17];
  assign o_bpu_rs1idx[1] = i_data[16];
  assign o_bpu_rs1idx[0] = i_data[15];
  assign o_bpu_rs2idx[4] = i_data[24];
  assign o_bpu_rs2idx[3] = i_data[23];
  assign o_bpu_rs2idx[2] = i_data[22];
  assign o_bpu_rs2idx[1] = i_data[21];
  assign o_bpu_rs2idx[0] = i_data[20];
  assign o_csr_ren = \u_DECODE/n57 [0];
  assign o_csr_zimm[31] = 1'b0;
  assign o_csr_zimm[30] = 1'b0;
  assign o_csr_zimm[29] = 1'b0;
  assign o_csr_zimm[28] = 1'b0;
  assign o_csr_zimm[27] = 1'b0;
  assign o_csr_zimm[26] = 1'b0;
  assign o_csr_zimm[25] = 1'b0;
  assign o_csr_zimm[24] = 1'b0;
  assign o_csr_zimm[23] = 1'b0;
  assign o_csr_zimm[22] = 1'b0;
  assign o_csr_zimm[21] = 1'b0;
  assign o_csr_zimm[20] = 1'b0;
  assign o_csr_zimm[19] = 1'b0;
  assign o_csr_zimm[18] = 1'b0;
  assign o_csr_zimm[17] = 1'b0;
  assign o_csr_zimm[16] = 1'b0;
  assign o_csr_zimm[15] = 1'b0;
  assign o_csr_zimm[14] = 1'b0;
  assign o_csr_zimm[13] = 1'b0;
  assign o_csr_zimm[12] = 1'b0;
  assign o_csr_zimm[11] = 1'b0;
  assign o_csr_zimm[10] = 1'b0;
  assign o_csr_zimm[9] = 1'b0;
  assign o_csr_zimm[8] = 1'b0;
  assign o_csr_zimm[7] = 1'b0;
  assign o_csr_zimm[6] = 1'b0;
  assign o_csr_zimm[5] = 1'b0;
  assign o_decinfo[9] = \u_DECODE/aluinfo [9];
  assign o_decinfo[8] = \u_DECODE/n71 [8];
  assign o_rdidx[4] = i_data[11];
  assign o_rdidx[3] = i_data[10];
  assign o_rdidx[2] = i_data[9];
  assign o_rdidx[1] = i_data[8];
  assign o_rdidx[0] = i_data[7];
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u100 (
    .a(i_data[14]),
    .b(i_data[13]),
    .c(i_data[12]),
    .o(\u_DECODE/func_011_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u101 (
    .a(_al_u99_o),
    .b(\u_DECODE/func_011_lutinv ),
    .o(\u_DECODE/aluinfo [9]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*B*~(C*A))"),
    .INIT(32'h0000004c))
    _al_u102 (
    .a(i_data[6]),
    .b(i_data[5]),
    .c(i_data[4]),
    .d(i_data[3]),
    .e(i_data[2]),
    .o(\u_DECODE/n48_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u103 (
    .a(i_data[22]),
    .b(i_data[21]),
    .c(i_data[20]),
    .o(_al_u103_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*B))"),
    .INIT(16'haaa2))
    _al_u104 (
    .a(\u_DECODE/n48_lutinv ),
    .b(_al_u103_o),
    .c(i_data[24]),
    .d(i_data[23]),
    .o(rs2ren));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    _al_u105 (
    .a(i_data[6]),
    .b(i_data[5]),
    .c(i_data[4]),
    .d(i_data[3]),
    .e(i_data[2]),
    .o(\u_DECODE/n3_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u106 (
    .a(i_data_vld),
    .b(\u_DECODE/n3_lutinv ),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[31]),
    .o(\u_DECODE/n7 [31]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(D*C*B))"),
    .INIT(16'heaaa))
    _al_u107 (
    .a(\u_DECODE/n7 [31]),
    .b(i_data_vld),
    .c(\u_DECODE/bjuinfo [1]),
    .d(\u_DECODE/opc_rv32 ),
    .o(o_bpu_taken));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~C*~(B*~A))"),
    .INIT(16'hfff4))
    _al_u108 (
    .a(\u_DECODE/func7_0000001_lutinv ),
    .b(\u_DECODE/opc_op_lutinv ),
    .c(\u_DECODE/opc_opimm_lutinv ),
    .d(\u_DECODE/n21_lutinv ),
    .o(o_decinfo_grp[0]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(~D*A)))"),
    .INIT(16'hc0e0))
    _al_u109 (
    .a(\u_DECODE/n47_lutinv ),
    .b(_al_u95_o),
    .c(i_data[31]),
    .d(i_data[6]),
    .o(_al_u109_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u110 (
    .a(\u_DECODE/n3_lutinv ),
    .b(i_data[7]),
    .o(\u_DECODE/n23 [11]));
  AL_MAP_LUT2 #(
    .EQN("~(~B*~A)"),
    .INIT(4'he))
    _al_u111 (
    .a(_al_u109_o),
    .b(\u_DECODE/n23 [11]),
    .o(o_imm[11]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u112 (
    .a(\u_DECODE/n47_lutinv ),
    .b(_al_u95_o),
    .o(_al_u112_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u113 (
    .a(_al_u112_o),
    .b(i_data[29]),
    .o(o_imm[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u114 (
    .a(_al_u112_o),
    .b(i_data[28]),
    .o(o_imm[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u115 (
    .a(_al_u112_o),
    .b(i_data[27]),
    .o(o_imm[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u116 (
    .a(_al_u112_o),
    .b(i_data[26]),
    .o(o_imm[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u117 (
    .a(_al_u112_o),
    .b(i_data[25]),
    .o(o_imm[5]));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u118 (
    .a(\u_DECODE/n47_lutinv ),
    .b(_al_u95_o),
    .c(i_data[24]),
    .d(i_data[11]),
    .o(o_imm[4]));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u119 (
    .a(\u_DECODE/n47_lutinv ),
    .b(_al_u95_o),
    .c(i_data[23]),
    .d(i_data[10]),
    .o(o_imm[3]));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u120 (
    .a(\u_DECODE/n47_lutinv ),
    .b(_al_u95_o),
    .c(i_data[22]),
    .d(i_data[9]),
    .o(o_imm[2]));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u121 (
    .a(\u_DECODE/n47_lutinv ),
    .b(_al_u95_o),
    .c(i_data[21]),
    .d(i_data[8]),
    .o(o_imm[1]));
  AL_MAP_LUT5 #(
    .EQN("(B*A*~(~E*~D*C))"),
    .INIT(32'h88888808))
    _al_u122 (
    .a(i_data_vld),
    .b(\u_DECODE/n48_lutinv ),
    .c(_al_u103_o),
    .d(i_data[24]),
    .e(i_data[23]),
    .o(o_bpu_rs2ren));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u123 (
    .a(i_data_vld),
    .b(\u_DECODE/bjuinfo [1]),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[3]),
    .o(inst_jalr_lutinv));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    _al_u124 (
    .a(i_data[19]),
    .b(i_data[18]),
    .c(i_data[17]),
    .d(i_data[16]),
    .e(i_data[15]),
    .o(_al_u124_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u125 (
    .a(inst_jalr_lutinv),
    .b(_al_u124_o),
    .o(jalr_rs1ren));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u126 (
    .a(\u_BPU_BP/n2 [0]),
    .b(\u_BPU_BP/n4 [0]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[20]),
    .o(o_bpu_jaddr[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u127 (
    .a(i_data_vld),
    .b(o_decinfo_grp[2]),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[31]),
    .o(bp_imm[31]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u128 (
    .a(i_data[6]),
    .b(i_data[5]),
    .c(i_data[4]),
    .d(i_data[3]),
    .o(\u_DECODE/n38_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u129 (
    .a(i_data_vld),
    .b(\u_DECODE/n38_lutinv ),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[31]),
    .o(_al_u129_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u130 (
    .a(_al_u27_o),
    .b(i_data[4]),
    .c(i_data[3]),
    .d(i_data[2]),
    .o(\u_DECODE/n1_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    _al_u131 (
    .a(_al_u129_o),
    .b(i_data_vld),
    .c(\u_DECODE/n1_lutinv ),
    .d(\u_DECODE/opc_rv32 ),
    .e(i_data[19]),
    .o(bp_imm[19]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    _al_u132 (
    .a(_al_u129_o),
    .b(i_data_vld),
    .c(\u_DECODE/n1_lutinv ),
    .d(\u_DECODE/opc_rv32 ),
    .e(i_data[18]),
    .o(bp_imm[18]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    _al_u133 (
    .a(_al_u129_o),
    .b(i_data_vld),
    .c(\u_DECODE/n1_lutinv ),
    .d(\u_DECODE/opc_rv32 ),
    .e(i_data[17]),
    .o(bp_imm[17]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    _al_u134 (
    .a(_al_u129_o),
    .b(i_data_vld),
    .c(\u_DECODE/n1_lutinv ),
    .d(\u_DECODE/opc_rv32 ),
    .e(i_data[16]),
    .o(bp_imm[16]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    _al_u135 (
    .a(_al_u129_o),
    .b(i_data_vld),
    .c(\u_DECODE/n1_lutinv ),
    .d(\u_DECODE/opc_rv32 ),
    .e(i_data[15]),
    .o(bp_imm[15]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    _al_u136 (
    .a(_al_u129_o),
    .b(i_data_vld),
    .c(\u_DECODE/n1_lutinv ),
    .d(\u_DECODE/opc_rv32 ),
    .e(i_data[14]),
    .o(bp_imm[14]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    _al_u137 (
    .a(_al_u129_o),
    .b(i_data_vld),
    .c(\u_DECODE/n1_lutinv ),
    .d(\u_DECODE/opc_rv32 ),
    .e(i_data[13]),
    .o(bp_imm[13]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    _al_u138 (
    .a(_al_u129_o),
    .b(i_data_vld),
    .c(\u_DECODE/n1_lutinv ),
    .d(\u_DECODE/opc_rv32 ),
    .e(i_data[12]),
    .o(bp_imm[12]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u139 (
    .a(i_data_vld),
    .b(\u_DECODE/n1_lutinv ),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[20]),
    .o(\u_DECODE/n4 [11]));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u140 (
    .a(i_data_vld),
    .b(\u_DECODE/n38_lutinv ),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[31]),
    .e(i_data[2]),
    .o(\u_DECODE/n5 [31]));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~A*~(E*D*C))"),
    .INIT(32'hfeeeeeee))
    _al_u141 (
    .a(\u_DECODE/n4 [11]),
    .b(\u_DECODE/n5 [31]),
    .c(\u_DECODE/n23 [11]),
    .d(i_data_vld),
    .e(\u_DECODE/opc_rv32 ),
    .o(bp_imm[11]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u142 (
    .a(i_data_vld),
    .b(o_decinfo_grp[2]),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[30]),
    .o(bp_imm[10]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u143 (
    .a(i_data_vld),
    .b(o_decinfo_grp[2]),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[29]),
    .o(bp_imm[9]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u144 (
    .a(i_data_vld),
    .b(o_decinfo_grp[2]),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[28]),
    .o(bp_imm[8]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u145 (
    .a(i_data_vld),
    .b(o_decinfo_grp[2]),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[27]),
    .o(bp_imm[7]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u146 (
    .a(i_data_vld),
    .b(o_decinfo_grp[2]),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[26]),
    .o(bp_imm[6]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u147 (
    .a(i_data_vld),
    .b(o_decinfo_grp[2]),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[25]),
    .o(bp_imm[5]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u148 (
    .a(i_data_vld),
    .b(\u_DECODE/n3_lutinv ),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[11]),
    .o(\u_DECODE/n7 [4]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    _al_u149 (
    .a(\u_DECODE/n7 [4]),
    .b(i_data_vld),
    .c(\u_DECODE/bjuinfo [1]),
    .d(\u_DECODE/opc_rv32 ),
    .e(i_data[24]),
    .o(bp_imm[4]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u150 (
    .a(i_data_vld),
    .b(\u_DECODE/n3_lutinv ),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[10]),
    .o(\u_DECODE/n7 [3]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    _al_u151 (
    .a(\u_DECODE/n7 [3]),
    .b(i_data_vld),
    .c(\u_DECODE/bjuinfo [1]),
    .d(\u_DECODE/opc_rv32 ),
    .e(i_data[23]),
    .o(bp_imm[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u152 (
    .a(i_data_vld),
    .b(\u_DECODE/n3_lutinv ),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[9]),
    .o(\u_DECODE/n7 [2]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    _al_u153 (
    .a(\u_DECODE/n7 [2]),
    .b(i_data_vld),
    .c(\u_DECODE/bjuinfo [1]),
    .d(\u_DECODE/opc_rv32 ),
    .e(i_data[22]),
    .o(bp_imm[2]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u154 (
    .a(i_data_vld),
    .b(\u_DECODE/n3_lutinv ),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[8]),
    .o(\u_DECODE/n7 [1]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~(E*D*C*B))"),
    .INIT(32'heaaaaaaa))
    _al_u155 (
    .a(\u_DECODE/n7 [1]),
    .b(i_data_vld),
    .c(\u_DECODE/bjuinfo [1]),
    .d(\u_DECODE/opc_rv32 ),
    .e(i_data[21]),
    .o(bp_imm[1]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u156 (
    .a(\u_DECODE/opc_opimm_lutinv ),
    .b(o_decinfo_grp[1]),
    .c(\u_DECODE/n21_lutinv ),
    .o(_al_u156_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    _al_u157 (
    .a(o_rs2rdata[0]),
    .b(o_imm[0]),
    .c(_al_u156_o),
    .o(o_exu_op2[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u158 (
    .a(i_data[14]),
    .b(i_data[13]),
    .o(_al_u158_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u159 (
    .a(_al_u158_o),
    .b(i_data[12]),
    .o(\u_DECODE/func_111_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u160 (
    .a(i_data[14]),
    .b(i_data[13]),
    .c(i_data[12]),
    .o(\u_DECODE/func_010_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(E*~B)*~(D*A))"),
    .INIT(32'hfbf3faf0))
    _al_u161 (
    .a(o_decinfo_grp[3]),
    .b(_al_u99_o),
    .c(\u_DECODE/n7 [31]),
    .d(\u_DECODE/func_111_lutinv ),
    .e(\u_DECODE/func_010_lutinv ),
    .o(\u_DECODE/n71 [8]));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    _al_u162 (
    .a(o_rs2rdata[11]),
    .b(_al_u109_o),
    .c(_al_u156_o),
    .o(o_exu_op2[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u163 (
    .a(o_rs2rdata[9]),
    .b(o_imm[9]),
    .c(_al_u156_o),
    .o(o_exu_op2[9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u164 (
    .a(o_rs2rdata[8]),
    .b(o_imm[8]),
    .c(_al_u156_o),
    .o(o_exu_op2[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u165 (
    .a(o_rs2rdata[7]),
    .b(o_imm[7]),
    .c(_al_u156_o),
    .o(o_exu_op2[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u166 (
    .a(o_rs2rdata[6]),
    .b(o_imm[6]),
    .c(_al_u156_o),
    .o(o_exu_op2[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u167 (
    .a(o_rs2rdata[5]),
    .b(o_imm[5]),
    .c(_al_u156_o),
    .o(o_exu_op2[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u168 (
    .a(o_rs2rdata[4]),
    .b(o_imm[4]),
    .c(_al_u156_o),
    .o(o_exu_op2[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u169 (
    .a(o_rs2rdata[3]),
    .b(o_imm[3]),
    .c(_al_u156_o),
    .o(o_exu_op2[3]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u170 (
    .a(o_rs2rdata[2]),
    .b(o_imm[2]),
    .c(_al_u156_o),
    .o(o_exu_op2[2]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u171 (
    .a(o_rs2rdata[1]),
    .b(o_imm[1]),
    .c(_al_u156_o),
    .o(o_exu_op2[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u172 (
    .a(_al_u112_o),
    .b(i_data[31]),
    .o(_al_u172_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u173 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[14]),
    .o(o_imm[14]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u174 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[13]),
    .o(o_imm[13]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u175 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[12]),
    .o(o_imm[12]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u176 (
    .a(_al_u112_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[31]),
    .o(o_imm[31]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u177 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[30]),
    .o(o_imm[30]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u178 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[29]),
    .o(o_imm[29]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u179 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[28]),
    .o(o_imm[28]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u180 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[27]),
    .o(o_imm[27]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u181 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[26]),
    .o(o_imm[26]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u182 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[25]),
    .o(o_imm[25]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u183 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[24]),
    .o(o_imm[24]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u184 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[23]),
    .o(o_imm[23]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u185 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[22]),
    .o(o_imm[22]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u186 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[21]),
    .o(o_imm[21]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u187 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[20]),
    .o(o_imm[20]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u188 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[19]),
    .o(o_imm[19]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u189 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[18]),
    .o(o_imm[18]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u190 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[17]),
    .o(o_imm[17]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u191 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[16]),
    .o(o_imm[16]));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(C*B))"),
    .INIT(8'hea))
    _al_u192 (
    .a(_al_u172_o),
    .b(\u_DECODE/n21_lutinv ),
    .c(i_data[15]),
    .o(o_imm[15]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~A*~(~E*D*B)))"),
    .INIT(32'ha0a0e0a0))
    _al_u193 (
    .a(o_decinfo_grp[4]),
    .b(\u_DECODE/n3_lutinv ),
    .c(i_data[14]),
    .d(i_data[13]),
    .e(i_data[12]),
    .o(_al_u193_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u194 (
    .a(i_data[14]),
    .b(i_data[13]),
    .o(\u_DECODE/lsuinfo [5]));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*C*A))"),
    .INIT(16'h1333))
    _al_u195 (
    .a(o_decinfo_grp[3]),
    .b(_al_u193_o),
    .c(\u_DECODE/lsuinfo [5]),
    .d(i_data[12]),
    .o(_al_u195_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*~B))"),
    .INIT(8'h75))
    _al_u196 (
    .a(_al_u195_o),
    .b(_al_u99_o),
    .c(\u_DECODE/func_111_lutinv ),
    .o(o_decinfo[6]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u197 (
    .a(i_data[31]),
    .b(i_data[30]),
    .c(i_data[29]),
    .d(i_data[28]),
    .o(_al_u197_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u198 (
    .a(_al_u197_o),
    .b(i_data[27]),
    .c(i_data[26]),
    .d(i_data[25]),
    .o(\u_DECODE/func7_0100000_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(~B*~A))"),
    .INIT(16'he000))
    _al_u199 (
    .a(\u_DECODE/func7_0000001_lutinv ),
    .b(\u_DECODE/func7_0100000_lutinv ),
    .c(\u_DECODE/opc_op_lutinv ),
    .d(\u_DECODE/func_000_lutinv ),
    .o(_al_u199_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(~D*B))"),
    .INIT(16'h0501))
    _al_u200 (
    .a(_al_u199_o),
    .b(\u_DECODE/n47_lutinv ),
    .c(\u_DECODE/bjuinfo [1]),
    .d(i_data[6]),
    .o(_al_u200_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    _al_u201 (
    .a(o_decinfo_grp[4]),
    .b(\u_DECODE/func_000_lutinv ),
    .c(i_data[25]),
    .d(i_data[24]),
    .e(i_data[23]),
    .o(_al_u201_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(D*C*B))"),
    .INIT(16'hd555))
    _al_u202 (
    .a(_al_u200_o),
    .b(_al_u201_o),
    .c(_al_u66_o),
    .d(_al_u103_o),
    .o(o_decinfo[1]));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~B*~(C*~A))"),
    .INIT(16'hffdc))
    _al_u203 (
    .a(_al_u99_o),
    .b(o_decinfo_grp[1]),
    .c(\u_DECODE/func_000_lutinv ),
    .d(\u_DECODE/n21_lutinv ),
    .o(o_decinfo_grp[5]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u204 (
    .a(\u_BPU_BP/n2 [31]),
    .b(\u_BPU_BP/n4 [31]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[31]),
    .o(o_bpu_jaddr[31]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u205 (
    .a(\u_BPU_BP/n2 [30]),
    .b(\u_BPU_BP/n4 [30]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[31]),
    .o(o_bpu_jaddr[30]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u206 (
    .a(\u_BPU_BP/n2 [29]),
    .b(\u_BPU_BP/n4 [29]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[31]),
    .o(o_bpu_jaddr[29]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u207 (
    .a(\u_BPU_BP/n2 [28]),
    .b(\u_BPU_BP/n4 [28]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[31]),
    .o(o_bpu_jaddr[28]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u208 (
    .a(\u_BPU_BP/n2 [27]),
    .b(\u_BPU_BP/n4 [27]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[31]),
    .o(o_bpu_jaddr[27]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u209 (
    .a(\u_BPU_BP/n2 [26]),
    .b(\u_BPU_BP/n4 [26]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[31]),
    .o(o_bpu_jaddr[26]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u210 (
    .a(\u_BPU_BP/n2 [25]),
    .b(\u_BPU_BP/n4 [25]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[31]),
    .o(o_bpu_jaddr[25]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u211 (
    .a(\u_BPU_BP/n2 [24]),
    .b(\u_BPU_BP/n4 [24]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[31]),
    .o(o_bpu_jaddr[24]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u212 (
    .a(\u_BPU_BP/n2 [23]),
    .b(\u_BPU_BP/n4 [23]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[31]),
    .o(o_bpu_jaddr[23]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u213 (
    .a(\u_BPU_BP/n2 [22]),
    .b(\u_BPU_BP/n4 [22]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[31]),
    .o(o_bpu_jaddr[22]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u214 (
    .a(\u_BPU_BP/n2 [21]),
    .b(\u_BPU_BP/n4 [21]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[31]),
    .o(o_bpu_jaddr[21]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafeca0ec))
    _al_u215 (
    .a(\u_BPU_BP/n2 [20]),
    .b(\u_BPU_BP/n4 [20]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[31]),
    .o(o_bpu_jaddr[20]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u216 (
    .a(jalr_rs1ren),
    .b(\u_DECODE/n5 [31]),
    .o(_al_u216_o));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(~E*B)*~(D*A))"),
    .INIT(32'hfaf0fefc))
    _al_u217 (
    .a(\u_BPU_BP/n2 [19]),
    .b(\u_BPU_BP/n4 [19]),
    .c(_al_u216_o),
    .d(jalr_rs1ren),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[19]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(~E*B)*~(D*A))"),
    .INIT(32'hfaf0fefc))
    _al_u218 (
    .a(\u_BPU_BP/n2 [18]),
    .b(\u_BPU_BP/n4 [18]),
    .c(_al_u216_o),
    .d(jalr_rs1ren),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[18]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(~E*B)*~(D*A))"),
    .INIT(32'hfaf0fefc))
    _al_u219 (
    .a(\u_BPU_BP/n2 [17]),
    .b(\u_BPU_BP/n4 [17]),
    .c(_al_u216_o),
    .d(jalr_rs1ren),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[17]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(~E*B)*~(D*A))"),
    .INIT(32'hfaf0fefc))
    _al_u220 (
    .a(\u_BPU_BP/n2 [16]),
    .b(\u_BPU_BP/n4 [16]),
    .c(_al_u216_o),
    .d(jalr_rs1ren),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[16]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(~E*B)*~(D*A))"),
    .INIT(32'hfaf0fefc))
    _al_u221 (
    .a(\u_BPU_BP/n2 [15]),
    .b(\u_BPU_BP/n4 [15]),
    .c(_al_u216_o),
    .d(jalr_rs1ren),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[15]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(~E*B)*~(D*A))"),
    .INIT(32'hfaf0fefc))
    _al_u222 (
    .a(\u_BPU_BP/n2 [14]),
    .b(\u_BPU_BP/n4 [14]),
    .c(_al_u216_o),
    .d(jalr_rs1ren),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[14]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(~E*B)*~(D*A))"),
    .INIT(32'hfaf0fefc))
    _al_u223 (
    .a(\u_BPU_BP/n2 [13]),
    .b(\u_BPU_BP/n4 [13]),
    .c(_al_u216_o),
    .d(jalr_rs1ren),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[13]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(~E*B)*~(D*A))"),
    .INIT(32'hfaf0fefc))
    _al_u224 (
    .a(\u_BPU_BP/n2 [12]),
    .b(\u_BPU_BP/n4 [12]),
    .c(_al_u216_o),
    .d(jalr_rs1ren),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[12]));
  AL_MAP_LUT5 #(
    .EQN("~(~C*~(~E*B)*~(D*A))"),
    .INIT(32'hfaf0fefc))
    _al_u225 (
    .a(\u_BPU_BP/n2 [11]),
    .b(\u_BPU_BP/n4 [11]),
    .c(_al_u216_o),
    .d(jalr_rs1ren),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[11]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haf8ca08c))
    _al_u226 (
    .a(\u_BPU_BP/n2 [10]),
    .b(\u_BPU_BP/n4 [10]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[30]),
    .o(o_bpu_jaddr[10]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haf8ca08c))
    _al_u227 (
    .a(\u_BPU_BP/n2 [9]),
    .b(\u_BPU_BP/n4 [9]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[29]),
    .o(o_bpu_jaddr[9]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haf8ca08c))
    _al_u228 (
    .a(\u_BPU_BP/n2 [8]),
    .b(\u_BPU_BP/n4 [8]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[28]),
    .o(o_bpu_jaddr[8]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haf8ca08c))
    _al_u229 (
    .a(\u_BPU_BP/n2 [7]),
    .b(\u_BPU_BP/n4 [7]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[27]),
    .o(o_bpu_jaddr[7]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haf8ca08c))
    _al_u230 (
    .a(\u_BPU_BP/n2 [6]),
    .b(\u_BPU_BP/n4 [6]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[26]),
    .o(o_bpu_jaddr[6]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haf8ca08c))
    _al_u231 (
    .a(\u_BPU_BP/n2 [5]),
    .b(\u_BPU_BP/n4 [5]),
    .c(jalr_rs1ren),
    .d(inst_jalr_lutinv),
    .e(i_data[25]),
    .o(o_bpu_jaddr[5]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*B*C*D*~(E)+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafa08c8c))
    _al_u232 (
    .a(\u_BPU_BP/n2 [4]),
    .b(\u_BPU_BP/n4 [4]),
    .c(jalr_rs1ren),
    .d(bp_imm[4]),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[4]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*B*C*D*~(E)+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafa08c8c))
    _al_u233 (
    .a(\u_BPU_BP/n2 [3]),
    .b(\u_BPU_BP/n4 [3]),
    .c(jalr_rs1ren),
    .d(bp_imm[3]),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[3]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*B*C*D*~(E)+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafa08c8c))
    _al_u234 (
    .a(\u_BPU_BP/n2 [2]),
    .b(\u_BPU_BP/n4 [2]),
    .c(jalr_rs1ren),
    .d(bp_imm[2]),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[2]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*B*C*D*~(E)+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hafa08c8c))
    _al_u235 (
    .a(\u_BPU_BP/n2 [1]),
    .b(\u_BPU_BP/n4 [1]),
    .c(jalr_rs1ren),
    .d(bp_imm[1]),
    .e(inst_jalr_lutinv),
    .o(o_bpu_jaddr[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u236 (
    .a(\u_DECODE/func7_0100000_lutinv ),
    .b(\u_DECODE/lsuinfo [5]),
    .c(i_data[12]),
    .o(_al_u236_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u237 (
    .a(_al_u236_o),
    .b(\u_DECODE/opc_opimm_lutinv ),
    .o(_al_u237_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u238 (
    .a(_al_u237_o),
    .b(o_decinfo_grp[1]),
    .c(\u_DECODE/n47_lutinv ),
    .d(i_data[30]),
    .o(o_imm[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u239 (
    .a(o_rs2rdata[14]),
    .b(o_imm[14]),
    .c(_al_u156_o),
    .o(o_exu_op2[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u240 (
    .a(o_rs2rdata[13]),
    .b(o_imm[13]),
    .c(_al_u156_o),
    .o(o_exu_op2[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u241 (
    .a(o_rs2rdata[12]),
    .b(o_imm[12]),
    .c(_al_u156_o),
    .o(o_exu_op2[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u242 (
    .a(o_rs2rdata[31]),
    .b(o_imm[31]),
    .c(_al_u156_o),
    .o(o_exu_op2[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u243 (
    .a(o_rs2rdata[30]),
    .b(o_imm[30]),
    .c(_al_u156_o),
    .o(o_exu_op2[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u244 (
    .a(o_rs2rdata[29]),
    .b(o_imm[29]),
    .c(_al_u156_o),
    .o(o_exu_op2[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u245 (
    .a(o_rs2rdata[28]),
    .b(o_imm[28]),
    .c(_al_u156_o),
    .o(o_exu_op2[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u246 (
    .a(o_rs2rdata[27]),
    .b(o_imm[27]),
    .c(_al_u156_o),
    .o(o_exu_op2[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u247 (
    .a(o_rs2rdata[26]),
    .b(o_imm[26]),
    .c(_al_u156_o),
    .o(o_exu_op2[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u248 (
    .a(o_rs2rdata[25]),
    .b(o_imm[25]),
    .c(_al_u156_o),
    .o(o_exu_op2[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u249 (
    .a(o_rs2rdata[24]),
    .b(o_imm[24]),
    .c(_al_u156_o),
    .o(o_exu_op2[24]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u25 (
    .a(i_stop),
    .b(i_data_vld),
    .o(o_inst_vld));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u250 (
    .a(o_rs2rdata[23]),
    .b(o_imm[23]),
    .c(_al_u156_o),
    .o(o_exu_op2[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u251 (
    .a(o_rs2rdata[22]),
    .b(o_imm[22]),
    .c(_al_u156_o),
    .o(o_exu_op2[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u252 (
    .a(o_rs2rdata[21]),
    .b(o_imm[21]),
    .c(_al_u156_o),
    .o(o_exu_op2[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u253 (
    .a(o_rs2rdata[20]),
    .b(o_imm[20]),
    .c(_al_u156_o),
    .o(o_exu_op2[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u254 (
    .a(o_rs2rdata[19]),
    .b(o_imm[19]),
    .c(_al_u156_o),
    .o(o_exu_op2[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u255 (
    .a(o_rs2rdata[18]),
    .b(o_imm[18]),
    .c(_al_u156_o),
    .o(o_exu_op2[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u256 (
    .a(o_rs2rdata[17]),
    .b(o_imm[17]),
    .c(_al_u156_o),
    .o(o_exu_op2[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u257 (
    .a(o_rs2rdata[16]),
    .b(o_imm[16]),
    .c(_al_u156_o),
    .o(o_exu_op2[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u258 (
    .a(o_rs2rdata[15]),
    .b(o_imm[15]),
    .c(_al_u156_o),
    .o(o_exu_op2[15]));
  AL_MAP_LUT5 #(
    .EQN("(~D*C*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E))"),
    .INIT(32'h00a000c0))
    _al_u259 (
    .a(_al_u236_o),
    .b(\u_DECODE/func_010_lutinv ),
    .c(_al_u63_o),
    .d(i_data[6]),
    .e(i_data[4]),
    .o(\u_DECODE/n67 [4]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u26 (
    .a(i_data[4]),
    .b(i_data[3]),
    .c(i_data[2]),
    .o(_al_u26_o));
  AL_MAP_LUT4 #(
    .EQN("~((C*B)*~(A)*~(D)+(C*B)*A*~(D)+~((C*B))*A*D+(C*B)*A*D)"),
    .INIT(16'h553f))
    _al_u260 (
    .a(o_decinfo_grp[4]),
    .b(\u_DECODE/n3_lutinv ),
    .c(i_data[14]),
    .d(i_data[13]),
    .o(_al_u260_o));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(~E*~C)*~(D*A))"),
    .INIT(32'heeccefcf))
    _al_u261 (
    .a(o_decinfo_grp[3]),
    .b(\u_DECODE/n67 [4]),
    .c(_al_u260_o),
    .d(\u_DECODE/func_011_lutinv ),
    .e(i_data[12]),
    .o(o_decinfo[4]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~(~B*~A))"),
    .INIT(16'h0e00))
    _al_u262 (
    .a(o_decinfo_grp[4]),
    .b(o_decinfo_grp[1]),
    .c(i_data[13]),
    .d(i_data[12]),
    .o(_al_u262_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u263 (
    .a(i_data[14]),
    .b(i_data[13]),
    .c(i_data[12]),
    .o(\u_DECODE/func_001_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u264 (
    .a(_al_u262_o),
    .b(\u_DECODE/n3_lutinv ),
    .c(\u_DECODE/func_001_lutinv ),
    .o(_al_u264_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u265 (
    .a(\u_DECODE/func7_0000000_lutinv ),
    .b(_al_u26_o),
    .c(i_data[6]),
    .o(_al_u265_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u266 (
    .a(_al_u264_o),
    .b(_al_u265_o),
    .c(\u_DECODE/lsuinfo [5]),
    .d(i_data[12]),
    .o(_al_u266_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(C*B))"),
    .INIT(8'hd5))
    _al_u267 (
    .a(_al_u266_o),
    .b(o_decinfo_grp[3]),
    .c(\u_DECODE/func_010_lutinv ),
    .o(o_decinfo[3]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u268 (
    .a(_al_u66_o),
    .b(\u_DECODE/opc_op_lutinv ),
    .c(\u_DECODE/opc_opimm_lutinv ),
    .o(_al_u268_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hf333f500))
    _al_u269 (
    .a(_al_u268_o),
    .b(_al_u260_o),
    .c(o_decinfo_grp[1]),
    .d(\u_DECODE/lsuinfo [5]),
    .e(i_data[12]),
    .o(o_decinfo[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u27 (
    .a(i_data[6]),
    .b(i_data[5]),
    .o(_al_u27_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'h00080000))
    _al_u270 (
    .a(_al_u201_o),
    .b(_al_u66_o),
    .c(i_data[22]),
    .d(i_data[21]),
    .e(i_data[20]),
    .o(\u_DECODE/inst_ebreak ));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~(~B*~(~E*C))))"),
    .INIT(32'h11550155))
    _al_u271 (
    .a(\u_DECODE/inst_ebreak ),
    .b(o_decinfo_grp[1]),
    .c(\u_DECODE/n3_lutinv ),
    .d(\u_DECODE/lsuinfo [2]),
    .e(i_data[14]),
    .o(_al_u271_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(D*~(~C*~B)))"),
    .INIT(16'hfd55))
    _al_u272 (
    .a(_al_u271_o),
    .b(o_decinfo_grp[3]),
    .c(_al_u265_o),
    .d(\u_DECODE/func_001_lutinv ),
    .o(o_decinfo[2]));
  AL_MAP_LUT4 #(
    .EQN("(C*(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D))"),
    .INIT(16'hc050))
    _al_u273 (
    .a(_al_u268_o),
    .b(\u_DECODE/n3_lutinv ),
    .c(_al_u158_o),
    .d(i_data[12]),
    .o(\u_DECODE/n71 [7]));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(B*~(D*C)))"),
    .INIT(16'haeee))
    _al_u274 (
    .a(\u_DECODE/n71 [7]),
    .b(\u_DECODE/n57 [0]),
    .c(_al_u124_o),
    .d(i_data[13]),
    .o(o_decinfo[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u275 (
    .a(o_rs2rdata[10]),
    .b(o_imm[10]),
    .c(_al_u156_o),
    .o(o_exu_op2[10]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hf7a7ff2e))
    _al_u276 (
    .a(i_data[6]),
    .b(i_data[5]),
    .c(i_data[4]),
    .d(i_data[3]),
    .e(i_data[2]),
    .o(_al_u276_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u277 (
    .a(i_data[11]),
    .b(i_data[10]),
    .c(i_data[9]),
    .d(i_data[7]),
    .o(_al_u277_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u278 (
    .a(_al_u276_o),
    .b(_al_u277_o),
    .c(i_data[8]),
    .o(o_rdwen));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*A*~(~E*~D))"),
    .INIT(32'h08080800))
    _al_u279 (
    .a(_al_u26_o),
    .b(_al_u27_o),
    .c(i_data[14]),
    .d(i_data[13]),
    .e(i_data[12]),
    .o(_al_u279_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u28 (
    .a(_al_u26_o),
    .b(_al_u27_o),
    .o(o_decinfo_grp[4]));
  AL_MAP_LUT5 #(
    .EQN("(~D*(~E*~((~C*B))*~(A)+~E*(~C*B)*~(A)+~(~E)*(~C*B)*A+~E*(~C*B)*A))"),
    .INIT(32'h0008005d))
    _al_u280 (
    .a(i_data[6]),
    .b(i_data[5]),
    .c(i_data[4]),
    .d(i_data[3]),
    .e(i_data[2]),
    .o(\u_DECODE/n42_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(~C*~A))"),
    .INIT(8'h32))
    _al_u281 (
    .a(_al_u279_o),
    .b(_al_u124_o),
    .c(\u_DECODE/n42_lutinv ),
    .o(rs1ren));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(~D*~A))"),
    .INIT(16'h0c08))
    _al_u282 (
    .a(_al_u279_o),
    .b(i_data_vld),
    .c(_al_u124_o),
    .d(\u_DECODE/n42_lutinv ),
    .o(o_bpu_rs1ren));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u29 (
    .a(i_data[6]),
    .b(i_data[4]),
    .c(i_data[3]),
    .d(i_data[2]),
    .o(\u_DECODE/n21_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u30 (
    .a(\u_DECODE/n21_lutinv ),
    .b(i_data[5]),
    .o(rs1topc_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u31 (
    .a(rs1_rdata[9]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[9]),
    .o(o_exu_op1[9]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u32 (
    .a(rs1_rdata[8]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[8]),
    .o(o_exu_op1[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u33 (
    .a(rs1_rdata[7]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[7]),
    .o(o_exu_op1[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u34 (
    .a(rs1_rdata[6]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[6]),
    .o(o_exu_op1[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u35 (
    .a(rs1_rdata[5]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[5]),
    .o(o_exu_op1[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u36 (
    .a(rs1_rdata[4]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[4]),
    .o(o_exu_op1[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u37 (
    .a(rs1_rdata[31]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[31]),
    .o(o_exu_op1[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u38 (
    .a(rs1_rdata[30]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[30]),
    .o(o_exu_op1[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u39 (
    .a(rs1_rdata[3]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[3]),
    .o(o_exu_op1[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u40 (
    .a(rs1_rdata[29]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[29]),
    .o(o_exu_op1[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u41 (
    .a(rs1_rdata[28]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[28]),
    .o(o_exu_op1[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u42 (
    .a(rs1_rdata[27]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[27]),
    .o(o_exu_op1[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u43 (
    .a(rs1_rdata[26]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[26]),
    .o(o_exu_op1[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u44 (
    .a(rs1_rdata[25]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[25]),
    .o(o_exu_op1[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u45 (
    .a(rs1_rdata[24]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[24]),
    .o(o_exu_op1[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u46 (
    .a(rs1_rdata[23]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[23]),
    .o(o_exu_op1[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u47 (
    .a(rs1_rdata[22]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[22]),
    .o(o_exu_op1[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u48 (
    .a(rs1_rdata[21]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[21]),
    .o(o_exu_op1[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u49 (
    .a(rs1_rdata[20]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[20]),
    .o(o_exu_op1[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u50 (
    .a(rs1_rdata[2]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[2]),
    .o(o_exu_op1[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u51 (
    .a(rs1_rdata[19]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[19]),
    .o(o_exu_op1[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u52 (
    .a(rs1_rdata[18]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[18]),
    .o(o_exu_op1[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u53 (
    .a(rs1_rdata[17]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[17]),
    .o(o_exu_op1[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u54 (
    .a(rs1_rdata[16]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[16]),
    .o(o_exu_op1[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u55 (
    .a(rs1_rdata[15]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[15]),
    .o(o_exu_op1[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u56 (
    .a(rs1_rdata[14]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[14]),
    .o(o_exu_op1[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u57 (
    .a(rs1_rdata[13]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[13]),
    .o(o_exu_op1[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u58 (
    .a(rs1_rdata[12]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[12]),
    .o(o_exu_op1[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u59 (
    .a(rs1_rdata[11]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[11]),
    .o(o_exu_op1[11]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u60 (
    .a(rs1_rdata[10]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[10]),
    .o(o_exu_op1[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u61 (
    .a(rs1_rdata[1]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[1]),
    .o(o_exu_op1[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u62 (
    .a(rs1_rdata[0]),
    .b(rs1topc_lutinv),
    .c(o_iaddr[0]),
    .o(o_exu_op1[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u63 (
    .a(i_data[3]),
    .b(i_data[2]),
    .o(_al_u63_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u64 (
    .a(_al_u63_o),
    .b(i_data[6]),
    .c(i_data[4]),
    .o(o_decinfo_grp[1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u65 (
    .a(i_data[31]),
    .b(i_data[30]),
    .c(i_data[29]),
    .d(i_data[28]),
    .o(_al_u65_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u66 (
    .a(_al_u65_o),
    .b(i_data[27]),
    .c(i_data[26]),
    .o(_al_u66_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u67 (
    .a(_al_u66_o),
    .b(i_data[25]),
    .o(\u_DECODE/func7_0000001_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u68 (
    .a(_al_u26_o),
    .b(i_data[6]),
    .c(i_data[5]),
    .o(\u_DECODE/opc_op_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u69 (
    .a(\u_DECODE/func7_0000001_lutinv ),
    .b(\u_DECODE/opc_op_lutinv ),
    .o(o_decinfo_grp[3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u70 (
    .a(i_data[13]),
    .b(i_data[12]),
    .o(\u_DECODE/lsuinfo [2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u71 (
    .a(\u_DECODE/lsuinfo [2]),
    .b(i_data[14]),
    .o(\u_DECODE/func_000_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u72 (
    .a(o_decinfo_grp[4]),
    .b(\u_DECODE/func_000_lutinv ),
    .o(\u_DECODE/n57 [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u73 (
    .a(\u_DECODE/n57 [0]),
    .b(i_data[31]),
    .o(o_csridx[11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u74 (
    .a(\u_DECODE/n57 [0]),
    .b(i_data[30]),
    .o(o_csridx[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u75 (
    .a(\u_DECODE/n57 [0]),
    .b(i_data[29]),
    .o(o_csridx[9]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u76 (
    .a(\u_DECODE/n57 [0]),
    .b(i_data[28]),
    .o(o_csridx[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u77 (
    .a(\u_DECODE/n57 [0]),
    .b(i_data[27]),
    .o(o_csridx[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u78 (
    .a(\u_DECODE/n57 [0]),
    .b(i_data[26]),
    .o(o_csridx[6]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u79 (
    .a(\u_DECODE/n57 [0]),
    .b(i_data[25]),
    .o(o_csridx[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u80 (
    .a(\u_DECODE/n57 [0]),
    .b(i_data[24]),
    .o(o_csridx[4]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u81 (
    .a(\u_DECODE/n57 [0]),
    .b(i_data[23]),
    .o(o_csridx[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u82 (
    .a(\u_DECODE/n57 [0]),
    .b(i_data[22]),
    .o(o_csridx[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u83 (
    .a(\u_DECODE/n57 [0]),
    .b(i_data[21]),
    .o(o_csridx[1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u84 (
    .a(\u_DECODE/n57 [0]),
    .b(i_data[20]),
    .o(o_csridx[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u85 (
    .a(o_decinfo_grp[4]),
    .b(i_data[19]),
    .c(i_data[14]),
    .o(o_csr_zimm[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u86 (
    .a(o_decinfo_grp[4]),
    .b(i_data[18]),
    .c(i_data[14]),
    .o(o_csr_zimm[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u87 (
    .a(o_decinfo_grp[4]),
    .b(i_data[17]),
    .c(i_data[14]),
    .o(o_csr_zimm[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u88 (
    .a(o_decinfo_grp[4]),
    .b(i_data[16]),
    .c(i_data[14]),
    .o(o_csr_zimm[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u89 (
    .a(o_decinfo_grp[4]),
    .b(i_data[15]),
    .c(i_data[14]),
    .o(o_csr_zimm[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u90 (
    .a(i_data[6]),
    .b(i_data[5]),
    .c(i_data[4]),
    .d(i_data[2]),
    .o(\u_DECODE/bjuinfo [1]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u91 (
    .a(i_data[1]),
    .b(i_data[0]),
    .o(\u_DECODE/opc_rv32 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    _al_u92 (
    .a(i_data_vld),
    .b(\u_DECODE/bjuinfo [1]),
    .c(\u_DECODE/opc_rv32 ),
    .d(i_data[20]),
    .e(i_data[3]),
    .o(\u_DECODE/n5 [0]));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*A*~(~E*D))"),
    .INIT(32'h08080008))
    _al_u93 (
    .a(i_data[6]),
    .b(i_data[5]),
    .c(i_data[4]),
    .d(i_data[3]),
    .e(i_data[2]),
    .o(o_decinfo_grp[2]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u94 (
    .a(_al_u63_o),
    .b(i_data[5]),
    .c(i_data[4]),
    .o(\u_DECODE/n47_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u95 (
    .a(_al_u63_o),
    .b(i_data[6]),
    .c(i_data[5]),
    .o(_al_u95_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(C*B)*~(~E*D*A))"),
    .INIT(32'hc0c0eac0))
    _al_u96 (
    .a(\u_DECODE/n47_lutinv ),
    .b(_al_u95_o),
    .c(i_data[20]),
    .d(i_data[7]),
    .e(i_data[6]),
    .o(o_imm[0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u97 (
    .a(_al_u65_o),
    .b(i_data[27]),
    .c(i_data[26]),
    .d(i_data[25]),
    .o(\u_DECODE/func7_0000000_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u98 (
    .a(_al_u26_o),
    .b(i_data[6]),
    .c(i_data[5]),
    .o(\u_DECODE/opc_opimm_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u99 (
    .a(\u_DECODE/func7_0000000_lutinv ),
    .b(\u_DECODE/opc_op_lutinv ),
    .c(\u_DECODE/opc_opimm_lutinv ),
    .o(_al_u99_o));
  EG_PHY_LSLICE #(
    //.MACRO("u_BPU_BP/add0/ucin_al_u283"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_BPU_BP/add0/u11_al_u286  (
    .a({rs1_rdata[13],rs1_rdata[11]}),
    .b({rs1_rdata[14],rs1_rdata[12]}),
    .c(2'b00),
    .d({bp_imm[13],bp_imm[11]}),
    .e({bp_imm[14],bp_imm[12]}),
    .fci(\u_BPU_BP/add0/c11 ),
    .f({\u_BPU_BP/n2 [13],\u_BPU_BP/n2 [11]}),
    .fco(\u_BPU_BP/add0/c15 ),
    .fx({\u_BPU_BP/n2 [14],\u_BPU_BP/n2 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_BPU_BP/add0/ucin_al_u283"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_BPU_BP/add0/u15_al_u287  (
    .a({rs1_rdata[17],rs1_rdata[15]}),
    .b({rs1_rdata[18],rs1_rdata[16]}),
    .c(2'b00),
    .d({bp_imm[17],bp_imm[15]}),
    .e({bp_imm[18],bp_imm[16]}),
    .fci(\u_BPU_BP/add0/c15 ),
    .f({\u_BPU_BP/n2 [17],\u_BPU_BP/n2 [15]}),
    .fco(\u_BPU_BP/add0/c19 ),
    .fx({\u_BPU_BP/n2 [18],\u_BPU_BP/n2 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_BPU_BP/add0/ucin_al_u283"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_BPU_BP/add0/u19_al_u288  (
    .a({rs1_rdata[21],rs1_rdata[19]}),
    .b({rs1_rdata[22],rs1_rdata[20]}),
    .c(2'b00),
    .d({bp_imm[31],bp_imm[19]}),
    .e({bp_imm[31],bp_imm[31]}),
    .fci(\u_BPU_BP/add0/c19 ),
    .f({\u_BPU_BP/n2 [21],\u_BPU_BP/n2 [19]}),
    .fco(\u_BPU_BP/add0/c23 ),
    .fx({\u_BPU_BP/n2 [22],\u_BPU_BP/n2 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_BPU_BP/add0/ucin_al_u283"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_BPU_BP/add0/u23_al_u289  (
    .a({rs1_rdata[25],rs1_rdata[23]}),
    .b({rs1_rdata[26],rs1_rdata[24]}),
    .c(2'b00),
    .d({bp_imm[31],bp_imm[31]}),
    .e({bp_imm[31],bp_imm[31]}),
    .fci(\u_BPU_BP/add0/c23 ),
    .f({\u_BPU_BP/n2 [25],\u_BPU_BP/n2 [23]}),
    .fco(\u_BPU_BP/add0/c27 ),
    .fx({\u_BPU_BP/n2 [26],\u_BPU_BP/n2 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_BPU_BP/add0/ucin_al_u283"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_BPU_BP/add0/u27_al_u290  (
    .a({rs1_rdata[29],rs1_rdata[27]}),
    .b({rs1_rdata[30],rs1_rdata[28]}),
    .c(2'b00),
    .d({bp_imm[31],bp_imm[31]}),
    .e({bp_imm[31],bp_imm[31]}),
    .fci(\u_BPU_BP/add0/c27 ),
    .f({\u_BPU_BP/n2 [29],\u_BPU_BP/n2 [27]}),
    .fco(\u_BPU_BP/add0/c31 ),
    .fx({\u_BPU_BP/n2 [30],\u_BPU_BP/n2 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_BPU_BP/add0/ucin_al_u283"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_BPU_BP/add0/u31_al_u291  (
    .a({open_n90,rs1_rdata[31]}),
    .c(2'b00),
    .d({open_n95,bp_imm[31]}),
    .fci(\u_BPU_BP/add0/c31 ),
    .f({open_n112,\u_BPU_BP/n2 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_BPU_BP/add0/ucin_al_u283"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_BPU_BP/add0/u3_al_u284  (
    .a({rs1_rdata[5],rs1_rdata[3]}),
    .b({rs1_rdata[6],rs1_rdata[4]}),
    .c(2'b00),
    .d({bp_imm[5],bp_imm[3]}),
    .e({bp_imm[6],bp_imm[4]}),
    .fci(\u_BPU_BP/add0/c3 ),
    .f({\u_BPU_BP/n2 [5],\u_BPU_BP/n2 [3]}),
    .fco(\u_BPU_BP/add0/c7 ),
    .fx({\u_BPU_BP/n2 [6],\u_BPU_BP/n2 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_BPU_BP/add0/ucin_al_u283"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_BPU_BP/add0/u7_al_u285  (
    .a({rs1_rdata[9],rs1_rdata[7]}),
    .b({rs1_rdata[10],rs1_rdata[8]}),
    .c(2'b00),
    .d({bp_imm[9],bp_imm[7]}),
    .e({bp_imm[10],bp_imm[8]}),
    .fci(\u_BPU_BP/add0/c7 ),
    .f({\u_BPU_BP/n2 [9],\u_BPU_BP/n2 [7]}),
    .fco(\u_BPU_BP/add0/c11 ),
    .fx({\u_BPU_BP/n2 [10],\u_BPU_BP/n2 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_BPU_BP/add0/ucin_al_u283"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_BPU_BP/add0/ucin_al_u283  (
    .a({rs1_rdata[1],1'b0}),
    .b({rs1_rdata[2],rs1_rdata[0]}),
    .c(2'b00),
    .d({bp_imm[1],1'b1}),
    .e({bp_imm[2],\u_DECODE/n5 [0]}),
    .f({\u_BPU_BP/n2 [1],open_n171}),
    .fco(\u_BPU_BP/add0/c3 ),
    .fx({\u_BPU_BP/n2 [2],\u_BPU_BP/n2 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin  (
    .a({o_iaddr[0],1'b0}),
    .b({\u_DECODE/n5 [0],open_n174}),
    .f({\u_BPU_BP/n4 [0],open_n194}),
    .fco(\u_BPU_BP/add1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u10|u_BPU_BP/add1/u9  (
    .a(o_iaddr[10:9]),
    .b(bp_imm[10:9]),
    .fci(\u_BPU_BP/add1/c9 ),
    .f(\u_BPU_BP/n4 [10:9]),
    .fco(\u_BPU_BP/add1/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u12|u_BPU_BP/add1/u11  (
    .a(o_iaddr[12:11]),
    .b(bp_imm[12:11]),
    .fci(\u_BPU_BP/add1/c11 ),
    .f(\u_BPU_BP/n4 [12:11]),
    .fco(\u_BPU_BP/add1/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u14|u_BPU_BP/add1/u13  (
    .a(o_iaddr[14:13]),
    .b(bp_imm[14:13]),
    .fci(\u_BPU_BP/add1/c13 ),
    .f(\u_BPU_BP/n4 [14:13]),
    .fco(\u_BPU_BP/add1/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u16|u_BPU_BP/add1/u15  (
    .a(o_iaddr[16:15]),
    .b(bp_imm[16:15]),
    .fci(\u_BPU_BP/add1/c15 ),
    .f(\u_BPU_BP/n4 [16:15]),
    .fco(\u_BPU_BP/add1/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u18|u_BPU_BP/add1/u17  (
    .a(o_iaddr[18:17]),
    .b(bp_imm[18:17]),
    .fci(\u_BPU_BP/add1/c17 ),
    .f(\u_BPU_BP/n4 [18:17]),
    .fco(\u_BPU_BP/add1/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u20|u_BPU_BP/add1/u19  (
    .a(o_iaddr[20:19]),
    .b({bp_imm[31],bp_imm[19]}),
    .fci(\u_BPU_BP/add1/c19 ),
    .f(\u_BPU_BP/n4 [20:19]),
    .fco(\u_BPU_BP/add1/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u22|u_BPU_BP/add1/u21  (
    .a(o_iaddr[22:21]),
    .b({bp_imm[31],bp_imm[31]}),
    .fci(\u_BPU_BP/add1/c21 ),
    .f(\u_BPU_BP/n4 [22:21]),
    .fco(\u_BPU_BP/add1/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u24|u_BPU_BP/add1/u23  (
    .a(o_iaddr[24:23]),
    .b({bp_imm[31],bp_imm[31]}),
    .fci(\u_BPU_BP/add1/c23 ),
    .f(\u_BPU_BP/n4 [24:23]),
    .fco(\u_BPU_BP/add1/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u26|u_BPU_BP/add1/u25  (
    .a(o_iaddr[26:25]),
    .b({bp_imm[31],bp_imm[31]}),
    .fci(\u_BPU_BP/add1/c25 ),
    .f(\u_BPU_BP/n4 [26:25]),
    .fco(\u_BPU_BP/add1/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u28|u_BPU_BP/add1/u27  (
    .a(o_iaddr[28:27]),
    .b({bp_imm[31],bp_imm[31]}),
    .fci(\u_BPU_BP/add1/c27 ),
    .f(\u_BPU_BP/n4 [28:27]),
    .fco(\u_BPU_BP/add1/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u2|u_BPU_BP/add1/u1  (
    .a(o_iaddr[2:1]),
    .b(bp_imm[2:1]),
    .fci(\u_BPU_BP/add1/c1 ),
    .f(\u_BPU_BP/n4 [2:1]),
    .fco(\u_BPU_BP/add1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u30|u_BPU_BP/add1/u29  (
    .a(o_iaddr[30:29]),
    .b({bp_imm[31],bp_imm[31]}),
    .fci(\u_BPU_BP/add1/c29 ),
    .f(\u_BPU_BP/n4 [30:29]),
    .fco(\u_BPU_BP/add1/c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u31_al_u292  (
    .a({open_n463,o_iaddr[31]}),
    .b({open_n464,bp_imm[31]}),
    .fci(\u_BPU_BP/add1/c31 ),
    .f({open_n483,\u_BPU_BP/n4 [31]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u4|u_BPU_BP/add1/u3  (
    .a(o_iaddr[4:3]),
    .b(bp_imm[4:3]),
    .fci(\u_BPU_BP/add1/c3 ),
    .f(\u_BPU_BP/n4 [4:3]),
    .fco(\u_BPU_BP/add1/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u6|u_BPU_BP/add1/u5  (
    .a(o_iaddr[6:5]),
    .b(bp_imm[6:5]),
    .fci(\u_BPU_BP/add1/c5 ),
    .f(\u_BPU_BP/n4 [6:5]),
    .fco(\u_BPU_BP/add1/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_BPU_BP/add1/u0|u_BPU_BP/add1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_BPU_BP/add1/u8|u_BPU_BP/add1/u7  (
    .a(o_iaddr[8:7]),
    .b(bp_imm[8:7]),
    .fci(\u_BPU_BP/add1/c7 ),
    .f(\u_BPU_BP/n4 [8:7]),
    .fco(\u_BPU_BP/add1/c9 ));
  REGFILE u_REGFILE (
    .i_clk(i_clk),
    .i_rd_wdata(i_rd_wdata),
    .i_rdidx(i_rdidx),
    .i_rdwen(i_rdwen),
    .i_rs1idx(i_data[19:15]),
    .i_rs1ren(rs1ren),
    .i_rs2idx(i_data[24:20]),
    .i_rs2ren(rs2ren),
    .i_rstn(1'b0),
    .o_rs1_rdata(rs1_rdata),
    .o_rs2_rdata(o_rs2rdata));  // ../RTL/core/bpu.v(186)

endmodule 

module CSR_REGFILE  // ../RTL/core/csr_regfile.v(21)
  (
  i_clk,
  i_csr_ren,
  i_csr_ridx,
  i_csr_wdata,
  i_csr_wen,
  i_csr_widx,
  i_rstn,
  o_csr_rdata
  );

  input i_clk;  // ../RTL/core/csr_regfile.v(22)
  input i_csr_ren;  // ../RTL/core/csr_regfile.v(26)
  input [11:0] i_csr_ridx;  // ../RTL/core/csr_regfile.v(27)
  input [31:0] i_csr_wdata;  // ../RTL/core/csr_regfile.v(32)
  input i_csr_wen;  // ../RTL/core/csr_regfile.v(30)
  input [11:0] i_csr_widx;  // ../RTL/core/csr_regfile.v(31)
  input i_rstn;  // ../RTL/core/csr_regfile.v(23)
  output [31:0] o_csr_rdata;  // ../RTL/core/csr_regfile.v(28)

  wire [31:0] fctrl;  // ../RTL/core/csr_regfile.v(128)
  wire [31:0] fop1;  // ../RTL/core/csr_regfile.v(129)
  wire [31:0] fop2;  // ../RTL/core/csr_regfile.v(130)
  wire [31:0] fres0_add;  // ../RTL/core/csr_regfile.v(131)
  wire [31:0] fres0_mul;  // ../RTL/core/csr_regfile.v(133)
  wire [31:0] fres0_sub;  // ../RTL/core/csr_regfile.v(132)
  wire [31:2] mtvec_base;  // ../RTL/core/csr_regfile.v(60)
  wire [1:0] mtvec_mode;  // ../RTL/core/csr_regfile.v(61)
  wire [31:0] n39;
  wire _al_u100_o;
  wire _al_u101_o;
  wire _al_u103_o;
  wire _al_u104_o;
  wire _al_u105_o;
  wire _al_u107_o;
  wire _al_u108_o;
  wire _al_u110_o;
  wire _al_u111_o;
  wire _al_u112_o;
  wire _al_u114_o;
  wire _al_u115_o;
  wire _al_u117_o;
  wire _al_u118_o;
  wire _al_u119_o;
  wire _al_u121_o;
  wire _al_u122_o;
  wire _al_u124_o;
  wire _al_u125_o;
  wire _al_u126_o;
  wire _al_u128_o;
  wire _al_u129_o;
  wire _al_u130_o;
  wire _al_u132_o;
  wire _al_u133_o;
  wire _al_u134_o;
  wire _al_u136_o;
  wire _al_u137_o;
  wire _al_u139_o;
  wire _al_u140_o;
  wire _al_u141_o;
  wire _al_u143_o;
  wire _al_u144_o;
  wire _al_u145_o;
  wire _al_u147_o;
  wire _al_u148_o;
  wire _al_u150_o;
  wire _al_u151_o;
  wire _al_u152_o;
  wire _al_u155_o;
  wire _al_u156_o;
  wire _al_u157_o;
  wire _al_u159_o;
  wire _al_u160_o;
  wire _al_u161_o;
  wire _al_u24_o;
  wire _al_u25_o;
  wire _al_u26_o;
  wire _al_u27_o;
  wire _al_u29_o;
  wire _al_u31_o;
  wire _al_u34_o;
  wire _al_u35_o;
  wire _al_u36_o;
  wire _al_u37_o;
  wire _al_u39_o;
  wire _al_u42_o;
  wire _al_u44_o;
  wire _al_u45_o;
  wire _al_u46_o;
  wire _al_u48_o;
  wire _al_u49_o;
  wire _al_u50_o;
  wire _al_u52_o;
  wire _al_u53_o;
  wire _al_u54_o;
  wire _al_u56_o;
  wire _al_u57_o;
  wire _al_u58_o;
  wire _al_u60_o;
  wire _al_u61_o;
  wire _al_u62_o;
  wire _al_u64_o;
  wire _al_u65_o;
  wire _al_u66_o;
  wire _al_u68_o;
  wire _al_u69_o;
  wire _al_u70_o;
  wire _al_u72_o;
  wire _al_u73_o;
  wire _al_u74_o;
  wire _al_u76_o;
  wire _al_u77_o;
  wire _al_u79_o;
  wire _al_u80_o;
  wire _al_u81_o;
  wire _al_u83_o;
  wire _al_u84_o;
  wire _al_u86_o;
  wire _al_u87_o;
  wire _al_u89_o;
  wire _al_u90_o;
  wire _al_u92_o;
  wire _al_u93_o;
  wire _al_u95_o;
  wire _al_u96_o;
  wire _al_u97_o;
  wire _al_u99_o;
  wire n1;
  wire n11;
  wire n14;
  wire n17;
  wire n22_lutinv;
  wire n26_lutinv;
  wire n27_lutinv;
  wire n28_lutinv;
  wire n29_lutinv;

  assign o_csr_rdata[31] = n39[31];
  assign o_csr_rdata[30] = n39[30];
  assign o_csr_rdata[29] = n39[29];
  assign o_csr_rdata[28] = n39[28];
  assign o_csr_rdata[27] = n39[27];
  assign o_csr_rdata[26] = n39[26];
  assign o_csr_rdata[25] = n39[25];
  assign o_csr_rdata[24] = n39[24];
  assign o_csr_rdata[23] = n39[23];
  assign o_csr_rdata[22] = n39[22];
  assign o_csr_rdata[21] = n39[21];
  assign o_csr_rdata[20] = n39[20];
  assign o_csr_rdata[19] = n39[19];
  assign o_csr_rdata[18] = n39[18];
  assign o_csr_rdata[17] = n39[17];
  assign o_csr_rdata[16] = n39[16];
  assign o_csr_rdata[15] = n39[15];
  assign o_csr_rdata[14] = n39[14];
  assign o_csr_rdata[13] = n39[13];
  assign o_csr_rdata[12] = n39[12];
  assign o_csr_rdata[11] = n39[11];
  assign o_csr_rdata[10] = n39[10];
  assign o_csr_rdata[9] = n39[9];
  assign o_csr_rdata[8] = n39[8];
  assign o_csr_rdata[7] = n39[7];
  assign o_csr_rdata[6] = n39[6];
  assign o_csr_rdata[5] = n39[5];
  assign o_csr_rdata[4] = n39[4];
  assign o_csr_rdata[3] = n39[3];
  assign o_csr_rdata[2] = n39[2];
  assign o_csr_rdata[1] = n39[1];
  assign o_csr_rdata[0] = n39[0];
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u100 (
    .a(fres0_add[23]),
    .b(fres0_mul[23]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u100_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u101 (
    .a(_al_u99_o),
    .b(n29_lutinv),
    .c(fop2[23]),
    .o(_al_u101_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u102 (
    .a(_al_u100_o),
    .b(fres0_sub[23]),
    .c(_al_u101_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[23]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u103 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[22]),
    .d(mtvec_base[22]),
    .o(_al_u103_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u104 (
    .a(fres0_add[22]),
    .b(fres0_mul[22]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u104_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u105 (
    .a(_al_u103_o),
    .b(n29_lutinv),
    .c(fop2[22]),
    .o(_al_u105_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u106 (
    .a(_al_u104_o),
    .b(fres0_sub[22]),
    .c(_al_u105_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[22]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u107 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[21]),
    .d(mtvec_base[21]),
    .o(_al_u107_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    _al_u108 (
    .a(fres0_add[21]),
    .b(fres0_sub[21]),
    .c(fres0_mul[21]),
    .d(fctrl[0]),
    .e(fctrl[1]),
    .o(_al_u108_o));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(E*C)*~(D*~A))"),
    .INIT(32'hf7f37733))
    _al_u109 (
    .a(_al_u108_o),
    .b(_al_u107_o),
    .c(n29_lutinv),
    .d(n27_lutinv),
    .e(fop2[21]),
    .o(n39[21]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u110 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[20]),
    .d(mtvec_base[20]),
    .o(_al_u110_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u111 (
    .a(fres0_add[20]),
    .b(fres0_mul[20]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u111_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u112 (
    .a(_al_u110_o),
    .b(n29_lutinv),
    .c(fop2[20]),
    .o(_al_u112_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u113 (
    .a(_al_u111_o),
    .b(fres0_sub[20]),
    .c(_al_u112_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[20]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u114 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[2]),
    .d(mtvec_base[2]),
    .o(_al_u114_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    _al_u115 (
    .a(fres0_add[2]),
    .b(fres0_sub[2]),
    .c(fres0_mul[2]),
    .d(fctrl[0]),
    .e(fctrl[1]),
    .o(_al_u115_o));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(E*C)*~(D*~A))"),
    .INIT(32'hf7f37733))
    _al_u116 (
    .a(_al_u115_o),
    .b(_al_u114_o),
    .c(n29_lutinv),
    .d(n27_lutinv),
    .e(fop2[2]),
    .o(n39[2]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u117 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[19]),
    .d(mtvec_base[19]),
    .o(_al_u117_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u118 (
    .a(fres0_add[19]),
    .b(fres0_mul[19]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u118_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u119 (
    .a(_al_u117_o),
    .b(n29_lutinv),
    .c(fop2[19]),
    .o(_al_u119_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u120 (
    .a(_al_u118_o),
    .b(fres0_sub[19]),
    .c(_al_u119_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[19]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u121 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[18]),
    .d(mtvec_base[18]),
    .o(_al_u121_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    _al_u122 (
    .a(fres0_add[18]),
    .b(fres0_sub[18]),
    .c(fres0_mul[18]),
    .d(fctrl[0]),
    .e(fctrl[1]),
    .o(_al_u122_o));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(E*C)*~(D*~A))"),
    .INIT(32'hf7f37733))
    _al_u123 (
    .a(_al_u122_o),
    .b(_al_u121_o),
    .c(n29_lutinv),
    .d(n27_lutinv),
    .e(fop2[18]),
    .o(n39[18]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u124 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[17]),
    .d(mtvec_base[17]),
    .o(_al_u124_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u125 (
    .a(fres0_add[17]),
    .b(fres0_mul[17]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u125_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u126 (
    .a(_al_u124_o),
    .b(n29_lutinv),
    .c(fop2[17]),
    .o(_al_u126_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u127 (
    .a(_al_u125_o),
    .b(fres0_sub[17]),
    .c(_al_u126_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[17]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u128 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[16]),
    .d(mtvec_base[16]),
    .o(_al_u128_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u129 (
    .a(fres0_add[16]),
    .b(fres0_mul[16]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u129_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u130 (
    .a(_al_u128_o),
    .b(n29_lutinv),
    .c(fop2[16]),
    .o(_al_u130_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u131 (
    .a(_al_u129_o),
    .b(fres0_sub[16]),
    .c(_al_u130_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[16]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u132 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[15]),
    .d(mtvec_base[15]),
    .o(_al_u132_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u133 (
    .a(fres0_add[15]),
    .b(fres0_mul[15]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u133_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u134 (
    .a(_al_u132_o),
    .b(n29_lutinv),
    .c(fop2[15]),
    .o(_al_u134_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u135 (
    .a(_al_u133_o),
    .b(fres0_sub[15]),
    .c(_al_u134_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[15]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u136 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[14]),
    .d(mtvec_base[14]),
    .o(_al_u136_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    _al_u137 (
    .a(fres0_add[14]),
    .b(fres0_sub[14]),
    .c(fres0_mul[14]),
    .d(fctrl[0]),
    .e(fctrl[1]),
    .o(_al_u137_o));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(E*C)*~(D*~A))"),
    .INIT(32'hf7f37733))
    _al_u138 (
    .a(_al_u137_o),
    .b(_al_u136_o),
    .c(n29_lutinv),
    .d(n27_lutinv),
    .e(fop2[14]),
    .o(n39[14]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u139 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[13]),
    .d(mtvec_base[13]),
    .o(_al_u139_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u140 (
    .a(fres0_add[13]),
    .b(fres0_mul[13]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u140_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u141 (
    .a(_al_u139_o),
    .b(n29_lutinv),
    .c(fop2[13]),
    .o(_al_u141_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u142 (
    .a(_al_u140_o),
    .b(fres0_sub[13]),
    .c(_al_u141_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[13]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u143 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[12]),
    .d(mtvec_base[12]),
    .o(_al_u143_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u144 (
    .a(fres0_add[12]),
    .b(fres0_mul[12]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u144_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u145 (
    .a(_al_u143_o),
    .b(n29_lutinv),
    .c(fop2[12]),
    .o(_al_u145_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u146 (
    .a(_al_u144_o),
    .b(fres0_sub[12]),
    .c(_al_u145_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[12]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u147 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[11]),
    .d(mtvec_base[11]),
    .o(_al_u147_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    _al_u148 (
    .a(fres0_add[11]),
    .b(fres0_sub[11]),
    .c(fres0_mul[11]),
    .d(fctrl[0]),
    .e(fctrl[1]),
    .o(_al_u148_o));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(E*C)*~(D*~A))"),
    .INIT(32'hf7f37733))
    _al_u149 (
    .a(_al_u148_o),
    .b(_al_u147_o),
    .c(n29_lutinv),
    .d(n27_lutinv),
    .e(fop2[11]),
    .o(n39[11]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u150 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[10]),
    .d(mtvec_base[10]),
    .o(_al_u150_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u151 (
    .a(fres0_add[10]),
    .b(fres0_mul[10]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u151_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u152 (
    .a(_al_u150_o),
    .b(n29_lutinv),
    .c(fop2[10]),
    .o(_al_u152_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u153 (
    .a(_al_u151_o),
    .b(fres0_sub[10]),
    .c(_al_u152_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[10]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    _al_u154 (
    .a(_al_u35_o),
    .b(_al_u36_o),
    .c(i_csr_ridx[2]),
    .d(i_csr_ridx[1]),
    .e(i_csr_ridx[0]),
    .o(n26_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u155 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(mtvec_mode[1]),
    .d(fop1[1]),
    .o(_al_u155_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u156 (
    .a(_al_u155_o),
    .b(n26_lutinv),
    .c(fctrl[1]),
    .o(_al_u156_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    _al_u157 (
    .a(fres0_add[1]),
    .b(fres0_sub[1]),
    .c(fres0_mul[1]),
    .d(fctrl[0]),
    .e(fctrl[1]),
    .o(_al_u157_o));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(E*C)*~(D*~A))"),
    .INIT(32'hf7f37733))
    _al_u158 (
    .a(_al_u157_o),
    .b(_al_u156_o),
    .c(n29_lutinv),
    .d(n27_lutinv),
    .e(fop2[1]),
    .o(n39[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u159 (
    .a(n28_lutinv),
    .b(n26_lutinv),
    .c(fctrl[0]),
    .d(fop1[0]),
    .o(_al_u159_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u160 (
    .a(_al_u159_o),
    .b(n22_lutinv),
    .c(mtvec_mode[0]),
    .o(_al_u160_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    _al_u161 (
    .a(fres0_add[0]),
    .b(fres0_sub[0]),
    .c(fres0_mul[0]),
    .d(fctrl[0]),
    .e(fctrl[1]),
    .o(_al_u161_o));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(E*C)*~(D*~A))"),
    .INIT(32'hf7f37733))
    _al_u162 (
    .a(_al_u161_o),
    .b(_al_u160_o),
    .c(n29_lutinv),
    .d(n27_lutinv),
    .e(fop2[0]),
    .o(n39[0]));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u24 (
    .a(i_csr_widx[5]),
    .b(i_csr_widx[4]),
    .c(i_csr_widx[3]),
    .o(_al_u24_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u25 (
    .a(_al_u24_o),
    .b(i_csr_wen),
    .c(i_csr_widx[0]),
    .o(_al_u25_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u26 (
    .a(i_csr_widx[9]),
    .b(i_csr_widx[8]),
    .c(i_csr_widx[7]),
    .d(i_csr_widx[6]),
    .o(_al_u26_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u27 (
    .a(_al_u26_o),
    .b(i_csr_widx[11]),
    .c(i_csr_widx[10]),
    .o(_al_u27_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u28 (
    .a(_al_u27_o),
    .b(_al_u25_o),
    .c(i_csr_widx[2]),
    .d(i_csr_widx[1]),
    .o(n11));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u29 (
    .a(i_csr_wen),
    .b(i_csr_widx[5]),
    .c(i_csr_widx[4]),
    .d(i_csr_widx[0]),
    .o(_al_u29_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    _al_u30 (
    .a(_al_u27_o),
    .b(_al_u29_o),
    .c(i_csr_widx[3]),
    .d(i_csr_widx[2]),
    .e(i_csr_widx[1]),
    .o(n1));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u31 (
    .a(_al_u24_o),
    .b(i_csr_wen),
    .c(i_csr_widx[0]),
    .o(_al_u31_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u32 (
    .a(_al_u27_o),
    .b(_al_u31_o),
    .c(i_csr_widx[2]),
    .d(i_csr_widx[1]),
    .o(n17));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u33 (
    .a(_al_u27_o),
    .b(_al_u25_o),
    .c(i_csr_widx[2]),
    .d(i_csr_widx[1]),
    .o(n14));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u34 (
    .a(i_csr_ridx[9]),
    .b(i_csr_ridx[8]),
    .c(i_csr_ridx[7]),
    .d(i_csr_ridx[6]),
    .o(_al_u34_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u35 (
    .a(_al_u34_o),
    .b(i_csr_ridx[11]),
    .c(i_csr_ridx[10]),
    .o(_al_u35_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u36 (
    .a(i_csr_ridx[5]),
    .b(i_csr_ridx[4]),
    .c(i_csr_ridx[3]),
    .o(_al_u36_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u37 (
    .a(_al_u35_o),
    .b(_al_u36_o),
    .c(i_csr_ridx[0]),
    .o(_al_u37_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u38 (
    .a(_al_u37_o),
    .b(i_csr_ridx[2]),
    .c(i_csr_ridx[1]),
    .o(n29_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u39 (
    .a(i_csr_ridx[3]),
    .b(i_csr_ridx[2]),
    .c(i_csr_ridx[1]),
    .d(i_csr_ridx[0]),
    .o(_al_u39_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u40 (
    .a(_al_u35_o),
    .b(_al_u39_o),
    .c(i_csr_ridx[5]),
    .d(i_csr_ridx[4]),
    .o(n22_lutinv));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    _al_u41 (
    .a(_al_u35_o),
    .b(_al_u36_o),
    .c(i_csr_ridx[2]),
    .d(i_csr_ridx[1]),
    .e(i_csr_ridx[0]),
    .o(n28_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u42 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[9]),
    .d(mtvec_base[9]),
    .o(_al_u42_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u43 (
    .a(_al_u37_o),
    .b(i_csr_ridx[2]),
    .c(i_csr_ridx[1]),
    .o(n27_lutinv));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u44 (
    .a(fctrl[0]),
    .b(fctrl[1]),
    .o(_al_u44_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u45 (
    .a(fres0_add[9]),
    .b(fres0_mul[9]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u45_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u46 (
    .a(_al_u42_o),
    .b(n29_lutinv),
    .c(fop2[9]),
    .o(_al_u46_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u47 (
    .a(_al_u45_o),
    .b(fres0_sub[9]),
    .c(_al_u46_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[9]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u48 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[8]),
    .d(mtvec_base[8]),
    .o(_al_u48_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u49 (
    .a(fres0_add[8]),
    .b(fres0_mul[8]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u49_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u50 (
    .a(_al_u48_o),
    .b(n29_lutinv),
    .c(fop2[8]),
    .o(_al_u50_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u51 (
    .a(_al_u49_o),
    .b(fres0_sub[8]),
    .c(_al_u50_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[8]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u52 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[7]),
    .d(mtvec_base[7]),
    .o(_al_u52_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u53 (
    .a(fres0_add[7]),
    .b(fres0_mul[7]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u53_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u54 (
    .a(_al_u52_o),
    .b(n29_lutinv),
    .c(fop2[7]),
    .o(_al_u54_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u55 (
    .a(_al_u53_o),
    .b(fres0_sub[7]),
    .c(_al_u54_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[7]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u56 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[6]),
    .d(mtvec_base[6]),
    .o(_al_u56_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u57 (
    .a(fres0_add[6]),
    .b(fres0_mul[6]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u57_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u58 (
    .a(_al_u56_o),
    .b(n29_lutinv),
    .c(fop2[6]),
    .o(_al_u58_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u59 (
    .a(_al_u57_o),
    .b(fres0_sub[6]),
    .c(_al_u58_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[6]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u60 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[5]),
    .d(mtvec_base[5]),
    .o(_al_u60_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u61 (
    .a(fres0_add[5]),
    .b(fres0_mul[5]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u61_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u62 (
    .a(_al_u60_o),
    .b(n29_lutinv),
    .c(fop2[5]),
    .o(_al_u62_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u63 (
    .a(_al_u61_o),
    .b(fres0_sub[5]),
    .c(_al_u62_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[5]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u64 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[4]),
    .d(mtvec_base[4]),
    .o(_al_u64_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u65 (
    .a(fres0_add[4]),
    .b(fres0_mul[4]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u65_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u66 (
    .a(_al_u64_o),
    .b(n29_lutinv),
    .c(fop2[4]),
    .o(_al_u66_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u67 (
    .a(_al_u65_o),
    .b(fres0_sub[4]),
    .c(_al_u66_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[4]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u68 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[31]),
    .d(mtvec_base[31]),
    .o(_al_u68_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u69 (
    .a(fres0_add[31]),
    .b(fres0_mul[31]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u69_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u70 (
    .a(_al_u68_o),
    .b(n29_lutinv),
    .c(fop2[31]),
    .o(_al_u70_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u71 (
    .a(_al_u69_o),
    .b(fres0_sub[31]),
    .c(_al_u70_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[31]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u72 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[30]),
    .d(mtvec_base[30]),
    .o(_al_u72_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u73 (
    .a(fres0_add[30]),
    .b(fres0_mul[30]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u73_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u74 (
    .a(_al_u72_o),
    .b(n29_lutinv),
    .c(fop2[30]),
    .o(_al_u74_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u75 (
    .a(_al_u73_o),
    .b(fres0_sub[30]),
    .c(_al_u74_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[30]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u76 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[3]),
    .d(mtvec_base[3]),
    .o(_al_u76_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    _al_u77 (
    .a(fres0_add[3]),
    .b(fres0_sub[3]),
    .c(fres0_mul[3]),
    .d(fctrl[0]),
    .e(fctrl[1]),
    .o(_al_u77_o));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(E*C)*~(D*~A))"),
    .INIT(32'hf7f37733))
    _al_u78 (
    .a(_al_u77_o),
    .b(_al_u76_o),
    .c(n29_lutinv),
    .d(n27_lutinv),
    .e(fop2[3]),
    .o(n39[3]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u79 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[29]),
    .d(mtvec_base[29]),
    .o(_al_u79_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u80 (
    .a(fres0_add[29]),
    .b(fres0_mul[29]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u80_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u81 (
    .a(_al_u79_o),
    .b(n29_lutinv),
    .c(fop2[29]),
    .o(_al_u81_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u82 (
    .a(_al_u80_o),
    .b(fres0_sub[29]),
    .c(_al_u81_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[29]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u83 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[28]),
    .d(mtvec_base[28]),
    .o(_al_u83_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    _al_u84 (
    .a(fres0_add[28]),
    .b(fres0_sub[28]),
    .c(fres0_mul[28]),
    .d(fctrl[0]),
    .e(fctrl[1]),
    .o(_al_u84_o));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(E*C)*~(D*~A))"),
    .INIT(32'hf7f37733))
    _al_u85 (
    .a(_al_u84_o),
    .b(_al_u83_o),
    .c(n29_lutinv),
    .d(n27_lutinv),
    .e(fop2[28]),
    .o(n39[28]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u86 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[27]),
    .d(mtvec_base[27]),
    .o(_al_u86_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    _al_u87 (
    .a(fres0_add[27]),
    .b(fres0_sub[27]),
    .c(fres0_mul[27]),
    .d(fctrl[0]),
    .e(fctrl[1]),
    .o(_al_u87_o));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(E*C)*~(D*~A))"),
    .INIT(32'hf7f37733))
    _al_u88 (
    .a(_al_u87_o),
    .b(_al_u86_o),
    .c(n29_lutinv),
    .d(n27_lutinv),
    .e(fop2[27]),
    .o(n39[27]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u89 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[26]),
    .d(mtvec_base[26]),
    .o(_al_u89_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    _al_u90 (
    .a(fres0_add[26]),
    .b(fres0_sub[26]),
    .c(fres0_mul[26]),
    .d(fctrl[0]),
    .e(fctrl[1]),
    .o(_al_u90_o));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(E*C)*~(D*~A))"),
    .INIT(32'hf7f37733))
    _al_u91 (
    .a(_al_u90_o),
    .b(_al_u89_o),
    .c(n29_lutinv),
    .d(n27_lutinv),
    .e(fop2[26]),
    .o(n39[26]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u92 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[25]),
    .d(mtvec_base[25]),
    .o(_al_u92_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff0f3355))
    _al_u93 (
    .a(fres0_add[25]),
    .b(fres0_sub[25]),
    .c(fres0_mul[25]),
    .d(fctrl[0]),
    .e(fctrl[1]),
    .o(_al_u93_o));
  AL_MAP_LUT5 #(
    .EQN("~(B*~(E*C)*~(D*~A))"),
    .INIT(32'hf7f37733))
    _al_u94 (
    .a(_al_u93_o),
    .b(_al_u92_o),
    .c(n29_lutinv),
    .d(n27_lutinv),
    .e(fop2[25]),
    .o(n39[25]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u95 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[24]),
    .d(mtvec_base[24]),
    .o(_al_u95_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u96 (
    .a(fres0_add[24]),
    .b(fres0_mul[24]),
    .c(fctrl[0]),
    .d(fctrl[1]),
    .o(_al_u96_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u97 (
    .a(_al_u95_o),
    .b(n29_lutinv),
    .c(fop2[24]),
    .o(_al_u97_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~(D*~(~A*~(E*B))))"),
    .INIT(32'hef0faf0f))
    _al_u98 (
    .a(_al_u96_o),
    .b(fres0_sub[24]),
    .c(_al_u97_o),
    .d(n27_lutinv),
    .e(_al_u44_o),
    .o(n39[24]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u99 (
    .a(n22_lutinv),
    .b(n28_lutinv),
    .c(fop1[23]),
    .d(mtvec_base[23]),
    .o(_al_u99_o));
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg0_b0 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[0]),
    .sr(i_rstn),
    .q(mtvec_mode[0]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg0_b1 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[1]),
    .sr(i_rstn),
    .q(mtvec_mode[1]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg1_b0 (
    .ce(n11),
    .clk(i_clk),
    .d(i_csr_wdata[0]),
    .sr(i_rstn),
    .q(fctrl[0]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg1_b1 (
    .ce(n11),
    .clk(i_clk),
    .d(i_csr_wdata[1]),
    .sr(i_rstn),
    .q(fctrl[1]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b0 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[0]),
    .sr(i_rstn),
    .q(fop1[0]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b1 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[1]),
    .sr(i_rstn),
    .q(fop1[1]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b10 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[10]),
    .sr(i_rstn),
    .q(fop1[10]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b11 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[11]),
    .sr(i_rstn),
    .q(fop1[11]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b12 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[12]),
    .sr(i_rstn),
    .q(fop1[12]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b13 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[13]),
    .sr(i_rstn),
    .q(fop1[13]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b14 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[14]),
    .sr(i_rstn),
    .q(fop1[14]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b15 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[15]),
    .sr(i_rstn),
    .q(fop1[15]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b16 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[16]),
    .sr(i_rstn),
    .q(fop1[16]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b17 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[17]),
    .sr(i_rstn),
    .q(fop1[17]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b18 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[18]),
    .sr(i_rstn),
    .q(fop1[18]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b19 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[19]),
    .sr(i_rstn),
    .q(fop1[19]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b2 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[2]),
    .sr(i_rstn),
    .q(fop1[2]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b20 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[20]),
    .sr(i_rstn),
    .q(fop1[20]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b21 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[21]),
    .sr(i_rstn),
    .q(fop1[21]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b22 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[22]),
    .sr(i_rstn),
    .q(fop1[22]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b23 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[23]),
    .sr(i_rstn),
    .q(fop1[23]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b24 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[24]),
    .sr(i_rstn),
    .q(fop1[24]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b25 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[25]),
    .sr(i_rstn),
    .q(fop1[25]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b26 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[26]),
    .sr(i_rstn),
    .q(fop1[26]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b27 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[27]),
    .sr(i_rstn),
    .q(fop1[27]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b28 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[28]),
    .sr(i_rstn),
    .q(fop1[28]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b29 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[29]),
    .sr(i_rstn),
    .q(fop1[29]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b3 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[3]),
    .sr(i_rstn),
    .q(fop1[3]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b30 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[30]),
    .sr(i_rstn),
    .q(fop1[30]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b31 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[31]),
    .sr(i_rstn),
    .q(fop1[31]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b4 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[4]),
    .sr(i_rstn),
    .q(fop1[4]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b5 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[5]),
    .sr(i_rstn),
    .q(fop1[5]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b6 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[6]),
    .sr(i_rstn),
    .q(fop1[6]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b7 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[7]),
    .sr(i_rstn),
    .q(fop1[7]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b8 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[8]),
    .sr(i_rstn),
    .q(fop1[8]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b9 (
    .ce(n14),
    .clk(i_clk),
    .d(i_csr_wdata[9]),
    .sr(i_rstn),
    .q(fop1[9]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b0 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[0]),
    .sr(i_rstn),
    .q(fop2[0]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b1 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[1]),
    .sr(i_rstn),
    .q(fop2[1]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b10 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[10]),
    .sr(i_rstn),
    .q(fop2[10]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b11 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[11]),
    .sr(i_rstn),
    .q(fop2[11]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b12 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[12]),
    .sr(i_rstn),
    .q(fop2[12]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b13 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[13]),
    .sr(i_rstn),
    .q(fop2[13]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b14 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[14]),
    .sr(i_rstn),
    .q(fop2[14]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b15 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[15]),
    .sr(i_rstn),
    .q(fop2[15]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b16 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[16]),
    .sr(i_rstn),
    .q(fop2[16]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b17 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[17]),
    .sr(i_rstn),
    .q(fop2[17]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b18 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[18]),
    .sr(i_rstn),
    .q(fop2[18]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b19 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[19]),
    .sr(i_rstn),
    .q(fop2[19]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b2 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[2]),
    .sr(i_rstn),
    .q(fop2[2]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b20 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[20]),
    .sr(i_rstn),
    .q(fop2[20]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b21 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[21]),
    .sr(i_rstn),
    .q(fop2[21]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b22 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[22]),
    .sr(i_rstn),
    .q(fop2[22]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b23 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[23]),
    .sr(i_rstn),
    .q(fop2[23]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b24 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[24]),
    .sr(i_rstn),
    .q(fop2[24]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b25 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[25]),
    .sr(i_rstn),
    .q(fop2[25]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b26 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[26]),
    .sr(i_rstn),
    .q(fop2[26]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b27 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[27]),
    .sr(i_rstn),
    .q(fop2[27]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b28 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[28]),
    .sr(i_rstn),
    .q(fop2[28]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b29 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[29]),
    .sr(i_rstn),
    .q(fop2[29]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b3 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[3]),
    .sr(i_rstn),
    .q(fop2[3]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b30 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[30]),
    .sr(i_rstn),
    .q(fop2[30]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b31 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[31]),
    .sr(i_rstn),
    .q(fop2[31]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b4 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[4]),
    .sr(i_rstn),
    .q(fop2[4]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b5 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[5]),
    .sr(i_rstn),
    .q(fop2[5]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b6 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[6]),
    .sr(i_rstn),
    .q(fop2[6]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b7 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[7]),
    .sr(i_rstn),
    .q(fop2[7]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b8 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[8]),
    .sr(i_rstn),
    .q(fop2[8]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg3_b9 (
    .ce(n17),
    .clk(i_clk),
    .d(i_csr_wdata[9]),
    .sr(i_rstn),
    .q(fop2[9]));  // ../RTL/core/csr_regfile.v(139)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b0 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[2]),
    .sr(i_rstn),
    .q(mtvec_base[2]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b1 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[3]),
    .sr(i_rstn),
    .q(mtvec_base[3]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b10 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[12]),
    .sr(i_rstn),
    .q(mtvec_base[12]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b11 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[13]),
    .sr(i_rstn),
    .q(mtvec_base[13]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b12 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[14]),
    .sr(i_rstn),
    .q(mtvec_base[14]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b13 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[15]),
    .sr(i_rstn),
    .q(mtvec_base[15]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b14 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[16]),
    .sr(i_rstn),
    .q(mtvec_base[16]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b15 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[17]),
    .sr(i_rstn),
    .q(mtvec_base[17]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b16 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[18]),
    .sr(i_rstn),
    .q(mtvec_base[18]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b17 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[19]),
    .sr(i_rstn),
    .q(mtvec_base[19]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b18 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[20]),
    .sr(i_rstn),
    .q(mtvec_base[20]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b19 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[21]),
    .sr(i_rstn),
    .q(mtvec_base[21]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b2 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[4]),
    .sr(i_rstn),
    .q(mtvec_base[4]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b20 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[22]),
    .sr(i_rstn),
    .q(mtvec_base[22]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b21 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[23]),
    .sr(i_rstn),
    .q(mtvec_base[23]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b22 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[24]),
    .sr(i_rstn),
    .q(mtvec_base[24]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b23 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[25]),
    .sr(i_rstn),
    .q(mtvec_base[25]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b24 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[26]),
    .sr(i_rstn),
    .q(mtvec_base[26]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b25 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[27]),
    .sr(i_rstn),
    .q(mtvec_base[27]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b26 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[28]),
    .sr(i_rstn),
    .q(mtvec_base[28]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b27 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[29]),
    .sr(i_rstn),
    .q(mtvec_base[29]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b28 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[30]),
    .sr(i_rstn),
    .q(mtvec_base[30]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b29 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[31]),
    .sr(i_rstn),
    .q(mtvec_base[31]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b3 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[5]),
    .sr(i_rstn),
    .q(mtvec_base[5]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b4 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[6]),
    .sr(i_rstn),
    .q(mtvec_base[6]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b5 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[7]),
    .sr(i_rstn),
    .q(mtvec_base[7]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b6 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[8]),
    .sr(i_rstn),
    .q(mtvec_base[8]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b7 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[9]),
    .sr(i_rstn),
    .q(mtvec_base[9]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b8 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[10]),
    .sr(i_rstn),
    .q(mtvec_base[10]));  // ../RTL/core/csr_regfile.v(64)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg4_b9 (
    .ce(n1),
    .clk(i_clk),
    .d(i_csr_wdata[11]),
    .sr(i_rstn),
    .q(mtvec_base[11]));  // ../RTL/core/csr_regfile.v(64)
  FPU32 u_FPU1 (
    .i_clk(i_clk),
    .i_op1(fop1),
    .i_op2(fop2),
    .i_rsn(1'b0),
    .o_addres(fres0_add),
    .o_mulres(fres0_mul),
    .o_subres(fres0_sub));  // ../RTL/core/csr_regfile.v(157)

endmodule 

module EXU  // ../RTL/core/exu.v(14)
  (
  i_clk,
  i_csr_rdata,
  i_csr_zimm,
  i_csridx,
  i_decinfo,
  i_decinfo_grp,
  i_exu_op1,
  i_exu_op2,
  i_iaddr,
  i_imm,
  i_rdidx,
  i_rdwen,
  i_ribm_gnt,
  i_ribm_rdata,
  i_ribm_rsp,
  i_rs2rdata,
  i_rstn,
  i_vld,
  o_csr_wdata,
  o_csr_wen,
  o_csridx,
  o_exu_jaddr,
  o_exu_rdidx0,
  o_exu_rdidx1,
  o_exu_rdidx2,
  o_exu_rdwen0,
  o_exu_rdwen1,
  o_exu_rdwen2,
  o_exu_resource_match,
  o_exu_taken,
  o_lsu_working,
  o_mdu_working,
  o_rdidx0,
  o_rdidx1,
  o_rdidx2,
  o_rdwdata0,
  o_rdwdata1,
  o_rdwdata2,
  o_rdwen0,
  o_rdwen1,
  o_rdwen2,
  o_ribm_addr,
  o_ribm_mask,
  o_ribm_rdy,
  o_ribm_req,
  o_ribm_wdata,
  o_ribm_wrcs
  );

  input i_clk;  // ../RTL/core/exu.v(15)
  input [31:0] i_csr_rdata;  // ../RTL/core/exu.v(29)
  input [31:0] i_csr_zimm;  // ../RTL/core/exu.v(30)
  input [11:0] i_csridx;  // ../RTL/core/exu.v(28)
  input [9:0] i_decinfo;  // ../RTL/core/exu.v(33)
  input [5:0] i_decinfo_grp;  // ../RTL/core/exu.v(32)
  input [31:0] i_exu_op1;  // ../RTL/core/exu.v(21)
  input [31:0] i_exu_op2;  // ../RTL/core/exu.v(22)
  input [31:0] i_iaddr;  // ../RTL/core/exu.v(34)
  input [31:0] i_imm;  // ../RTL/core/exu.v(24)
  input [4:0] i_rdidx;  // ../RTL/core/exu.v(26)
  input i_rdwen;  // ../RTL/core/exu.v(25)
  input i_ribm_gnt;  // ../RTL/core/exu.v(76)
  input [31:0] i_ribm_rdata;  // ../RTL/core/exu.v(74)
  input i_ribm_rsp;  // ../RTL/core/exu.v(77)
  input [31:0] i_rs2rdata;  // ../RTL/core/exu.v(23)
  input i_rstn;  // ../RTL/core/exu.v(16)
  input i_vld;  // ../RTL/core/exu.v(18)
  output [31:0] o_csr_wdata;  // ../RTL/core/exu.v(62)
  output o_csr_wen;  // ../RTL/core/exu.v(60)
  output [11:0] o_csridx;  // ../RTL/core/exu.v(61)
  output [31:0] o_exu_jaddr;  // ../RTL/core/exu.v(66)
  output [4:0] o_exu_rdidx0;  // ../RTL/core/exu.v(39)
  output [4:0] o_exu_rdidx1;  // ../RTL/core/exu.v(41)
  output [4:0] o_exu_rdidx2;  // ../RTL/core/exu.v(43)
  output o_exu_rdwen0;  // ../RTL/core/exu.v(38)
  output o_exu_rdwen1;  // ../RTL/core/exu.v(40)
  output o_exu_rdwen2;  // ../RTL/core/exu.v(42)
  output o_exu_resource_match;  // ../RTL/core/exu.v(44)
  output o_exu_taken;  // ../RTL/core/exu.v(65)
  output o_lsu_working;  // ../RTL/core/exu.v(55)
  output o_mdu_working;  // ../RTL/core/exu.v(51)
  output [4:0] o_rdidx0;  // ../RTL/core/exu.v(49)
  output [4:0] o_rdidx1;  // ../RTL/core/exu.v(53)
  output [4:0] o_rdidx2;  // ../RTL/core/exu.v(57)
  output [31:0] o_rdwdata0;  // ../RTL/core/exu.v(50)
  output [31:0] o_rdwdata1;  // ../RTL/core/exu.v(54)
  output [31:0] o_rdwdata2;  // ../RTL/core/exu.v(58)
  output o_rdwen0;  // ../RTL/core/exu.v(48)
  output o_rdwen1;  // ../RTL/core/exu.v(52)
  output o_rdwen2;  // ../RTL/core/exu.v(56)
  output [31:0] o_ribm_addr;  // ../RTL/core/exu.v(70)
  output [3:0] o_ribm_mask;  // ../RTL/core/exu.v(72)
  output o_ribm_rdy;  // ../RTL/core/exu.v(78)
  output o_ribm_req;  // ../RTL/core/exu.v(75)
  output [31:0] o_ribm_wdata;  // ../RTL/core/exu.v(73)
  output o_ribm_wrcs;  // ../RTL/core/exu.v(71)

  wire [31:0] alu2lsu_result;  // ../RTL/core/exu.v(90)
  wire [31:0] bju_rdwdata;  // ../RTL/core/exu.v(109)
  wire [31:0] \u_EXU_ALU/alu_and ;  // ../RTL/core/exu_alu.v(51)
  wire [31:0] \u_EXU_ALU/alu_or ;  // ../RTL/core/exu_alu.v(53)
  wire [31:0] \u_EXU_ALU/alu_sll ;  // ../RTL/core/exu_alu.v(43)
  wire [31:0] \u_EXU_ALU/alu_srl ;  // ../RTL/core/exu_alu.v(45)
  wire [31:0] \u_EXU_ALU/alu_xor ;  // ../RTL/core/exu_alu.v(49)
  wire [31:0] \u_EXU_ALU/n0 ;
  wire [31:0] \u_EXU_ALU/n168 ;
  wire [31:0] \u_EXU_ALU/n33 ;
  wire [31:0] \u_EXU_BJU/bxx_nxtpc ;  // ../RTL/core/exu_bju.v(57)
  wire [63:0] \u_EXU_LSU/access2_data ;  // ../RTL/core/exu_lsu.v(209)
  wire [1:0] \u_EXU_LSU/align_mode_reg ;  // ../RTL/core/exu_lsu.v(98)
  wire [9:0] \u_EXU_LSU/lsuinfo ;  // ../RTL/core/exu_lsu.v(94)
  wire [31:0] \u_EXU_LSU/n54 ;
  wire [31:0] \u_EXU_LSU/n55 ;
  wire [29:0] \u_EXU_LSU/n59 ;
  wire [3:0] \u_EXU_LSU/n65 ;
  wire [3:0] \u_EXU_LSU/n66 ;
  wire [31:0] \u_EXU_LSU/n67 ;
  wire [31:0] \u_EXU_LSU/n76 ;
  wire [3:0] \u_EXU_LSU/n78 ;
  wire [31:0] \u_EXU_LSU/n79 ;
  wire [31:0] \u_EXU_LSU/overleft_buffer ;  // ../RTL/core/exu_lsu.v(100)
  wire [31:0] \u_EXU_LSU/rs2rdata_reg ;  // ../RTL/core/exu_lsu.v(99)
  wire [31:0] \u_EXU_SCU/n0 ;
  wire _al_u1002_o;
  wire _al_u1003_o;
  wire _al_u1004_o;
  wire _al_u1005_o;
  wire _al_u1006_o;
  wire _al_u1007_o;
  wire _al_u1009_o;
  wire _al_u1012_o;
  wire _al_u1013_o;
  wire _al_u1014_o;
  wire _al_u1015_o;
  wire _al_u1016_o;
  wire _al_u1017_o;
  wire _al_u1018_o;
  wire _al_u1019_o;
  wire _al_u1020_o;
  wire _al_u1022_o;
  wire _al_u1023_o;
  wire _al_u1024_o;
  wire _al_u1026_o;
  wire _al_u1027_o;
  wire _al_u1028_o;
  wire _al_u1029_o;
  wire _al_u1030_o;
  wire _al_u1031_o;
  wire _al_u1032_o;
  wire _al_u1033_o;
  wire _al_u1035_o;
  wire _al_u1036_o;
  wire _al_u1037_o;
  wire _al_u1038_o;
  wire _al_u1039_o;
  wire _al_u1040_o;
  wire _al_u1041_o;
  wire _al_u1043_o;
  wire _al_u1045_o;
  wire _al_u1046_o;
  wire _al_u1047_o;
  wire _al_u1048_o;
  wire _al_u1049_o;
  wire _al_u1051_o;
  wire _al_u1052_o;
  wire _al_u1055_o;
  wire _al_u1056_o;
  wire _al_u1057_o;
  wire _al_u1058_o;
  wire _al_u1059_o;
  wire _al_u1060_o;
  wire _al_u1061_o;
  wire _al_u1063_o;
  wire _al_u1064_o;
  wire _al_u1065_o;
  wire _al_u1066_o;
  wire _al_u1067_o;
  wire _al_u1068_o;
  wire _al_u1069_o;
  wire _al_u1072_o;
  wire _al_u1073_o;
  wire _al_u1075_o;
  wire _al_u1076_o;
  wire _al_u1078_o;
  wire _al_u1079_o;
  wire _al_u1080_o;
  wire _al_u1082_o;
  wire _al_u1086_o;
  wire _al_u1087_o;
  wire _al_u1088_o;
  wire _al_u1089_o;
  wire _al_u1090_o;
  wire _al_u1092_o;
  wire _al_u1093_o;
  wire _al_u1094_o;
  wire _al_u1095_o;
  wire _al_u1096_o;
  wire _al_u1097_o;
  wire _al_u1098_o;
  wire _al_u1100_o;
  wire _al_u1101_o;
  wire _al_u1102_o;
  wire _al_u1103_o;
  wire _al_u1104_o;
  wire _al_u1105_o;
  wire _al_u1106_o;
  wire _al_u1107_o;
  wire _al_u1108_o;
  wire _al_u1109_o;
  wire _al_u1110_o;
  wire _al_u1111_o;
  wire _al_u1112_o;
  wire _al_u1114_o;
  wire _al_u1115_o;
  wire _al_u1117_o;
  wire _al_u1118_o;
  wire _al_u1119_o;
  wire _al_u1120_o;
  wire _al_u1121_o;
  wire _al_u1122_o;
  wire _al_u1123_o;
  wire _al_u1124_o;
  wire _al_u1126_o;
  wire _al_u1127_o;
  wire _al_u1128_o;
  wire _al_u1129_o;
  wire _al_u1130_o;
  wire _al_u1132_o;
  wire _al_u1133_o;
  wire _al_u1134_o;
  wire _al_u1135_o;
  wire _al_u1136_o;
  wire _al_u1137_o;
  wire _al_u1138_o;
  wire _al_u1139_o;
  wire _al_u1140_o;
  wire _al_u1141_o;
  wire _al_u1142_o;
  wire _al_u1144_o;
  wire _al_u1146_o;
  wire _al_u1147_o;
  wire _al_u1149_o;
  wire _al_u1150_o;
  wire _al_u1152_o;
  wire _al_u1154_o;
  wire _al_u1156_o;
  wire _al_u1157_o;
  wire _al_u1158_o;
  wire _al_u1159_o;
  wire _al_u1160_o;
  wire _al_u1161_o;
  wire _al_u1162_o;
  wire _al_u1163_o;
  wire _al_u1164_o;
  wire _al_u1167_o;
  wire _al_u1168_o;
  wire _al_u1169_o;
  wire _al_u1172_o;
  wire _al_u1174_o;
  wire _al_u1176_o;
  wire _al_u1177_o;
  wire _al_u1178_o;
  wire _al_u1179_o;
  wire _al_u1180_o;
  wire _al_u1181_o;
  wire _al_u1182_o;
  wire _al_u1184_o;
  wire _al_u1185_o;
  wire _al_u1186_o;
  wire _al_u1187_o;
  wire _al_u1188_o;
  wire _al_u1189_o;
  wire _al_u1191_o;
  wire _al_u1193_o;
  wire _al_u1194_o;
  wire _al_u1195_o;
  wire _al_u1196_o;
  wire _al_u1197_o;
  wire _al_u1199_o;
  wire _al_u1200_o;
  wire _al_u1201_o;
  wire _al_u1203_o;
  wire _al_u1204_o;
  wire _al_u1205_o;
  wire _al_u1206_o;
  wire _al_u1207_o;
  wire _al_u1209_o;
  wire _al_u1210_o;
  wire _al_u1212_o;
  wire _al_u1213_o;
  wire _al_u1215_o;
  wire _al_u1216_o;
  wire _al_u1217_o;
  wire _al_u1218_o;
  wire _al_u1219_o;
  wire _al_u1221_o;
  wire _al_u1223_o;
  wire _al_u1224_o;
  wire _al_u1225_o;
  wire _al_u1226_o;
  wire _al_u1227_o;
  wire _al_u1228_o;
  wire _al_u1229_o;
  wire _al_u1230_o;
  wire _al_u1232_o;
  wire _al_u1233_o;
  wire _al_u1234_o;
  wire _al_u1235_o;
  wire _al_u1237_o;
  wire _al_u1238_o;
  wire _al_u1239_o;
  wire _al_u1240_o;
  wire _al_u1241_o;
  wire _al_u1242_o;
  wire _al_u1243_o;
  wire _al_u1244_o;
  wire _al_u1245_o;
  wire _al_u1247_o;
  wire _al_u1249_o;
  wire _al_u1250_o;
  wire _al_u1251_o;
  wire _al_u1252_o;
  wire _al_u1253_o;
  wire _al_u1255_o;
  wire _al_u1256_o;
  wire _al_u1257_o;
  wire _al_u1258_o;
  wire _al_u1260_o;
  wire _al_u1261_o;
  wire _al_u1262_o;
  wire _al_u1263_o;
  wire _al_u1265_o;
  wire _al_u1266_o;
  wire _al_u1267_o;
  wire _al_u1268_o;
  wire _al_u1269_o;
  wire _al_u1270_o;
  wire _al_u1271_o;
  wire _al_u1272_o;
  wire _al_u1273_o;
  wire _al_u1274_o;
  wire _al_u1275_o;
  wire _al_u1276_o;
  wire _al_u1277_o;
  wire _al_u1278_o;
  wire _al_u1279_o;
  wire _al_u1280_o;
  wire _al_u1281_o;
  wire _al_u1284_o;
  wire _al_u1285_o;
  wire _al_u1286_o;
  wire _al_u1287_o;
  wire _al_u1288_o;
  wire _al_u1289_o;
  wire _al_u1290_o;
  wire _al_u1291_o;
  wire _al_u1292_o;
  wire _al_u1293_o;
  wire _al_u1294_o;
  wire _al_u1295_o;
  wire _al_u1296_o;
  wire _al_u1297_o;
  wire _al_u1298_o;
  wire _al_u1301_o;
  wire _al_u1302_o;
  wire _al_u1304_o;
  wire _al_u1305_o;
  wire _al_u1306_o;
  wire _al_u1308_o;
  wire _al_u1309_o;
  wire _al_u1310_o;
  wire _al_u1311_o;
  wire _al_u1312_o;
  wire _al_u1313_o;
  wire _al_u1314_o;
  wire _al_u1316_o;
  wire _al_u1317_o;
  wire _al_u1318_o;
  wire _al_u1319_o;
  wire _al_u1320_o;
  wire _al_u1321_o;
  wire _al_u1322_o;
  wire _al_u1323_o;
  wire _al_u1324_o;
  wire _al_u1325_o;
  wire _al_u1326_o;
  wire _al_u1327_o;
  wire _al_u1328_o;
  wire _al_u1329_o;
  wire _al_u1330_o;
  wire _al_u1331_o;
  wire _al_u1332_o;
  wire _al_u1334_o;
  wire _al_u1335_o;
  wire _al_u1336_o;
  wire _al_u1337_o;
  wire _al_u1338_o;
  wire _al_u1339_o;
  wire _al_u1340_o;
  wire _al_u1341_o;
  wire _al_u1342_o;
  wire _al_u1343_o;
  wire _al_u1344_o;
  wire _al_u1346_o;
  wire _al_u1347_o;
  wire _al_u1348_o;
  wire _al_u1349_o;
  wire _al_u1350_o;
  wire _al_u1351_o;
  wire _al_u1353_o;
  wire _al_u1354_o;
  wire _al_u1355_o;
  wire _al_u1356_o;
  wire _al_u1358_o;
  wire _al_u1359_o;
  wire _al_u1360_o;
  wire _al_u1361_o;
  wire _al_u1362_o;
  wire _al_u1363_o;
  wire _al_u1364_o;
  wire _al_u1365_o;
  wire _al_u1366_o;
  wire _al_u1368_o;
  wire _al_u1369_o;
  wire _al_u1370_o;
  wire _al_u1371_o;
  wire _al_u1374_o;
  wire _al_u1375_o;
  wire _al_u1376_o;
  wire _al_u1377_o;
  wire _al_u1378_o;
  wire _al_u1379_o;
  wire _al_u1380_o;
  wire _al_u1382_o;
  wire _al_u1383_o;
  wire _al_u1384_o;
  wire _al_u1385_o;
  wire _al_u1387_o;
  wire _al_u1388_o;
  wire _al_u1389_o;
  wire _al_u1390_o;
  wire _al_u1392_o;
  wire _al_u1393_o;
  wire _al_u1394_o;
  wire _al_u1396_o;
  wire _al_u1397_o;
  wire _al_u1398_o;
  wire _al_u1399_o;
  wire _al_u1400_o;
  wire _al_u1401_o;
  wire _al_u1402_o;
  wire _al_u1404_o;
  wire _al_u1405_o;
  wire _al_u1406_o;
  wire _al_u1407_o;
  wire _al_u1408_o;
  wire _al_u1410_o;
  wire _al_u1411_o;
  wire _al_u1412_o;
  wire _al_u1416_o;
  wire _al_u1417_o;
  wire _al_u1418_o;
  wire _al_u1419_o;
  wire _al_u1420_o;
  wire _al_u1421_o;
  wire _al_u1423_o;
  wire _al_u1424_o;
  wire _al_u1426_o;
  wire _al_u1427_o;
  wire _al_u1428_o;
  wire _al_u1429_o;
  wire _al_u1430_o;
  wire _al_u1431_o;
  wire _al_u1432_o;
  wire _al_u1433_o;
  wire _al_u1434_o;
  wire _al_u1436_o;
  wire _al_u1437_o;
  wire _al_u1438_o;
  wire _al_u1439_o;
  wire _al_u1440_o;
  wire _al_u1441_o;
  wire _al_u1442_o;
  wire _al_u1443_o;
  wire _al_u1444_o;
  wire _al_u1446_o;
  wire _al_u1447_o;
  wire _al_u1448_o;
  wire _al_u1449_o;
  wire _al_u1451_o;
  wire _al_u1452_o;
  wire _al_u1453_o;
  wire _al_u1454_o;
  wire _al_u1455_o;
  wire _al_u1456_o;
  wire _al_u1458_o;
  wire _al_u1459_o;
  wire _al_u1461_o;
  wire _al_u1462_o;
  wire _al_u1463_o;
  wire _al_u1465_o;
  wire _al_u1466_o;
  wire _al_u1467_o;
  wire _al_u422_o;
  wire _al_u426_o;
  wire _al_u428_o;
  wire _al_u429_o;
  wire _al_u430_o;
  wire _al_u431_o;
  wire _al_u432_o;
  wire _al_u433_o;
  wire _al_u435_o;
  wire _al_u436_o;
  wire _al_u437_o;
  wire _al_u438_o;
  wire _al_u439_o;
  wire _al_u440_o;
  wire _al_u442_o;
  wire _al_u443_o;
  wire _al_u444_o;
  wire _al_u445_o;
  wire _al_u446_o;
  wire _al_u447_o;
  wire _al_u449_o;
  wire _al_u450_o;
  wire _al_u451_o;
  wire _al_u452_o;
  wire _al_u453_o;
  wire _al_u455_o;
  wire _al_u456_o;
  wire _al_u457_o;
  wire _al_u458_o;
  wire _al_u459_o;
  wire _al_u460_o;
  wire _al_u462_o;
  wire _al_u463_o;
  wire _al_u464_o;
  wire _al_u465_o;
  wire _al_u466_o;
  wire _al_u467_o;
  wire _al_u469_o;
  wire _al_u470_o;
  wire _al_u471_o;
  wire _al_u472_o;
  wire _al_u473_o;
  wire _al_u475_o;
  wire _al_u476_o;
  wire _al_u477_o;
  wire _al_u478_o;
  wire _al_u479_o;
  wire _al_u481_o;
  wire _al_u482_o;
  wire _al_u485_o;
  wire _al_u487_o;
  wire _al_u489_o;
  wire _al_u491_o;
  wire _al_u493_o;
  wire _al_u495_o;
  wire _al_u497_o;
  wire _al_u499_o;
  wire _al_u501_o;
  wire _al_u503_o;
  wire _al_u505_o;
  wire _al_u507_o;
  wire _al_u509_o;
  wire _al_u511_o;
  wire _al_u513_o;
  wire _al_u515_o;
  wire _al_u517_o;
  wire _al_u519_o;
  wire _al_u521_o;
  wire _al_u523_o;
  wire _al_u525_o;
  wire _al_u527_o;
  wire _al_u529_o;
  wire _al_u531_o;
  wire _al_u533_o;
  wire _al_u535_o;
  wire _al_u537_o;
  wire _al_u539_o;
  wire _al_u541_o;
  wire _al_u543_o;
  wire _al_u548_o;
  wire _al_u549_o;
  wire _al_u550_o;
  wire _al_u551_o;
  wire _al_u552_o;
  wire _al_u553_o;
  wire _al_u556_o;
  wire _al_u557_o;
  wire _al_u558_o;
  wire _al_u561_o;
  wire _al_u562_o;
  wire _al_u563_o;
  wire _al_u565_o;
  wire _al_u566_o;
  wire _al_u568_o;
  wire _al_u569_o;
  wire _al_u570_o;
  wire _al_u571_o;
  wire _al_u574_o;
  wire _al_u575_o;
  wire _al_u576_o;
  wire _al_u577_o;
  wire _al_u579_o;
  wire _al_u580_o;
  wire _al_u581_o;
  wire _al_u582_o;
  wire _al_u584_o;
  wire _al_u585_o;
  wire _al_u586_o;
  wire _al_u587_o;
  wire _al_u589_o;
  wire _al_u590_o;
  wire _al_u591_o;
  wire _al_u592_o;
  wire _al_u594_o;
  wire _al_u595_o;
  wire _al_u596_o;
  wire _al_u597_o;
  wire _al_u599_o;
  wire _al_u600_o;
  wire _al_u601_o;
  wire _al_u602_o;
  wire _al_u604_o;
  wire _al_u605_o;
  wire _al_u606_o;
  wire _al_u607_o;
  wire _al_u609_o;
  wire _al_u610_o;
  wire _al_u611_o;
  wire _al_u612_o;
  wire _al_u613_o;
  wire _al_u615_o;
  wire _al_u616_o;
  wire _al_u617_o;
  wire _al_u619_o;
  wire _al_u620_o;
  wire _al_u623_o;
  wire _al_u624_o;
  wire _al_u625_o;
  wire _al_u626_o;
  wire _al_u628_o;
  wire _al_u629_o;
  wire _al_u630_o;
  wire _al_u632_o;
  wire _al_u633_o;
  wire _al_u634_o;
  wire _al_u635_o;
  wire _al_u637_o;
  wire _al_u638_o;
  wire _al_u639_o;
  wire _al_u641_o;
  wire _al_u642_o;
  wire _al_u643_o;
  wire _al_u644_o;
  wire _al_u646_o;
  wire _al_u648_o;
  wire _al_u649_o;
  wire _al_u650_o;
  wire _al_u653_o;
  wire _al_u654_o;
  wire _al_u656_o;
  wire _al_u657_o;
  wire _al_u659_o;
  wire _al_u660_o;
  wire _al_u661_o;
  wire _al_u664_o;
  wire _al_u665_o;
  wire _al_u667_o;
  wire _al_u668_o;
  wire _al_u670_o;
  wire _al_u671_o;
  wire _al_u672_o;
  wire _al_u673_o;
  wire _al_u675_o;
  wire _al_u676_o;
  wire _al_u677_o;
  wire _al_u680_o;
  wire _al_u683_o;
  wire _al_u687_o;
  wire _al_u695_o;
  wire _al_u698_o;
  wire _al_u701_o;
  wire _al_u704_o;
  wire _al_u706_o;
  wire _al_u707_o;
  wire _al_u709_o;
  wire _al_u710_o;
  wire _al_u713_o;
  wire _al_u715_o;
  wire _al_u716_o;
  wire _al_u718_o;
  wire _al_u719_o;
  wire _al_u721_o;
  wire _al_u722_o;
  wire _al_u724_o;
  wire _al_u725_o;
  wire _al_u727_o;
  wire _al_u728_o;
  wire _al_u730_o;
  wire _al_u731_o;
  wire _al_u733_o;
  wire _al_u736_o;
  wire _al_u739_o;
  wire _al_u742_o;
  wire _al_u746_o;
  wire _al_u748_o;
  wire _al_u751_o;
  wire _al_u754_o;
  wire _al_u757_o;
  wire _al_u779_o;
  wire _al_u782_o;
  wire _al_u788_o;
  wire _al_u794_o;
  wire _al_u799_o;
  wire _al_u801_o;
  wire _al_u805_o;
  wire _al_u807_o;
  wire _al_u809_o;
  wire _al_u815_o;
  wire _al_u817_o;
  wire _al_u819_o;
  wire _al_u821_o;
  wire _al_u823_o;
  wire _al_u825_o;
  wire _al_u827_o;
  wire _al_u837_o;
  wire _al_u839_o;
  wire _al_u841_o;
  wire _al_u851_o;
  wire _al_u858_o;
  wire _al_u859_o;
  wire _al_u860_o;
  wire _al_u863_o;
  wire _al_u864_o;
  wire _al_u865_o;
  wire _al_u866_o;
  wire _al_u867_o;
  wire _al_u869_o;
  wire _al_u870_o;
  wire _al_u871_o;
  wire _al_u872_o;
  wire _al_u873_o;
  wire _al_u874_o;
  wire _al_u875_o;
  wire _al_u877_o;
  wire _al_u878_o;
  wire _al_u879_o;
  wire _al_u882_o;
  wire _al_u883_o;
  wire _al_u885_o;
  wire _al_u887_o;
  wire _al_u890_o;
  wire _al_u891_o;
  wire _al_u892_o;
  wire _al_u897_o;
  wire _al_u898_o;
  wire _al_u899_o;
  wire _al_u900_o;
  wire _al_u902_o;
  wire _al_u903_o;
  wire _al_u904_o;
  wire _al_u905_o;
  wire _al_u906_o;
  wire _al_u907_o;
  wire _al_u908_o;
  wire _al_u909_o;
  wire _al_u910_o;
  wire _al_u911_o;
  wire _al_u912_o;
  wire _al_u913_o;
  wire _al_u914_o;
  wire _al_u915_o;
  wire _al_u916_o;
  wire _al_u917_o;
  wire _al_u918_o;
  wire _al_u919_o;
  wire _al_u920_o;
  wire _al_u921_o;
  wire _al_u922_o;
  wire _al_u923_o;
  wire _al_u924_o;
  wire _al_u925_o;
  wire _al_u926_o;
  wire _al_u927_o;
  wire _al_u928_o;
  wire _al_u929_o;
  wire _al_u930_o;
  wire _al_u931_o;
  wire _al_u933_o;
  wire _al_u934_o;
  wire _al_u935_o;
  wire _al_u936_o;
  wire _al_u937_o;
  wire _al_u938_o;
  wire _al_u939_o;
  wire _al_u940_o;
  wire _al_u941_o;
  wire _al_u942_o;
  wire _al_u943_o;
  wire _al_u944_o;
  wire _al_u945_o;
  wire _al_u946_o;
  wire _al_u948_o;
  wire _al_u950_o;
  wire _al_u951_o;
  wire _al_u954_o;
  wire _al_u955_o;
  wire _al_u956_o;
  wire _al_u958_o;
  wire _al_u960_o;
  wire _al_u961_o;
  wire _al_u963_o;
  wire _al_u965_o;
  wire _al_u967_o;
  wire _al_u969_o;
  wire _al_u970_o;
  wire _al_u971_o;
  wire _al_u972_o;
  wire _al_u973_o;
  wire _al_u974_o;
  wire _al_u975_o;
  wire _al_u976_o;
  wire _al_u977_o;
  wire _al_u979_o;
  wire _al_u980_o;
  wire _al_u981_o;
  wire _al_u982_o;
  wire _al_u983_o;
  wire _al_u985_o;
  wire _al_u986_o;
  wire _al_u987_o;
  wire _al_u988_o;
  wire _al_u989_o;
  wire _al_u990_o;
  wire _al_u991_o;
  wire _al_u994_o;
  wire _al_u995_o;
  wire _al_u996_o;
  wire _al_u997_o;
  wire _al_u998_o;
  wire _al_u999_o;
  wire bju_rdwen;  // ../RTL/core/exu.v(108)
  wire mdu_flush;  // ../RTL/core/exu.v(172)
  wire n7_lutinv;
  wire \u_EXU_ALU/add0/c11 ;  // ../RTL/core/exu_alu.v(39)
  wire \u_EXU_ALU/add0/c15 ;  // ../RTL/core/exu_alu.v(39)
  wire \u_EXU_ALU/add0/c19 ;  // ../RTL/core/exu_alu.v(39)
  wire \u_EXU_ALU/add0/c23 ;  // ../RTL/core/exu_alu.v(39)
  wire \u_EXU_ALU/add0/c27 ;  // ../RTL/core/exu_alu.v(39)
  wire \u_EXU_ALU/add0/c3 ;  // ../RTL/core/exu_alu.v(39)
  wire \u_EXU_ALU/add0/c31 ;  // ../RTL/core/exu_alu.v(39)
  wire \u_EXU_ALU/add0/c7 ;  // ../RTL/core/exu_alu.v(39)
  wire \u_EXU_ALU/lt0_c1 ;
  wire \u_EXU_ALU/lt0_c11 ;
  wire \u_EXU_ALU/lt0_c13 ;
  wire \u_EXU_ALU/lt0_c15 ;
  wire \u_EXU_ALU/lt0_c17 ;
  wire \u_EXU_ALU/lt0_c19 ;
  wire \u_EXU_ALU/lt0_c21 ;
  wire \u_EXU_ALU/lt0_c23 ;
  wire \u_EXU_ALU/lt0_c25 ;
  wire \u_EXU_ALU/lt0_c27 ;
  wire \u_EXU_ALU/lt0_c29 ;
  wire \u_EXU_ALU/lt0_c3 ;
  wire \u_EXU_ALU/lt0_c31 ;
  wire \u_EXU_ALU/lt0_c5 ;
  wire \u_EXU_ALU/lt0_c7 ;
  wire \u_EXU_ALU/lt0_c9 ;
  wire \u_EXU_ALU/lt1_c1 ;
  wire \u_EXU_ALU/lt1_c11 ;
  wire \u_EXU_ALU/lt1_c13 ;
  wire \u_EXU_ALU/lt1_c15 ;
  wire \u_EXU_ALU/lt1_c17 ;
  wire \u_EXU_ALU/lt1_c19 ;
  wire \u_EXU_ALU/lt1_c21 ;
  wire \u_EXU_ALU/lt1_c23 ;
  wire \u_EXU_ALU/lt1_c25 ;
  wire \u_EXU_ALU/lt1_c27 ;
  wire \u_EXU_ALU/lt1_c29 ;
  wire \u_EXU_ALU/lt1_c3 ;
  wire \u_EXU_ALU/lt1_c31 ;
  wire \u_EXU_ALU/lt1_c5 ;
  wire \u_EXU_ALU/lt1_c7 ;
  wire \u_EXU_ALU/lt1_c9 ;
  wire \u_EXU_ALU/n100_lutinv ;
  wire \u_EXU_ALU/n101_lutinv ;
  wire \u_EXU_ALU/n109_lutinv ;
  wire \u_EXU_ALU/n110_lutinv ;
  wire \u_EXU_ALU/n111_lutinv ;
  wire \u_EXU_ALU/n115_lutinv ;
  wire \u_EXU_ALU/n125_lutinv ;
  wire \u_EXU_ALU/n127_lutinv ;
  wire \u_EXU_ALU/n179_neg_lutinv ;
  wire \u_EXU_ALU/n226_lutinv ;
  wire \u_EXU_ALU/n227_lutinv ;
  wire \u_EXU_ALU/n228_lutinv ;
  wire \u_EXU_ALU/n229_lutinv ;
  wire \u_EXU_ALU/n235_lutinv ;
  wire \u_EXU_ALU/n236_lutinv ;
  wire \u_EXU_ALU/n237_lutinv ;
  wire \u_EXU_ALU/n241_lutinv ;
  wire \u_EXU_ALU/n249_lutinv ;
  wire \u_EXU_ALU/n253 ;
  wire \u_EXU_ALU/n255_lutinv ;
  wire \u_EXU_ALU/n256_lutinv ;
  wire \u_EXU_ALU/n261 ;
  wire \u_EXU_ALU/n281_neg_lutinv ;
  wire \u_EXU_ALU/n327_lutinv ;
  wire \u_EXU_ALU/n351_lutinv ;
  wire \u_EXU_ALU/n352_lutinv ;
  wire \u_EXU_ALU/n362_lutinv ;
  wire \u_EXU_ALU/n363_lutinv ;
  wire \u_EXU_ALU/n365_lutinv ;
  wire \u_EXU_ALU/n366_lutinv ;
  wire \u_EXU_ALU/n369_lutinv ;
  wire \u_EXU_ALU/n370_lutinv ;
  wire \u_EXU_ALU/n371_lutinv ;
  wire \u_EXU_ALU/n372_lutinv ;
  wire \u_EXU_ALU/n373_lutinv ;
  wire \u_EXU_ALU/n374_lutinv ;
  wire \u_EXU_ALU/n375_lutinv ;
  wire \u_EXU_ALU/n379_lutinv ;
  wire \u_EXU_ALU/n402_lutinv ;
  wire \u_EXU_ALU/n413_lutinv ;
  wire \u_EXU_ALU/n416_lutinv ;
  wire \u_EXU_ALU/n45_lutinv ;
  wire \u_EXU_ALU/n46_lutinv ;
  wire \u_EXU_ALU/n49_lutinv ;
  wire \u_EXU_ALU/n77_lutinv ;
  wire \u_EXU_ALU/n80_lutinv ;
  wire \u_EXU_ALU/n83_lutinv ;
  wire \u_EXU_ALU/n84_lutinv ;
  wire \u_EXU_ALU/n88_lutinv ;
  wire \u_EXU_ALU/n92_lutinv ;
  wire \u_EXU_ALU/n96_lutinv ;
  wire \u_EXU_ALU/n97_lutinv ;
  wire \u_EXU_ALU/sub0/c11 ;  // ../RTL/core/exu_alu.v(41)
  wire \u_EXU_ALU/sub0/c15 ;  // ../RTL/core/exu_alu.v(41)
  wire \u_EXU_ALU/sub0/c19 ;  // ../RTL/core/exu_alu.v(41)
  wire \u_EXU_ALU/sub0/c23 ;  // ../RTL/core/exu_alu.v(41)
  wire \u_EXU_ALU/sub0/c27 ;  // ../RTL/core/exu_alu.v(41)
  wire \u_EXU_ALU/sub0/c3 ;  // ../RTL/core/exu_alu.v(41)
  wire \u_EXU_ALU/sub0/c31 ;  // ../RTL/core/exu_alu.v(41)
  wire \u_EXU_ALU/sub0/c7 ;  // ../RTL/core/exu_alu.v(41)
  wire \u_EXU_ALU/u1029_sel_is_0_o ;
  wire \u_EXU_BJU/add0/c11 ;  // ../RTL/core/exu_bju.v(57)
  wire \u_EXU_BJU/add0/c15 ;  // ../RTL/core/exu_bju.v(57)
  wire \u_EXU_BJU/add0/c19 ;  // ../RTL/core/exu_bju.v(57)
  wire \u_EXU_BJU/add0/c23 ;  // ../RTL/core/exu_bju.v(57)
  wire \u_EXU_BJU/add0/c27 ;  // ../RTL/core/exu_bju.v(57)
  wire \u_EXU_BJU/add0/c3 ;  // ../RTL/core/exu_bju.v(57)
  wire \u_EXU_BJU/add0/c31 ;  // ../RTL/core/exu_bju.v(57)
  wire \u_EXU_BJU/add0/c7 ;  // ../RTL/core/exu_bju.v(57)
  wire \u_EXU_BJU/add1/c11 ;  // ../RTL/core/exu_bju.v(62)
  wire \u_EXU_BJU/add1/c15 ;  // ../RTL/core/exu_bju.v(62)
  wire \u_EXU_BJU/add1/c19 ;  // ../RTL/core/exu_bju.v(62)
  wire \u_EXU_BJU/add1/c23 ;  // ../RTL/core/exu_bju.v(62)
  wire \u_EXU_BJU/add1/c27 ;  // ../RTL/core/exu_bju.v(62)
  wire \u_EXU_BJU/add1/c3 ;  // ../RTL/core/exu_bju.v(62)
  wire \u_EXU_BJU/add1/c7 ;  // ../RTL/core/exu_bju.v(62)
  wire \u_EXU_BJU/bxx_beq ;  // ../RTL/core/exu_bju.v(42)
  wire \u_EXU_BJU/bxx_bne ;  // ../RTL/core/exu_bju.v(43)
  wire \u_EXU_LSU/access2_once ;  // ../RTL/core/exu_lsu.v(96)
  wire \u_EXU_LSU/access2_vld ;  // ../RTL/core/exu_lsu.v(95)
  wire \u_EXU_LSU/add0/c1 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c11 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c13 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c15 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c17 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c19 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c21 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c23 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c25 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c27 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c29 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c3 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c5 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c7 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/add0/c9 ;  // ../RTL/core/exu_lsu.v(185)
  wire \u_EXU_LSU/handshake_once ;  // ../RTL/core/exu_lsu.v(152)
  wire \u_EXU_LSU/handshake_rdy_last ;  // ../RTL/core/exu_lsu.v(69)
  wire \u_EXU_LSU/mux10_b2_sel_is_2_o ;
  wire \u_EXU_LSU/mux11_b0_sel_is_2_o ;
  wire \u_EXU_LSU/mux14_b1_sel_is_0_o ;
  wire \u_EXU_LSU/mux16_b3_sel_is_2_o ;
  wire \u_EXU_LSU/mux27_b16_sel_is_1_o ;
  wire \u_EXU_LSU/mux32_b0_sel_is_0_o ;
  wire \u_EXU_LSU/n1 ;
  wire \u_EXU_LSU/n155_lutinv ;
  wire \u_EXU_LSU/n157_lutinv ;
  wire \u_EXU_LSU/n18_lutinv ;
  wire \u_EXU_LSU/n20_lutinv ;
  wire \u_EXU_LSU/n23 ;
  wire \u_EXU_LSU/n25 ;
  wire \u_EXU_LSU/n26 ;
  wire \u_EXU_LSU/n30 ;
  wire \u_EXU_LSU/n57 ;
  wire \u_EXU_LSU/n75 ;
  wire \u_EXU_LSU/n8 ;
  wire \u_EXU_LSU/n80 ;
  wire \u_EXU_LSU/working ;  // ../RTL/core/exu_lsu.v(91)

  assign o_csridx[11] = i_csridx[11];
  assign o_csridx[10] = i_csridx[10];
  assign o_csridx[9] = i_csridx[9];
  assign o_csridx[8] = i_csridx[8];
  assign o_csridx[7] = i_csridx[7];
  assign o_csridx[6] = i_csridx[6];
  assign o_csridx[5] = i_csridx[5];
  assign o_csridx[4] = i_csridx[4];
  assign o_csridx[3] = i_csridx[3];
  assign o_csridx[2] = i_csridx[2];
  assign o_csridx[1] = i_csridx[1];
  assign o_csridx[0] = i_csridx[0];
  assign o_rdidx0[4] = i_rdidx[4];
  assign o_rdidx0[3] = i_rdidx[3];
  assign o_rdidx0[2] = i_rdidx[2];
  assign o_rdidx0[1] = i_rdidx[1];
  assign o_rdidx0[0] = i_rdidx[0];
  assign o_exu_rdwen0 = i_rdwen;
  assign o_exu_rdidx0[4] = i_rdidx[4];
  assign o_exu_rdidx0[3] = i_rdidx[3];
  assign o_exu_rdidx0[2] = i_rdidx[2];
  assign o_exu_rdidx0[1] = i_rdidx[1];
  assign o_exu_rdidx0[0] = i_rdidx[0];
  assign o_exu_rdidx2[4] = o_rdidx2[4];
  assign o_exu_rdidx2[3] = o_rdidx2[3];
  assign o_exu_rdidx2[2] = o_rdidx2[2];
  assign o_exu_rdidx2[1] = o_rdidx2[1];
  assign o_exu_rdidx2[0] = o_rdidx2[0];
  assign o_ribm_addr[1] = 1'b0;
  assign o_ribm_addr[0] = 1'b0;
  assign o_ribm_rdy = i_ribm_rsp;
  AL_MAP_LUT5 #(
    .EQN("(B*(~A*~((~E*C))*~(D)+~A*(~E*C)*~(D)+~(~A)*(~E*C)*D+~A*(~E*C)*D))"),
    .INIT(32'h0044c044))
    _al_u1000 (
    .a(_al_u999_o),
    .b(_al_u965_o),
    .c(i_exu_op1[31]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(\u_EXU_ALU/n46_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1001 (
    .a(_al_u998_o),
    .b(_al_u911_o),
    .c(\u_EXU_ALU/n46_lutinv ),
    .d(_al_u917_o),
    .e(i_decinfo[3]),
    .o(\u_EXU_ALU/alu_srl [29]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1002 (
    .a(_al_u946_o),
    .b(i_exu_op2[30]),
    .c(i_exu_op2[29]),
    .o(_al_u1002_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1003 (
    .a(i_exu_op2[22]),
    .b(i_exu_op2[21]),
    .o(_al_u1003_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1004 (
    .a(_al_u1003_o),
    .b(i_exu_op2[19]),
    .c(i_exu_op2[18]),
    .d(i_exu_op2[17]),
    .e(i_exu_op2[16]),
    .o(_al_u1004_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1005 (
    .a(i_exu_op2[31]),
    .b(i_exu_op2[28]),
    .c(i_exu_op2[23]),
    .d(i_exu_op2[20]),
    .o(_al_u1005_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1006 (
    .a(_al_u1002_o),
    .b(_al_u1004_o),
    .c(_al_u937_o),
    .d(_al_u938_o),
    .e(_al_u1005_o),
    .o(_al_u1006_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1007 (
    .a(i_exu_op2[1]),
    .b(i_exu_op2[0]),
    .o(_al_u1007_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*~A))"),
    .INIT(16'hf0b0))
    _al_u1008 (
    .a(_al_u1007_o),
    .b(_al_u965_o),
    .c(i_exu_op1[31]),
    .d(i_exu_op2[4]),
    .o(\u_EXU_ALU/n235_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*~(E*D*C))"),
    .INIT(32'h02222222))
    _al_u1009 (
    .a(_al_u996_o),
    .b(\u_EXU_ALU/alu_srl [29]),
    .c(_al_u1006_o),
    .d(\u_EXU_ALU/n235_lutinv ),
    .e(i_decinfo[4]),
    .o(_al_u1009_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u1010 (
    .a(i_exu_op1[1]),
    .b(i_exu_op1[0]),
    .c(i_exu_op2[1]),
    .d(i_exu_op2[0]),
    .o(\u_EXU_ALU/n351_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haa33aa0f))
    _al_u1011 (
    .a(\u_EXU_ALU/n351_lutinv ),
    .b(_al_u903_o),
    .c(_al_u905_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(\u_EXU_ALU/n379_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*~(D)+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(D)+~(~A)*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D)"),
    .INIT(32'h0faa33aa))
    _al_u1012 (
    .a(_al_u899_o),
    .b(i_exu_op1[7]),
    .c(i_exu_op1[6]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1012_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u1013 (
    .a(i_exu_op1[13]),
    .b(i_exu_op1[12]),
    .c(i_exu_op2[0]),
    .o(_al_u1013_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*~(D)+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(D)+~(~A)*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D)"),
    .INIT(32'h0faa33aa))
    _al_u1014 (
    .a(_al_u1013_o),
    .b(i_exu_op1[11]),
    .c(i_exu_op1[10]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1014_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'h55cc55f0))
    _al_u1015 (
    .a(\u_EXU_ALU/n379_lutinv ),
    .b(_al_u1012_o),
    .c(_al_u1014_o),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(_al_u1015_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u1016 (
    .a(i_exu_op1[29]),
    .b(i_exu_op1[28]),
    .c(i_exu_op2[0]),
    .o(_al_u1016_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1017 (
    .a(_al_u920_o),
    .b(_al_u1016_o),
    .c(i_exu_op2[1]),
    .d(i_exu_op2[2]),
    .o(_al_u1017_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcaf0))
    _al_u1018 (
    .a(_al_u919_o),
    .b(_al_u928_o),
    .c(_al_u1017_o),
    .d(i_exu_op2[2]),
    .o(_al_u1018_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcaf0))
    _al_u1019 (
    .a(i_exu_op1[19]),
    .b(i_exu_op1[18]),
    .c(i_exu_op2[0]),
    .d(i_exu_op2[1]),
    .o(_al_u1019_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1020 (
    .a(i_exu_op1[21]),
    .b(i_exu_op1[20]),
    .c(_al_u1019_o),
    .d(i_exu_op2[1]),
    .o(_al_u1020_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33550f55))
    _al_u1021 (
    .a(_al_u1020_o),
    .b(_al_u897_o),
    .c(_al_u926_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(\u_EXU_ALU/n363_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~(~B*~(C)*~(E)+~B*C*~(E)+~(~B)*C*E+~B*C*E)*~(A)*~(D)+~(~B*~(C)*~(E)+~B*C*~(E)+~(~B)*C*E+~B*C*E)*A*~(D)+~(~(~B*~(C)*~(E)+~B*C*~(E)+~(~B)*C*E+~B*C*E))*A*D+~(~B*~(C)*~(E)+~B*C*~(E)+~(~B)*C*E+~B*C*E)*A*D)"),
    .INIT(32'haa0faacc))
    _al_u1022 (
    .a(_al_u1015_o),
    .b(_al_u1018_o),
    .c(\u_EXU_ALU/n363_lutinv ),
    .d(i_exu_op2[4]),
    .e(i_exu_op2[3]),
    .o(_al_u1022_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1023 (
    .a(\u_EXU_ALU/u1029_sel_is_0_o ),
    .b(\u_EXU_ALU/n46_lutinv ),
    .c(i_decinfo[4]),
    .o(_al_u1023_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1024 (
    .a(bju_rdwdata[29]),
    .b(bju_rdwen),
    .c(i_csr_rdata[29]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1024_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~C*A*~(D*~B)))"),
    .INIT(32'h0000f7f5))
    _al_u1025 (
    .a(_al_u1009_o),
    .b(_al_u1022_o),
    .c(_al_u1023_o),
    .d(_al_u918_o),
    .e(_al_u1024_o),
    .o(o_rdwdata0[29]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1026 (
    .a(i_decinfo[2]),
    .b(i_exu_op2[4]),
    .o(_al_u1026_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1027 (
    .a(_al_u911_o),
    .b(_al_u915_o),
    .c(_al_u917_o),
    .d(_al_u1026_o),
    .o(_al_u1027_o));
  AL_MAP_LUT5 #(
    .EQN("(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'haa0faa33))
    _al_u1028 (
    .a(_al_u980_o),
    .b(i_exu_op1[24]),
    .c(i_exu_op1[23]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1028_o));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haaccaaf0))
    _al_u1029 (
    .a(_al_u1028_o),
    .b(_al_u985_o),
    .c(_al_u988_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1029_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcaf0))
    _al_u1030 (
    .a(i_exu_op1[14]),
    .b(i_exu_op1[13]),
    .c(i_exu_op2[0]),
    .d(i_exu_op2[1]),
    .o(_al_u1030_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1031 (
    .a(i_exu_op1[16]),
    .b(i_exu_op1[15]),
    .c(_al_u1030_o),
    .d(i_exu_op2[1]),
    .o(_al_u1031_o));
  AL_MAP_LUT5 #(
    .EQN("((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'haaf0aacc))
    _al_u1032 (
    .a(_al_u1031_o),
    .b(_al_u979_o),
    .c(_al_u982_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1032_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*~(C)*~(D)+B*C*~(D)+~(B)*C*D+B*C*D))"),
    .INIT(16'h0a22))
    _al_u1033 (
    .a(_al_u1027_o),
    .b(_al_u1029_o),
    .c(_al_u1032_o),
    .d(i_exu_op2[3]),
    .o(_al_u1033_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1034 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[28]),
    .c(i_exu_op2[28]),
    .o(\u_EXU_ALU/alu_and [28]));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(C*A))"),
    .INIT(16'h1300))
    _al_u1035 (
    .a(\u_EXU_ALU/n33 [28]),
    .b(\u_EXU_ALU/alu_and [28]),
    .c(i_decinfo[1]),
    .d(i_decinfo_grp[0]),
    .o(_al_u1035_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1036 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[28]),
    .d(i_exu_op2[28]),
    .o(_al_u1036_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u1037 (
    .a(\u_EXU_ALU/n0 [28]),
    .b(_al_u1036_o),
    .c(i_decinfo_grp[5]),
    .o(_al_u1037_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(~D*A))"),
    .INIT(16'hc040))
    _al_u1038 (
    .a(_al_u965_o),
    .b(i_decinfo[4]),
    .c(i_exu_op1[31]),
    .d(i_exu_op2[4]),
    .o(_al_u1038_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u1039 (
    .a(_al_u1035_o),
    .b(_al_u1037_o),
    .c(_al_u1038_o),
    .d(\u_EXU_ALU/n179_neg_lutinv ),
    .o(_al_u1039_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*~(D)+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(D)+~(~A)*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D)"),
    .INIT(32'h0faa33aa))
    _al_u1040 (
    .a(_al_u976_o),
    .b(i_exu_op1[10]),
    .c(i_exu_op1[9]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1040_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u1041 (
    .a(i_exu_op1[8]),
    .b(i_exu_op1[7]),
    .c(i_exu_op2[0]),
    .o(_al_u1041_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33550f55))
    _al_u1042 (
    .a(_al_u1040_o),
    .b(_al_u972_o),
    .c(_al_u1041_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(\u_EXU_ALU/n372_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u1043 (
    .a(i_exu_op1[2]),
    .b(i_exu_op1[1]),
    .c(i_exu_op2[0]),
    .o(_al_u1043_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1044 (
    .a(i_exu_op1[0]),
    .b(i_exu_op2[0]),
    .o(\u_EXU_ALU/n327_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hffaa0fcc))
    _al_u1045 (
    .a(_al_u1043_o),
    .b(_al_u971_o),
    .c(\u_EXU_ALU/n327_lutinv ),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1045_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1046 (
    .a(_al_u911_o),
    .b(_al_u915_o),
    .c(_al_u917_o),
    .d(i_decinfo[2]),
    .e(i_exu_op2[4]),
    .o(_al_u1046_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C))"),
    .INIT(16'h3a00))
    _al_u1047 (
    .a(\u_EXU_ALU/n372_lutinv ),
    .b(_al_u1045_o),
    .c(i_exu_op2[3]),
    .d(_al_u1046_o),
    .o(_al_u1047_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1048 (
    .a(i_exu_op1[31]),
    .b(i_exu_op1[30]),
    .c(i_exu_op2[0]),
    .o(_al_u1048_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1049 (
    .a(i_exu_op1[29]),
    .b(i_exu_op1[28]),
    .c(i_exu_op2[0]),
    .o(_al_u1049_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0503))
    _al_u1050 (
    .a(_al_u1048_o),
    .b(_al_u1049_o),
    .c(i_exu_op2[2]),
    .d(i_exu_op2[1]),
    .o(\u_EXU_ALU/n80_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1051 (
    .a(_al_u998_o),
    .b(_al_u911_o),
    .c(\u_EXU_ALU/n80_lutinv ),
    .d(_al_u917_o),
    .e(_al_u954_o),
    .o(_al_u1051_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1052 (
    .a(bju_rdwdata[28]),
    .b(bju_rdwen),
    .c(i_csr_rdata[28]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1052_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~D*~C*B*~A))"),
    .INIT(32'h0000fffb))
    _al_u1053 (
    .a(_al_u1033_o),
    .b(_al_u1039_o),
    .c(_al_u1047_o),
    .d(_al_u1051_o),
    .e(_al_u1052_o),
    .o(o_rdwdata0[28]));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33550f55))
    _al_u1054 (
    .a(_al_u927_o),
    .b(_al_u1013_o),
    .c(_al_u897_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(\u_EXU_ALU/n365_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'h55f055cc))
    _al_u1055 (
    .a(\u_EXU_ALU/n365_lutinv ),
    .b(_al_u921_o),
    .c(_al_u929_o),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(_al_u1055_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1056 (
    .a(_al_u899_o),
    .b(_al_u900_o),
    .c(i_exu_op2[1]),
    .o(_al_u1056_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1057 (
    .a(i_decinfo[2]),
    .b(i_exu_op2[3]),
    .o(_al_u1057_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*C*~(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E))"),
    .INIT(32'h00500030))
    _al_u1058 (
    .a(_al_u902_o),
    .b(_al_u903_o),
    .c(_al_u1057_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1058_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u1059 (
    .a(i_decinfo[2]),
    .b(i_exu_op2[3]),
    .o(_al_u1059_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(D*~(A*~(C)*~(E)+A*C*~(E)+~(A)*C*E+A*C*E)))"),
    .INIT(32'h30332233))
    _al_u1060 (
    .a(_al_u1056_o),
    .b(_al_u1058_o),
    .c(_al_u906_o),
    .d(_al_u1059_o),
    .e(i_exu_op2[2]),
    .o(_al_u1060_o));
  AL_MAP_LUT5 #(
    .EQN("(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haa33aa0f))
    _al_u1061 (
    .a(_al_u999_o),
    .b(i_exu_op1[28]),
    .c(i_exu_op1[27]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1061_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u1062 (
    .a(i_exu_op1[31]),
    .b(i_exu_op2[1]),
    .c(i_exu_op2[0]),
    .o(\u_EXU_ALU/n110_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D))"),
    .INIT(16'hc050))
    _al_u1063 (
    .a(_al_u1061_o),
    .b(\u_EXU_ALU/n110_lutinv ),
    .c(_al_u954_o),
    .d(i_exu_op2[2]),
    .o(_al_u1063_o));
  AL_MAP_LUT5 #(
    .EQN("((~C*~(D*~A))*~(B)*~(E)+(~C*~(D*~A))*B*~(E)+~((~C*~(D*~A)))*B*E+(~C*~(D*~A))*B*E)"),
    .INIT(32'hcccc0a0f))
    _al_u1064 (
    .a(_al_u1055_o),
    .b(_al_u1060_o),
    .c(_al_u1063_o),
    .d(i_decinfo[2]),
    .e(i_exu_op2[4]),
    .o(_al_u1064_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1065 (
    .a(_al_u937_o),
    .b(_al_u938_o),
    .c(_al_u940_o),
    .d(_al_u941_o),
    .e(_al_u942_o),
    .o(_al_u1065_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1066 (
    .a(_al_u1065_o),
    .b(_al_u961_o),
    .o(_al_u1066_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D*B)*~(C*A))"),
    .INIT(32'h135f5f5f))
    _al_u1067 (
    .a(\u_EXU_ALU/n33 [27]),
    .b(i_decinfo[6]),
    .c(i_decinfo[1]),
    .d(i_exu_op1[27]),
    .e(i_exu_op2[27]),
    .o(_al_u1067_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1068 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[27]),
    .d(i_exu_op2[27]),
    .o(_al_u1068_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~C*A*~(D*B))"),
    .INIT(32'h020a0000))
    _al_u1069 (
    .a(_al_u1067_o),
    .b(\u_EXU_ALU/n0 [27]),
    .c(_al_u1068_o),
    .d(i_decinfo_grp[5]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1069_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1070 (
    .a(_al_u924_o),
    .b(i_exu_op1[31]),
    .o(\u_EXU_ALU/n229_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(~D*~C))"),
    .INIT(16'h8880))
    _al_u1071 (
    .a(i_exu_op1[31]),
    .b(i_exu_op2[2]),
    .c(i_exu_op2[1]),
    .d(i_exu_op2[0]),
    .o(\u_EXU_ALU/n256_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(B*~(A*~(~D*~C)))"),
    .INIT(16'h444c))
    _al_u1072 (
    .a(_al_u1066_o),
    .b(_al_u1069_o),
    .c(\u_EXU_ALU/n229_lutinv ),
    .d(\u_EXU_ALU/n256_lutinv ),
    .o(_al_u1072_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1073 (
    .a(bju_rdwdata[27]),
    .b(bju_rdwen),
    .c(i_csr_rdata[27]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1073_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(C*~A)))"),
    .INIT(16'h0073))
    _al_u1074 (
    .a(_al_u1064_o),
    .b(_al_u1072_o),
    .c(\u_EXU_ALU/n281_neg_lutinv ),
    .d(_al_u1073_o),
    .o(o_rdwdata0[27]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u1075 (
    .a(\u_EXU_ALU/n0 [26]),
    .b(i_decinfo_grp[5]),
    .c(i_decinfo_grp[0]),
    .o(_al_u1075_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1076 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[26]),
    .d(i_exu_op2[26]),
    .o(_al_u1076_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1077 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[26]),
    .c(i_exu_op2[26]),
    .o(\u_EXU_ALU/alu_and [26]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*A*~(E*B))"),
    .INIT(32'h0002000a))
    _al_u1078 (
    .a(_al_u1075_o),
    .b(\u_EXU_ALU/n33 [26]),
    .c(_al_u1076_o),
    .d(\u_EXU_ALU/alu_and [26]),
    .e(i_decinfo[1]),
    .o(_al_u1078_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u1079 (
    .a(_al_u981_o),
    .b(_al_u986_o),
    .c(i_exu_op2[3]),
    .d(i_exu_op2[2]),
    .o(_al_u1079_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u1080 (
    .a(i_exu_op1[14]),
    .b(i_exu_op1[13]),
    .c(i_exu_op2[0]),
    .o(_al_u1080_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*~(D)+A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(D)+~(A)*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D+A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D)"),
    .INIT(32'h0f553355))
    _al_u1081 (
    .a(_al_u983_o),
    .b(_al_u1080_o),
    .c(_al_u976_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(\u_EXU_ALU/n366_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~C*A*~(E*~D)))"),
    .INIT(32'hc4ccc4c4))
    _al_u1082 (
    .a(_al_u1027_o),
    .b(_al_u1078_o),
    .c(_al_u1079_o),
    .d(\u_EXU_ALU/n366_lutinv ),
    .e(i_exu_op2[3]),
    .o(_al_u1082_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'h55cc55f0))
    _al_u1083 (
    .a(_al_u1049_o),
    .b(i_exu_op1[27]),
    .c(i_exu_op1[26]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(\u_EXU_ALU/n115_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u1084 (
    .a(\u_EXU_ALU/n115_lutinv ),
    .b(\u_EXU_ALU/n111_lutinv ),
    .c(i_exu_op2[3]),
    .d(i_exu_op2[2]),
    .o(\u_EXU_ALU/n49_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1085 (
    .a(i_exu_op1[31]),
    .b(i_exu_op2[2]),
    .c(i_exu_op2[1]),
    .o(\u_EXU_ALU/n255_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u1086 (
    .a(\u_EXU_ALU/n229_lutinv ),
    .b(\u_EXU_ALU/n255_lutinv ),
    .c(i_decinfo[4]),
    .o(_al_u1086_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~(C*B)*~(D*A)))"),
    .INIT(32'h0000eac0))
    _al_u1087 (
    .a(\u_EXU_ALU/n179_neg_lutinv ),
    .b(\u_EXU_ALU/u1029_sel_is_0_o ),
    .c(\u_EXU_ALU/n49_lutinv ),
    .d(_al_u1086_o),
    .e(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .o(_al_u1087_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*~(D)+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(D)+~(~A)*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D)"),
    .INIT(32'h0faa33aa))
    _al_u1088 (
    .a(_al_u972_o),
    .b(i_exu_op1[4]),
    .c(i_exu_op1[3]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1088_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hffaaf0cc))
    _al_u1089 (
    .a(_al_u1088_o),
    .b(_al_u975_o),
    .c(_al_u970_o),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(_al_u1089_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1090 (
    .a(bju_rdwdata[26]),
    .b(bju_rdwen),
    .c(i_csr_rdata[26]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1090_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~B*A*~(~D*C)))"),
    .INIT(32'h0000ddfd))
    _al_u1091 (
    .a(_al_u1082_o),
    .b(_al_u1087_o),
    .c(_al_u1046_o),
    .d(_al_u1089_o),
    .e(_al_u1090_o),
    .o(o_rdwdata0[26]));
  AL_MAP_LUT5 #(
    .EQN("(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'haa0faa33))
    _al_u1092 (
    .a(_al_u897_o),
    .b(i_exu_op1[17]),
    .c(i_exu_op1[16]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1092_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1093 (
    .a(_al_u1014_o),
    .b(_al_u1092_o),
    .c(_al_u930_o),
    .d(i_exu_op2[2]),
    .o(_al_u1093_o));
  AL_MAP_LUT5 #(
    .EQN("((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'haaf0aacc))
    _al_u1094 (
    .a(_al_u1020_o),
    .b(_al_u919_o),
    .c(_al_u928_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1094_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*~B)))"),
    .INIT(16'hba00))
    _al_u1095 (
    .a(_al_u1093_o),
    .b(_al_u1094_o),
    .c(_al_u924_o),
    .d(i_decinfo[2]),
    .o(_al_u1095_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff33550f))
    _al_u1096 (
    .a(i_exu_op1[31]),
    .b(i_exu_op1[30]),
    .c(i_exu_op1[29]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1096_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1097 (
    .a(i_exu_op1[28]),
    .b(i_exu_op1[27]),
    .c(i_exu_op2[0]),
    .o(_al_u1097_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1098 (
    .a(i_exu_op1[26]),
    .b(i_exu_op1[25]),
    .c(i_exu_op2[0]),
    .o(_al_u1098_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'h5533550f))
    _al_u1099 (
    .a(_al_u1096_o),
    .b(_al_u1097_o),
    .c(_al_u1098_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(\u_EXU_ALU/n83_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1100 (
    .a(\u_EXU_ALU/n83_lutinv ),
    .b(_al_u954_o),
    .c(i_exu_op2[4]),
    .o(_al_u1100_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u1101 (
    .a(\u_EXU_ALU/n351_lutinv ),
    .b(_al_u1057_o),
    .c(i_exu_op2[2]),
    .o(_al_u1101_o));
  AL_MAP_LUT5 #(
    .EQN("(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'haa0faa33))
    _al_u1102 (
    .a(_al_u903_o),
    .b(i_exu_op1[5]),
    .c(i_exu_op1[4]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1102_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)))"),
    .INIT(32'h44555055))
    _al_u1103 (
    .a(_al_u1101_o),
    .b(_al_u1102_o),
    .c(_al_u1012_o),
    .d(_al_u1059_o),
    .e(i_exu_op2[2]),
    .o(_al_u1103_o));
  AL_MAP_LUT5 #(
    .EQN("(D*~(~B*~A*~(E*~C)))"),
    .INIT(32'hef00ee00))
    _al_u1104 (
    .a(_al_u1095_o),
    .b(_al_u1100_o),
    .c(_al_u1103_o),
    .d(\u_EXU_ALU/n281_neg_lutinv ),
    .e(i_exu_op2[4]),
    .o(_al_u1104_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D*B)*~(C*A))"),
    .INIT(32'h135f5f5f))
    _al_u1105 (
    .a(\u_EXU_ALU/n33 [25]),
    .b(i_decinfo[6]),
    .c(i_decinfo[1]),
    .d(i_exu_op1[25]),
    .e(i_exu_op2[25]),
    .o(_al_u1105_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1106 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[25]),
    .d(i_exu_op2[25]),
    .o(_al_u1106_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u1107 (
    .a(_al_u1105_o),
    .b(\u_EXU_ALU/n0 [25]),
    .c(_al_u1106_o),
    .d(i_decinfo_grp[5]),
    .o(_al_u1107_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1108 (
    .a(i_exu_op1[31]),
    .b(i_exu_op2[3]),
    .o(_al_u1108_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u1109 (
    .a(\u_EXU_ALU/n255_lutinv ),
    .b(_al_u1108_o),
    .c(i_exu_op2[0]),
    .o(_al_u1109_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    _al_u1110 (
    .a(_al_u1109_o),
    .b(i_exu_op1[31]),
    .c(i_exu_op2[4]),
    .o(_al_u1110_o));
  AL_MAP_LUT4 #(
    .EQN("(D*B*~(~C*A))"),
    .INIT(16'hc400))
    _al_u1111 (
    .a(_al_u1066_o),
    .b(_al_u1107_o),
    .c(_al_u1110_o),
    .d(i_decinfo_grp[0]),
    .o(_al_u1111_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u1112 (
    .a(bju_rdwdata[25]),
    .b(bju_rdwen),
    .c(i_csr_rdata[25]),
    .d(i_decinfo_grp[4]),
    .o(_al_u1112_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*C)*~(B*~A))"),
    .INIT(16'hbb0b))
    _al_u1113 (
    .a(_al_u1104_o),
    .b(_al_u1111_o),
    .c(_al_u1112_o),
    .d(i_decinfo_grp[0]),
    .o(o_rdwdata0[25]));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*~(D)+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(D)+~(~A)*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D)"),
    .INIT(32'h0faa33aa))
    _al_u1114 (
    .a(_al_u971_o),
    .b(i_exu_op1[2]),
    .c(i_exu_op1[1]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1114_o));
  AL_MAP_LUT5 #(
    .EQN("(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'haa0faa33))
    _al_u1115 (
    .a(_al_u972_o),
    .b(i_exu_op1[8]),
    .c(i_exu_op1[7]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1115_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u1116 (
    .a(i_exu_op1[0]),
    .b(i_exu_op2[1]),
    .c(i_exu_op2[0]),
    .o(\u_EXU_ALU/n352_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hffaa0fcc))
    _al_u1117 (
    .a(_al_u1114_o),
    .b(_al_u1115_o),
    .c(\u_EXU_ALU/n352_lutinv ),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(_al_u1117_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D*B)*~(~C*A))"),
    .INIT(32'h31f5f5f5))
    _al_u1118 (
    .a(_al_u1046_o),
    .b(_al_u1006_o),
    .c(_al_u1117_o),
    .d(\u_EXU_ALU/n229_lutinv ),
    .e(i_decinfo[4]),
    .o(_al_u1118_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*~(D)+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(D)+~(~A)*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D)"),
    .INIT(32'h0faa33aa))
    _al_u1119 (
    .a(_al_u979_o),
    .b(i_exu_op1[18]),
    .c(i_exu_op1[17]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1119_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u1120 (
    .a(_al_u1028_o),
    .b(_al_u1119_o),
    .c(i_exu_op2[3]),
    .d(i_exu_op2[2]),
    .o(_al_u1120_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'hccaaf0aa))
    _al_u1121 (
    .a(_al_u1031_o),
    .b(_al_u974_o),
    .c(_al_u976_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1121_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u1122 (
    .a(_al_u1027_o),
    .b(_al_u1120_o),
    .c(_al_u1121_o),
    .d(i_exu_op2[3]),
    .o(_al_u1122_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1123 (
    .a(i_exu_op1[27]),
    .b(i_exu_op1[26]),
    .c(i_exu_op2[0]),
    .o(_al_u1123_o));
  AL_MAP_LUT5 #(
    .EQN("(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haa33aa0f))
    _al_u1124 (
    .a(_al_u1123_o),
    .b(i_exu_op1[25]),
    .c(i_exu_op1[24]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1124_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33550f55))
    _al_u1125 (
    .a(_al_u1124_o),
    .b(_al_u1048_o),
    .c(_al_u1049_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(\u_EXU_ALU/n84_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1126 (
    .a(\u_EXU_ALU/u1029_sel_is_0_o ),
    .b(\u_EXU_ALU/n84_lutinv ),
    .c(_al_u954_o),
    .o(_al_u1126_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(C*B)*~(D*A))"),
    .INIT(32'h153f0000))
    _al_u1127 (
    .a(\u_EXU_ALU/n0 [24]),
    .b(\u_EXU_ALU/n33 [24]),
    .c(i_decinfo[1]),
    .d(i_decinfo_grp[5]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1127_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h155f))
    _al_u1128 (
    .a(i_decinfo[7]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[24]),
    .d(i_exu_op2[24]),
    .o(_al_u1128_o));
  AL_MAP_LUT5 #(
    .EQN("(B*A*~(C*(E@D)))"),
    .INIT(32'h88080888))
    _al_u1129 (
    .a(_al_u1127_o),
    .b(_al_u1128_o),
    .c(i_decinfo[5]),
    .d(i_exu_op1[24]),
    .e(i_exu_op2[24]),
    .o(_al_u1129_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1130 (
    .a(bju_rdwdata[24]),
    .b(bju_rdwen),
    .c(i_csr_rdata[24]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1130_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*~C*~B*A))"),
    .INIT(32'h0000fdff))
    _al_u1131 (
    .a(_al_u1118_o),
    .b(_al_u1122_o),
    .c(_al_u1126_o),
    .d(_al_u1129_o),
    .e(_al_u1130_o),
    .o(o_rdwdata0[24]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1132 (
    .a(i_exu_op1[24]),
    .b(i_exu_op1[23]),
    .c(i_exu_op2[0]),
    .o(_al_u1132_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1133 (
    .a(_al_u1098_o),
    .b(_al_u1132_o),
    .c(i_exu_op2[1]),
    .o(_al_u1133_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u1134 (
    .a(i_decinfo[4]),
    .b(i_decinfo[3]),
    .c(i_exu_op2[3]),
    .o(_al_u1134_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1135 (
    .a(\u_EXU_ALU/n77_lutinv ),
    .b(_al_u1134_o),
    .o(_al_u1135_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(D*~(A*~(C)*~(E)+A*C*~(E)+~(A)*C*E+A*C*E)))"),
    .INIT(32'h30332233))
    _al_u1136 (
    .a(_al_u1133_o),
    .b(_al_u1135_o),
    .c(_al_u1061_o),
    .d(_al_u954_o),
    .e(i_exu_op2[2]),
    .o(_al_u1136_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1137 (
    .a(_al_u927_o),
    .b(_al_u929_o),
    .c(_al_u1059_o),
    .d(i_exu_op2[2]),
    .o(_al_u1137_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~B*A*~(D*C))"),
    .INIT(32'h00000222))
    _al_u1138 (
    .a(_al_u1136_o),
    .b(_al_u1137_o),
    .c(\u_EXU_ALU/n369_lutinv ),
    .d(_al_u1057_o),
    .e(i_exu_op2[4]),
    .o(_al_u1138_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1139 (
    .a(_al_u904_o),
    .b(_al_u906_o),
    .c(_al_u1059_o),
    .d(i_exu_op2[2]),
    .o(_al_u1139_o));
  AL_MAP_LUT5 #(
    .EQN("(D*C*B*~(E*~A))"),
    .INIT(32'h8000c000))
    _al_u1140 (
    .a(_al_u1139_o),
    .b(_al_u911_o),
    .c(_al_u915_o),
    .d(_al_u917_o),
    .e(i_exu_op2[4]),
    .o(_al_u1140_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1141 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[23]),
    .d(i_exu_op2[23]),
    .o(_al_u1141_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u1142 (
    .a(\u_EXU_ALU/n0 [23]),
    .b(_al_u1141_o),
    .c(i_decinfo_grp[5]),
    .o(_al_u1142_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1143 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[23]),
    .c(i_exu_op2[23]),
    .o(\u_EXU_ALU/alu_and [23]));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(C*A))"),
    .INIT(16'h1300))
    _al_u1144 (
    .a(\u_EXU_ALU/n33 [23]),
    .b(\u_EXU_ALU/alu_and [23]),
    .c(i_decinfo[1]),
    .d(i_decinfo_grp[0]),
    .o(_al_u1144_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~C*~(D*~(~E*A))))"),
    .INIT(32'hccc0c4c0))
    _al_u1145 (
    .a(_al_u948_o),
    .b(i_exu_op1[31]),
    .c(i_exu_op2[4]),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[0]),
    .o(\u_EXU_ALU/n228_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(C*B*~(E*D*A))"),
    .INIT(32'h40c0c0c0))
    _al_u1146 (
    .a(_al_u1065_o),
    .b(_al_u1142_o),
    .c(_al_u1144_o),
    .d(_al_u961_o),
    .e(\u_EXU_ALU/n228_lutinv ),
    .o(_al_u1146_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1147 (
    .a(bju_rdwdata[23]),
    .b(bju_rdwen),
    .c(i_csr_rdata[23]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1147_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(B*~A)))"),
    .INIT(16'h004f))
    _al_u1148 (
    .a(_al_u1138_o),
    .b(_al_u1140_o),
    .c(_al_u1146_o),
    .d(_al_u1147_o),
    .o(o_rdwdata0[23]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u1149 (
    .a(\u_EXU_ALU/n0 [22]),
    .b(i_decinfo_grp[5]),
    .c(i_decinfo_grp[0]),
    .o(_al_u1149_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h155f))
    _al_u1150 (
    .a(i_decinfo[7]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[22]),
    .d(i_exu_op2[22]),
    .o(_al_u1150_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u1151 (
    .a(i_decinfo[5]),
    .b(i_exu_op1[22]),
    .c(i_exu_op2[22]),
    .o(\u_EXU_ALU/alu_xor [22]));
  AL_MAP_LUT5 #(
    .EQN("(~D*C*A*~(E*B))"),
    .INIT(32'h002000a0))
    _al_u1152 (
    .a(_al_u1149_o),
    .b(\u_EXU_ALU/n33 [22]),
    .c(_al_u1150_o),
    .d(\u_EXU_ALU/alu_xor [22]),
    .e(i_decinfo[1]),
    .o(_al_u1152_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~C*~(D*~A)))"),
    .INIT(16'hc4c0))
    _al_u1153 (
    .a(_al_u948_o),
    .b(i_exu_op1[31]),
    .c(i_exu_op2[4]),
    .d(i_exu_op2[3]),
    .o(\u_EXU_ALU/n227_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u1154 (
    .a(_al_u1152_o),
    .b(_al_u1065_o),
    .c(_al_u961_o),
    .d(\u_EXU_ALU/n227_lutinv ),
    .o(_al_u1154_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33550f55))
    _al_u1155 (
    .a(_al_u977_o),
    .b(_al_u1041_o),
    .c(_al_u974_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(\u_EXU_ALU/n370_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(C*(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'h003f005f))
    _al_u1156 (
    .a(\u_EXU_ALU/n362_lutinv ),
    .b(\u_EXU_ALU/n370_lutinv ),
    .c(i_decinfo[2]),
    .d(i_exu_op2[4]),
    .e(i_exu_op2[3]),
    .o(_al_u1156_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h3050))
    _al_u1157 (
    .a(_al_u1088_o),
    .b(_al_u970_o),
    .c(_al_u1059_o),
    .d(i_exu_op2[2]),
    .o(_al_u1157_o));
  AL_MAP_LUT5 #(
    .EQN("(D*C*B*~(E*~A))"),
    .INIT(32'h8000c000))
    _al_u1158 (
    .a(_al_u1157_o),
    .b(_al_u911_o),
    .c(_al_u915_o),
    .d(_al_u917_o),
    .e(i_exu_op2[4]),
    .o(_al_u1158_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(~B*~A))"),
    .INIT(16'h00e0))
    _al_u1159 (
    .a(i_decinfo[4]),
    .b(i_decinfo[3]),
    .c(i_exu_op2[3]),
    .d(i_exu_op2[2]),
    .o(_al_u1159_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1160 (
    .a(\u_EXU_ALU/n111_lutinv ),
    .b(_al_u1159_o),
    .o(_al_u1160_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1161 (
    .a(i_exu_op1[23]),
    .b(i_exu_op1[22]),
    .c(i_exu_op2[0]),
    .o(_al_u1161_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(~A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33aa0faa))
    _al_u1162 (
    .a(_al_u1161_o),
    .b(i_exu_op1[25]),
    .c(i_exu_op1[24]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1162_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E)))"),
    .INIT(32'h11555055))
    _al_u1163 (
    .a(_al_u1160_o),
    .b(\u_EXU_ALU/n115_lutinv ),
    .c(_al_u1162_o),
    .d(_al_u954_o),
    .e(i_exu_op2[2]),
    .o(_al_u1163_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1164 (
    .a(bju_rdwdata[22]),
    .b(bju_rdwen),
    .c(i_csr_rdata[22]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1164_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(A*~(C*~(D*B))))"),
    .INIT(32'h000075f5))
    _al_u1165 (
    .a(_al_u1154_o),
    .b(_al_u1156_o),
    .c(_al_u1158_o),
    .d(_al_u1163_o),
    .e(_al_u1164_o),
    .o(o_rdwdata0[22]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1166 (
    .a(_al_u1012_o),
    .b(_al_u1014_o),
    .c(i_exu_op2[2]),
    .o(\u_EXU_ALU/n371_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(C*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'h005f003f))
    _al_u1167 (
    .a(\u_EXU_ALU/n371_lutinv ),
    .b(\u_EXU_ALU/n363_lutinv ),
    .c(i_decinfo[2]),
    .d(i_exu_op2[4]),
    .e(i_exu_op2[3]),
    .o(_al_u1167_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D))"),
    .INIT(16'hc050))
    _al_u1168 (
    .a(_al_u1102_o),
    .b(\u_EXU_ALU/n351_lutinv ),
    .c(_al_u1059_o),
    .d(i_exu_op2[2]),
    .o(_al_u1168_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u1169 (
    .a(\u_EXU_ALU/n281_neg_lutinv ),
    .b(_al_u1168_o),
    .c(i_exu_op2[4]),
    .o(_al_u1169_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u1170 (
    .a(i_decinfo[5]),
    .b(i_exu_op1[21]),
    .c(i_exu_op2[21]),
    .o(\u_EXU_ALU/alu_xor [21]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1171 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[21]),
    .c(i_exu_op2[21]),
    .o(\u_EXU_ALU/alu_and [21]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D*A))"),
    .INIT(16'h0103))
    _al_u1172 (
    .a(\u_EXU_ALU/n0 [21]),
    .b(\u_EXU_ALU/alu_xor [21]),
    .c(\u_EXU_ALU/alu_and [21]),
    .d(i_decinfo_grp[5]),
    .o(_al_u1172_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u1173 (
    .a(i_decinfo[7]),
    .b(i_exu_op1[21]),
    .c(i_exu_op2[21]),
    .o(\u_EXU_ALU/alu_or [21]));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(C*A))"),
    .INIT(16'h1300))
    _al_u1174 (
    .a(\u_EXU_ALU/n33 [21]),
    .b(\u_EXU_ALU/alu_or [21]),
    .c(i_decinfo[1]),
    .d(i_decinfo_grp[0]),
    .o(_al_u1174_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~C*~(D*~(~E*~A))))"),
    .INIT(32'hccc0c8c0))
    _al_u1175 (
    .a(_al_u1007_o),
    .b(i_exu_op1[31]),
    .c(i_exu_op2[4]),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(\u_EXU_ALU/n226_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(C*B*~(E*D*A))"),
    .INIT(32'h40c0c0c0))
    _al_u1176 (
    .a(_al_u1065_o),
    .b(_al_u1172_o),
    .c(_al_u1174_o),
    .d(_al_u961_o),
    .e(\u_EXU_ALU/n226_lutinv ),
    .o(_al_u1176_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1177 (
    .a(_al_u1096_o),
    .b(_al_u1159_o),
    .o(_al_u1177_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1178 (
    .a(i_exu_op1[22]),
    .b(i_exu_op1[21]),
    .c(i_exu_op2[0]),
    .o(_al_u1178_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1179 (
    .a(_al_u1132_o),
    .b(_al_u1178_o),
    .c(i_exu_op2[1]),
    .o(_al_u1179_o));
  AL_MAP_LUT5 #(
    .EQN("(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haa33aa0f))
    _al_u1180 (
    .a(_al_u1097_o),
    .b(i_exu_op1[26]),
    .c(i_exu_op1[25]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1180_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)))"),
    .INIT(32'h50554455))
    _al_u1181 (
    .a(_al_u1177_o),
    .b(_al_u1179_o),
    .c(_al_u1180_o),
    .d(_al_u954_o),
    .e(i_exu_op2[2]),
    .o(_al_u1181_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1182 (
    .a(bju_rdwdata[21]),
    .b(bju_rdwen),
    .c(i_csr_rdata[21]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1182_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*~(B*~(D*A))))"),
    .INIT(32'h00004fcf))
    _al_u1183 (
    .a(_al_u1167_o),
    .b(_al_u1169_o),
    .c(_al_u1176_o),
    .d(_al_u1181_o),
    .e(_al_u1182_o),
    .o(o_rdwdata0[21]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D))"),
    .INIT(16'h220a))
    _al_u1184 (
    .a(_al_u1159_o),
    .b(_al_u1048_o),
    .c(_al_u1049_o),
    .d(i_exu_op2[1]),
    .o(_al_u1184_o));
  AL_MAP_LUT5 #(
    .EQN("(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haa33aa0f))
    _al_u1185 (
    .a(_al_u1161_o),
    .b(i_exu_op1[21]),
    .c(i_exu_op1[20]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1185_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)))"),
    .INIT(32'h44555055))
    _al_u1186 (
    .a(_al_u1184_o),
    .b(_al_u1124_o),
    .c(_al_u1185_o),
    .d(_al_u954_o),
    .e(i_exu_op2[2]),
    .o(_al_u1186_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'hf050f030))
    _al_u1187 (
    .a(_al_u1031_o),
    .b(_al_u1119_o),
    .c(i_decinfo[2]),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(_al_u1187_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*A*~(B*~(E*~C)))"),
    .INIT(32'h002a0022))
    _al_u1188 (
    .a(_al_u1186_o),
    .b(_al_u1187_o),
    .c(\u_EXU_ALU/n372_lutinv ),
    .d(i_exu_op2[4]),
    .e(i_exu_op2[3]),
    .o(_al_u1188_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1189 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[20]),
    .d(i_exu_op2[20]),
    .o(_al_u1189_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1190 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[20]),
    .c(i_exu_op2[20]),
    .o(\u_EXU_ALU/alu_and [20]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~B*~A*~(E*C))"),
    .INIT(32'h00010011))
    _al_u1191 (
    .a(alu2lsu_result[20]),
    .b(_al_u1189_o),
    .c(\u_EXU_ALU/n33 [20]),
    .d(\u_EXU_ALU/alu_and [20]),
    .e(i_decinfo[1]),
    .o(_al_u1191_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1192 (
    .a(i_exu_op1[31]),
    .b(i_exu_op2[3]),
    .c(i_exu_op2[2]),
    .o(\u_EXU_ALU/n241_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1193 (
    .a(i_exu_op1[31]),
    .b(i_exu_op2[4]),
    .o(_al_u1193_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(C*B*~(~E*~D)))"),
    .INIT(32'h2a2a2aaa))
    _al_u1194 (
    .a(_al_u1191_o),
    .b(_al_u1065_o),
    .c(_al_u961_o),
    .d(\u_EXU_ALU/n241_lutinv ),
    .e(_al_u1193_o),
    .o(_al_u1194_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(~A*~(B)*~(D)+~A*B*~(D)+~(~A)*B*D+~A*B*D))"),
    .INIT(16'hc050))
    _al_u1195 (
    .a(_al_u1114_o),
    .b(\u_EXU_ALU/n352_lutinv ),
    .c(_al_u1059_o),
    .d(i_exu_op2[2]),
    .o(_al_u1195_o));
  AL_MAP_LUT5 #(
    .EQN("(D*C*B*~(E*~A))"),
    .INIT(32'h8000c000))
    _al_u1196 (
    .a(_al_u1195_o),
    .b(_al_u911_o),
    .c(_al_u915_o),
    .d(_al_u917_o),
    .e(i_exu_op2[4]),
    .o(_al_u1196_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u1197 (
    .a(bju_rdwdata[20]),
    .b(bju_rdwen),
    .c(i_csr_rdata[20]),
    .d(i_decinfo_grp[4]),
    .o(_al_u1197_o));
  AL_MAP_LUT5 #(
    .EQN("~(D*~((B*~(C*~A)))*~(E)+D*(B*~(C*~A))*~(E)+~(D)*(B*~(C*~A))*E+D*(B*~(C*~A))*E)"),
    .INIT(32'h737300ff))
    _al_u1198 (
    .a(_al_u1188_o),
    .b(_al_u1194_o),
    .c(_al_u1196_o),
    .d(_al_u1197_o),
    .e(i_decinfo_grp[0]),
    .o(o_rdwdata0[20]));
  AL_MAP_LUT5 #(
    .EQN("~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'h55cc55f0))
    _al_u1199 (
    .a(\u_EXU_ALU/n110_lutinv ),
    .b(_al_u999_o),
    .c(_al_u1097_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1199_o));
  AL_MAP_LUT5 #(
    .EQN("(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haa33aa0f))
    _al_u1200 (
    .a(_al_u1178_o),
    .b(i_exu_op1[20]),
    .c(i_exu_op1[19]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1200_o));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haaccaaf0))
    _al_u1201 (
    .a(_al_u1199_o),
    .b(_al_u1133_o),
    .c(_al_u1200_o),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(_al_u1201_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u1202 (
    .a(_al_u1056_o),
    .b(_al_u906_o),
    .c(i_exu_op2[2]),
    .o(\u_EXU_ALU/n373_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'hf050f030))
    _al_u1203 (
    .a(_al_u898_o),
    .b(_al_u927_o),
    .c(i_decinfo[2]),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(_al_u1203_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~(E*~B)*C)*~(~D*~A))"),
    .INIT(32'h3f2a0f0a))
    _al_u1204 (
    .a(_al_u1201_o),
    .b(\u_EXU_ALU/n373_lutinv ),
    .c(_al_u1203_o),
    .d(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .e(i_exu_op2[3]),
    .o(_al_u1204_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u1205 (
    .a(\u_EXU_ALU/n0 [19]),
    .b(i_decinfo_grp[5]),
    .c(i_decinfo_grp[0]),
    .o(_al_u1205_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h155f))
    _al_u1206 (
    .a(i_decinfo[7]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[19]),
    .d(i_exu_op2[19]),
    .o(_al_u1206_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u1207 (
    .a(_al_u1205_o),
    .b(_al_u1206_o),
    .c(\u_EXU_ALU/n33 [19]),
    .d(i_decinfo[1]),
    .o(_al_u1207_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1208 (
    .a(_al_u902_o),
    .b(_al_u903_o),
    .c(_al_u965_o),
    .d(i_exu_op2[1]),
    .o(\u_EXU_ALU/n413_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1209 (
    .a(_al_u1046_o),
    .b(_al_u1207_o),
    .c(\u_EXU_ALU/n413_lutinv ),
    .o(_al_u1209_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1210 (
    .a(\u_EXU_ALU/n256_lutinv ),
    .b(_al_u930_o),
    .o(_al_u1210_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u1211 (
    .a(i_decinfo[5]),
    .b(i_exu_op1[19]),
    .c(i_exu_op2[19]),
    .o(\u_EXU_ALU/alu_xor [19]));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(E*A*~(~D*~B)))"),
    .INIT(32'h05070f0f))
    _al_u1212 (
    .a(_al_u1006_o),
    .b(_al_u1210_o),
    .c(\u_EXU_ALU/alu_xor [19]),
    .d(_al_u1193_o),
    .e(i_decinfo[4]),
    .o(_al_u1212_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1213 (
    .a(bju_rdwdata[19]),
    .b(bju_rdwen),
    .c(i_csr_rdata[19]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1213_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*B*~(D*~A)))"),
    .INIT(32'h00007f3f))
    _al_u1214 (
    .a(_al_u1204_o),
    .b(_al_u1209_o),
    .c(_al_u1212_o),
    .d(\u_EXU_ALU/u1029_sel_is_0_o ),
    .e(_al_u1213_o),
    .o(o_rdwdata0[19]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hffccaaf0))
    _al_u1215 (
    .a(_al_u1048_o),
    .b(_al_u1049_o),
    .c(_al_u1123_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1215_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1216 (
    .a(i_exu_op1[19]),
    .b(i_exu_op1[18]),
    .c(i_exu_op2[0]),
    .o(_al_u1216_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(~A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33aa0faa))
    _al_u1217 (
    .a(_al_u1216_o),
    .b(i_exu_op1[21]),
    .c(i_exu_op1[20]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1217_o));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haaccaaf0))
    _al_u1218 (
    .a(_al_u1215_o),
    .b(_al_u1162_o),
    .c(_al_u1217_o),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(_al_u1218_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~D*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'hf050f030))
    _al_u1219 (
    .a(_al_u977_o),
    .b(_al_u983_o),
    .c(i_decinfo[2]),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(_al_u1219_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33550f55))
    _al_u1220 (
    .a(_al_u975_o),
    .b(_al_u971_o),
    .c(_al_u972_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(\u_EXU_ALU/n374_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~(~(E*~C)*B)*~(~D*~A))"),
    .INIT(32'h3f2a3322))
    _al_u1221 (
    .a(_al_u1218_o),
    .b(_al_u1219_o),
    .c(\u_EXU_ALU/n374_lutinv ),
    .d(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .e(i_exu_op2[3]),
    .o(_al_u1221_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1222 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[18]),
    .c(i_exu_op2[18]),
    .o(\u_EXU_ALU/alu_and [18]));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*B)*~(E*A))"),
    .INIT(32'h0105030f))
    _al_u1223 (
    .a(\u_EXU_ALU/n0 [18]),
    .b(\u_EXU_ALU/n33 [18]),
    .c(\u_EXU_ALU/alu_and [18]),
    .d(i_decinfo[1]),
    .e(i_decinfo_grp[5]),
    .o(_al_u1223_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*A)*~(B)*~(C)+(D*A)*B*~(C)+~((D*A))*B*C+(D*A)*B*C)"),
    .INIT(16'h353f))
    _al_u1224 (
    .a(\u_EXU_ALU/n241_lutinv ),
    .b(i_exu_op1[31]),
    .c(i_exu_op2[4]),
    .d(i_exu_op2[1]),
    .o(_al_u1224_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1225 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[18]),
    .d(i_exu_op2[18]),
    .o(_al_u1225_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*B*~(~D*C*A))"),
    .INIT(32'h0000cc4c))
    _al_u1226 (
    .a(_al_u1065_o),
    .b(_al_u1223_o),
    .c(_al_u961_o),
    .d(_al_u1224_o),
    .e(_al_u1225_o),
    .o(_al_u1226_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1227 (
    .a(i_decinfo[2]),
    .b(i_exu_op2[4]),
    .o(_al_u1227_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u1228 (
    .a(_al_u970_o),
    .b(_al_u965_o),
    .c(_al_u1227_o),
    .o(_al_u1228_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D*C*B*A))"),
    .INIT(32'h7fff0000))
    _al_u1229 (
    .a(_al_u1228_o),
    .b(_al_u911_o),
    .c(_al_u915_o),
    .d(_al_u917_o),
    .e(i_decinfo_grp[0]),
    .o(_al_u1229_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1230 (
    .a(bju_rdwdata[18]),
    .b(bju_rdwen),
    .c(i_csr_rdata[18]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1230_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*B*~(D*~A)))"),
    .INIT(32'h00007f3f))
    _al_u1231 (
    .a(_al_u1221_o),
    .b(_al_u1226_o),
    .c(_al_u1229_o),
    .d(\u_EXU_ALU/u1029_sel_is_0_o ),
    .e(_al_u1230_o),
    .o(o_rdwdata0[18]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1232 (
    .a(i_exu_op1[18]),
    .b(i_exu_op1[17]),
    .c(i_exu_op2[0]),
    .o(_al_u1232_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(~A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33aa0faa))
    _al_u1233 (
    .a(_al_u1232_o),
    .b(i_exu_op1[20]),
    .c(i_exu_op1[19]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1233_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'h55cc55f0))
    _al_u1234 (
    .a(\u_EXU_ALU/n83_lutinv ),
    .b(_al_u1179_o),
    .c(_al_u1233_o),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(_al_u1234_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1235 (
    .a(_al_u1014_o),
    .b(_al_u1092_o),
    .c(_al_u1059_o),
    .d(i_exu_op2[2]),
    .o(_al_u1235_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33550f55))
    _al_u1236 (
    .a(_al_u1012_o),
    .b(_al_u903_o),
    .c(_al_u905_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(\u_EXU_ALU/n375_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*C)*~(~D*~A))"),
    .INIT(32'h03023322))
    _al_u1237 (
    .a(_al_u1234_o),
    .b(_al_u1235_o),
    .c(\u_EXU_ALU/n375_lutinv ),
    .d(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .e(_al_u1057_o),
    .o(_al_u1237_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D*B)*~(C*A))"),
    .INIT(32'h135f5f5f))
    _al_u1238 (
    .a(\u_EXU_ALU/n33 [17]),
    .b(i_decinfo[6]),
    .c(i_decinfo[1]),
    .d(i_exu_op1[17]),
    .e(i_exu_op2[17]),
    .o(_al_u1238_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1239 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[17]),
    .d(i_exu_op2[17]),
    .o(_al_u1239_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u1240 (
    .a(_al_u1238_o),
    .b(_al_u1239_o),
    .c(\u_EXU_ALU/n0 [17]),
    .d(i_decinfo_grp[5]),
    .o(_al_u1240_o));
  AL_MAP_LUT5 #(
    .EQN("~((E*D*A)*~(B)*~(C)+(E*D*A)*B*~(C)+~((E*D*A))*B*C+(E*D*A)*B*C)"),
    .INIT(32'h353f3f3f))
    _al_u1241 (
    .a(\u_EXU_ALU/n255_lutinv ),
    .b(i_exu_op1[31]),
    .c(i_exu_op2[4]),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[0]),
    .o(_al_u1241_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*C*B))"),
    .INIT(16'haa2a))
    _al_u1242 (
    .a(_al_u1240_o),
    .b(_al_u1065_o),
    .c(_al_u961_o),
    .d(_al_u1241_o),
    .o(_al_u1242_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1243 (
    .a(\u_EXU_ALU/n351_lutinv ),
    .b(_al_u965_o),
    .c(_al_u1227_o),
    .o(_al_u1243_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D*C*B*A))"),
    .INIT(32'h7fff0000))
    _al_u1244 (
    .a(_al_u911_o),
    .b(_al_u915_o),
    .c(_al_u1243_o),
    .d(_al_u917_o),
    .e(i_decinfo_grp[0]),
    .o(_al_u1244_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1245 (
    .a(bju_rdwdata[17]),
    .b(bju_rdwen),
    .c(i_csr_rdata[17]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1245_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*B*~(D*~A)))"),
    .INIT(32'h00007f3f))
    _al_u1246 (
    .a(_al_u1237_o),
    .b(_al_u1242_o),
    .c(_al_u1244_o),
    .d(\u_EXU_ALU/u1029_sel_is_0_o ),
    .e(_al_u1245_o),
    .o(o_rdwdata0[17]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1247 (
    .a(i_exu_op1[17]),
    .b(i_exu_op1[16]),
    .c(i_exu_op2[0]),
    .o(_al_u1247_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1248 (
    .a(_al_u1216_o),
    .b(_al_u1247_o),
    .c(i_exu_op2[1]),
    .o(\u_EXU_ALU/n125_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("~(~(~B*~(C)*~(E)+~B*C*~(E)+~(~B)*C*E+~B*C*E)*~(A)*~(D)+~(~B*~(C)*~(E)+~B*C*~(E)+~(~B)*C*E+~B*C*E)*A*~(D)+~(~(~B*~(C)*~(E)+~B*C*~(E)+~(~B)*C*E+~B*C*E))*A*D+~(~B*~(C)*~(E)+~B*C*~(E)+~(~B)*C*E+~B*C*E)*A*D)"),
    .INIT(32'h55f05533))
    _al_u1249 (
    .a(\u_EXU_ALU/n84_lutinv ),
    .b(\u_EXU_ALU/n125_lutinv ),
    .c(_al_u1185_o),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(_al_u1249_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1250 (
    .a(_al_u1114_o),
    .b(_al_u1115_o),
    .c(_al_u1057_o),
    .d(i_exu_op2[2]),
    .o(_al_u1250_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~C)*~(~D*~A))"),
    .INIT(32'h30203322))
    _al_u1251 (
    .a(_al_u1249_o),
    .b(_al_u1250_o),
    .c(_al_u1121_o),
    .d(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .e(_al_u1059_o),
    .o(_al_u1251_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1252 (
    .a(\u_EXU_ALU/n352_lutinv ),
    .b(_al_u965_o),
    .c(_al_u1227_o),
    .o(_al_u1252_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D*C*B*A))"),
    .INIT(32'h7fff0000))
    _al_u1253 (
    .a(_al_u911_o),
    .b(_al_u915_o),
    .c(_al_u1252_o),
    .d(_al_u917_o),
    .e(i_decinfo_grp[0]),
    .o(_al_u1253_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1254 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[16]),
    .c(i_exu_op2[16]),
    .o(\u_EXU_ALU/alu_and [16]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*B))"),
    .INIT(16'h0105))
    _al_u1255 (
    .a(alu2lsu_result[16]),
    .b(\u_EXU_ALU/n33 [16]),
    .c(\u_EXU_ALU/alu_and [16]),
    .d(i_decinfo[1]),
    .o(_al_u1255_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1256 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[16]),
    .d(i_exu_op2[16]),
    .o(_al_u1256_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*C*B*~(E*A))"),
    .INIT(32'h004000c0))
    _al_u1257 (
    .a(_al_u1066_o),
    .b(_al_u1253_o),
    .c(_al_u1255_o),
    .d(_al_u1256_o),
    .e(_al_u1193_o),
    .o(_al_u1257_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1258 (
    .a(bju_rdwdata[16]),
    .b(bju_rdwen),
    .c(i_csr_rdata[16]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1258_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(C*~A)))"),
    .INIT(16'h0073))
    _al_u1259 (
    .a(_al_u1251_o),
    .b(_al_u1257_o),
    .c(\u_EXU_ALU/u1029_sel_is_0_o ),
    .d(_al_u1258_o),
    .o(o_rdwdata0[16]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1260 (
    .a(i_exu_op1[14]),
    .b(i_exu_op1[13]),
    .c(i_exu_op2[0]),
    .d(i_exu_op2[1]),
    .o(_al_u1260_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h530f))
    _al_u1261 (
    .a(i_exu_op1[16]),
    .b(i_exu_op1[15]),
    .c(_al_u1260_o),
    .d(i_exu_op2[1]),
    .o(_al_u1261_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1262 (
    .a(i_exu_op1[12]),
    .b(i_exu_op1[11]),
    .c(i_exu_op2[0]),
    .o(_al_u1262_o));
  AL_MAP_LUT5 #(
    .EQN("(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haa33aa0f))
    _al_u1263 (
    .a(_al_u1262_o),
    .b(i_exu_op1[10]),
    .c(i_exu_op1[9]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1263_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1264 (
    .a(_al_u1261_o),
    .b(_al_u1263_o),
    .c(i_exu_op2[2]),
    .o(\u_EXU_ALU/n100_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1265 (
    .a(i_exu_op1[2]),
    .b(i_exu_op1[1]),
    .c(i_exu_op2[0]),
    .o(_al_u1265_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1266 (
    .a(i_exu_op1[4]),
    .b(i_exu_op1[3]),
    .c(i_exu_op2[0]),
    .o(_al_u1266_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1267 (
    .a(i_exu_op1[8]),
    .b(i_exu_op1[7]),
    .c(i_exu_op2[0]),
    .o(_al_u1267_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1268 (
    .a(i_exu_op1[6]),
    .b(i_exu_op1[5]),
    .c(i_exu_op2[0]),
    .o(_al_u1268_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u1269 (
    .a(_al_u1267_o),
    .b(_al_u1268_o),
    .c(i_exu_op2[1]),
    .d(i_exu_op2[2]),
    .o(_al_u1269_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u1270 (
    .a(_al_u1265_o),
    .b(_al_u1266_o),
    .c(_al_u1269_o),
    .d(i_exu_op2[2]),
    .o(_al_u1270_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E)*~(A)*~(D)+~(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E)*A*~(D)+~(~(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E))*A*D+~(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E)*A*D)"),
    .INIT(32'haa33aaf0))
    _al_u1271 (
    .a(_al_u1234_o),
    .b(\u_EXU_ALU/n100_lutinv ),
    .c(_al_u1270_o),
    .d(i_exu_op2[4]),
    .e(i_exu_op2[3]),
    .o(_al_u1271_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D*B)*~(C*A))"),
    .INIT(32'h135f5f5f))
    _al_u1272 (
    .a(\u_EXU_ALU/n33 [1]),
    .b(i_decinfo[6]),
    .c(i_decinfo[1]),
    .d(i_exu_op1[1]),
    .e(i_exu_op2[1]),
    .o(_al_u1272_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1273 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[1]),
    .d(i_exu_op2[1]),
    .o(_al_u1273_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u1274 (
    .a(alu2lsu_result[1]),
    .b(_al_u1272_o),
    .c(_al_u1273_o),
    .d(i_decinfo_grp[0]),
    .o(_al_u1274_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(E*D*C*A))"),
    .INIT(32'h4ccccccc))
    _al_u1275 (
    .a(\u_EXU_ALU/n281_neg_lutinv ),
    .b(_al_u1274_o),
    .c(\u_EXU_ALU/n351_lutinv ),
    .d(_al_u965_o),
    .e(_al_u1026_o),
    .o(_al_u1275_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1276 (
    .a(_al_u937_o),
    .b(_al_u938_o),
    .c(_al_u1005_o),
    .o(_al_u1276_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1277 (
    .a(i_exu_op1[31]),
    .b(i_exu_op2[2]),
    .o(_al_u1277_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u1278 (
    .a(_al_u1007_o),
    .b(_al_u1277_o),
    .c(i_exu_op2[4]),
    .d(i_exu_op2[3]),
    .o(_al_u1278_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1279 (
    .a(_al_u1276_o),
    .b(_al_u1002_o),
    .c(_al_u1278_o),
    .d(_al_u1004_o),
    .e(i_decinfo[4]),
    .o(_al_u1279_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    _al_u1280 (
    .a(_al_u911_o),
    .b(_al_u917_o),
    .c(_al_u951_o),
    .d(_al_u912_o),
    .e(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .o(_al_u1280_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~((C*B)*~(E)*~(A)+(C*B)*E*~(A)+~((C*B))*E*A+(C*B)*E*A))"),
    .INIT(32'h001500bf))
    _al_u1281 (
    .a(bju_rdwen),
    .b(i_csr_rdata[1]),
    .c(i_decinfo_grp[4]),
    .d(i_decinfo_grp[0]),
    .e(i_iaddr[1]),
    .o(_al_u1281_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~C*B*~(D*~A)))"),
    .INIT(32'h0000f7f3))
    _al_u1282 (
    .a(_al_u1271_o),
    .b(_al_u1275_o),
    .c(_al_u1279_o),
    .d(_al_u1280_o),
    .e(_al_u1281_o),
    .o(o_rdwdata0[1]));
  AL_MAP_LUT5 #(
    .EQN("~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'h55cc55f0))
    _al_u1283 (
    .a(_al_u1247_o),
    .b(i_exu_op1[15]),
    .c(i_exu_op1[14]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(\u_EXU_ALU/n127_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1284 (
    .a(i_exu_op1[11]),
    .b(i_exu_op1[10]),
    .c(i_exu_op2[0]),
    .o(_al_u1284_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(~A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33aa0faa))
    _al_u1285 (
    .a(_al_u1284_o),
    .b(i_exu_op1[13]),
    .c(i_exu_op1[12]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1285_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(16'ha030))
    _al_u1286 (
    .a(\u_EXU_ALU/n127_lutinv ),
    .b(_al_u1285_o),
    .c(_al_u930_o),
    .d(i_exu_op2[2]),
    .o(_al_u1286_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1287 (
    .a(i_exu_op1[7]),
    .b(i_exu_op1[6]),
    .c(i_exu_op2[0]),
    .o(_al_u1287_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(~A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33aa0faa))
    _al_u1288 (
    .a(_al_u1287_o),
    .b(i_exu_op1[9]),
    .c(i_exu_op1[8]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1288_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~D*~(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'h0f0a0f0c))
    _al_u1289 (
    .a(i_exu_op1[3]),
    .b(i_exu_op1[2]),
    .c(i_exu_op2[2]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1289_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1290 (
    .a(i_exu_op1[5]),
    .b(i_exu_op1[4]),
    .c(i_exu_op2[1]),
    .d(i_exu_op2[0]),
    .o(_al_u1290_o));
  AL_MAP_LUT5 #(
    .EQN("(D*~(~(~C*B)*~(E*~A)))"),
    .INIT(32'h5d000c00))
    _al_u1291 (
    .a(_al_u1288_o),
    .b(_al_u1289_o),
    .c(_al_u1290_o),
    .d(_al_u924_o),
    .e(i_exu_op2[2]),
    .o(_al_u1291_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~D*~C*~(E*~A)))"),
    .INIT(32'hccc4ccc0))
    _al_u1292 (
    .a(_al_u1218_o),
    .b(_al_u1280_o),
    .c(_al_u1286_o),
    .d(_al_u1291_o),
    .e(i_exu_op2[4]),
    .o(_al_u1292_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h155f))
    _al_u1293 (
    .a(i_decinfo[7]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[2]),
    .d(i_exu_op2[2]),
    .o(_al_u1293_o));
  AL_MAP_LUT5 #(
    .EQN("(E*B*~A*~(D*C))"),
    .INIT(32'h04440000))
    _al_u1294 (
    .a(alu2lsu_result[2]),
    .b(_al_u1293_o),
    .c(\u_EXU_ALU/n33 [2]),
    .d(i_decinfo[1]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1294_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~C*A))"),
    .INIT(16'hc4cc))
    _al_u1295 (
    .a(_al_u1027_o),
    .b(_al_u1294_o),
    .c(_al_u970_o),
    .d(_al_u965_o),
    .o(_al_u1295_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1296 (
    .a(i_exu_op2[2]),
    .b(i_exu_op2[1]),
    .o(_al_u1296_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1297 (
    .a(_al_u1006_o),
    .b(_al_u1193_o),
    .c(_al_u1296_o),
    .d(i_decinfo[4]),
    .e(i_exu_op2[3]),
    .o(_al_u1297_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(B)*~(A)+(D*C)*B*~(A)+~((D*C))*B*A+(D*C)*B*A))"),
    .INIT(32'h00002777))
    _al_u1298 (
    .a(bju_rdwen),
    .b(bju_rdwdata[2]),
    .c(i_csr_rdata[2]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1298_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u1299 (
    .a(i_decinfo[5]),
    .b(i_exu_op1[2]),
    .c(i_exu_op2[2]),
    .o(\u_EXU_ALU/alu_xor [2]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~E*~C*B*~A))"),
    .INIT(32'h00ff00fb))
    _al_u1300 (
    .a(_al_u1292_o),
    .b(_al_u1295_o),
    .c(_al_u1297_o),
    .d(_al_u1298_o),
    .e(\u_EXU_ALU/alu_xor [2]),
    .o(o_rdwdata0[2]));
  AL_MAP_LUT5 #(
    .EQN("(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haa33aa0f))
    _al_u1301 (
    .a(_al_u1232_o),
    .b(i_exu_op1[16]),
    .c(i_exu_op1[15]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1301_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(~A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33aa0faa))
    _al_u1302 (
    .a(_al_u1262_o),
    .b(i_exu_op1[14]),
    .c(i_exu_op1[13]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1302_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1303 (
    .a(_al_u1301_o),
    .b(_al_u1302_o),
    .c(i_exu_op2[2]),
    .o(\u_EXU_ALU/n97_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(~A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33aa0faa))
    _al_u1304 (
    .a(_al_u1267_o),
    .b(i_exu_op1[10]),
    .c(i_exu_op1[9]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1304_o));
  AL_MAP_LUT5 #(
    .EQN("((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'haaf0aacc))
    _al_u1305 (
    .a(_al_u1304_o),
    .b(_al_u1266_o),
    .c(_al_u1268_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1305_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E)*~(A)*~(D)+~(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E)*A*~(D)+~(~(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E))*A*D+~(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E)*A*D)"),
    .INIT(32'haa33aaf0))
    _al_u1306 (
    .a(_al_u1201_o),
    .b(\u_EXU_ALU/n97_lutinv ),
    .c(_al_u1305_o),
    .d(i_exu_op2[4]),
    .e(i_exu_op2[3]),
    .o(_al_u1306_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1307 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[3]),
    .c(i_exu_op2[3]),
    .o(\u_EXU_ALU/alu_and [3]));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u1308 (
    .a(\u_EXU_ALU/alu_and [3]),
    .b(\u_EXU_ALU/n33 [3]),
    .c(i_decinfo[1]),
    .d(i_decinfo_grp[0]),
    .o(_al_u1308_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1309 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[3]),
    .d(i_exu_op2[3]),
    .o(_al_u1309_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u1310 (
    .a(_al_u1308_o),
    .b(alu2lsu_result[3]),
    .c(_al_u1309_o),
    .o(_al_u1310_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*A))"),
    .INIT(16'h4ccc))
    _al_u1311 (
    .a(\u_EXU_ALU/n281_neg_lutinv ),
    .b(_al_u1310_o),
    .c(\u_EXU_ALU/n413_lutinv ),
    .d(_al_u1026_o),
    .o(_al_u1311_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1312 (
    .a(\u_EXU_ALU/n256_lutinv ),
    .b(i_exu_op2[4]),
    .c(i_exu_op2[3]),
    .o(_al_u1312_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1313 (
    .a(_al_u1276_o),
    .b(_al_u1002_o),
    .c(_al_u1312_o),
    .d(_al_u1004_o),
    .e(i_decinfo[4]),
    .o(_al_u1313_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(B)*~(A)+(D*C)*B*~(A)+~((D*C))*B*A+(D*C)*B*A))"),
    .INIT(32'h00002777))
    _al_u1314 (
    .a(bju_rdwen),
    .b(bju_rdwdata[3]),
    .c(i_csr_rdata[3]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1314_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~C*B*~(D*~A)))"),
    .INIT(32'h0000f7f3))
    _al_u1315 (
    .a(_al_u1306_o),
    .b(_al_u1311_o),
    .c(_al_u1313_o),
    .d(_al_u1280_o),
    .e(_al_u1314_o),
    .o(o_rdwdata0[3]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(C*B)*~(D*A))"),
    .INIT(32'h153f0000))
    _al_u1316 (
    .a(\u_EXU_ALU/n0 [4]),
    .b(\u_EXU_ALU/n33 [4]),
    .c(i_decinfo[1]),
    .d(i_decinfo_grp[5]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1316_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h155f))
    _al_u1317 (
    .a(i_decinfo[7]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[4]),
    .d(i_exu_op2[4]),
    .o(_al_u1317_o));
  AL_MAP_LUT5 #(
    .EQN("(B*A*~(C*(E@D)))"),
    .INIT(32'h88080888))
    _al_u1318 (
    .a(_al_u1316_o),
    .b(_al_u1317_o),
    .c(i_decinfo[5]),
    .d(i_exu_op1[4]),
    .e(i_exu_op2[4]),
    .o(_al_u1318_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1319 (
    .a(i_decinfo[4]),
    .b(i_exu_op2[4]),
    .o(_al_u1319_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*A))"),
    .INIT(16'h4ccc))
    _al_u1320 (
    .a(\u_EXU_ALU/n179_neg_lutinv ),
    .b(_al_u1318_o),
    .c(\u_EXU_ALU/n241_lutinv ),
    .d(_al_u1319_o),
    .o(_al_u1320_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1321 (
    .a(i_exu_op1[13]),
    .b(i_exu_op1[12]),
    .c(i_exu_op2[0]),
    .d(i_exu_op2[1]),
    .o(_al_u1321_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h530f))
    _al_u1322 (
    .a(i_exu_op1[15]),
    .b(i_exu_op1[14]),
    .c(_al_u1321_o),
    .d(i_exu_op2[1]),
    .o(_al_u1322_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u1323 (
    .a(i_decinfo[4]),
    .b(i_decinfo[3]),
    .c(i_exu_op2[4]),
    .o(_al_u1323_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(C*(~B*~(A)*~(E)+~B*A*~(E)+~(~B)*A*E+~B*A*E)))"),
    .INIT(32'h005f00cf))
    _al_u1324 (
    .a(\u_EXU_ALU/n125_lutinv ),
    .b(_al_u1322_o),
    .c(_al_u1134_o),
    .d(_al_u1323_o),
    .e(i_exu_op2[2]),
    .o(_al_u1324_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1325 (
    .a(i_exu_op1[5]),
    .b(i_exu_op1[4]),
    .c(i_exu_op2[0]),
    .o(_al_u1325_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~D*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)))"),
    .INIT(32'haa22aa0a))
    _al_u1326 (
    .a(_al_u954_o),
    .b(_al_u1287_o),
    .c(_al_u1325_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1326_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1327 (
    .a(i_exu_op1[9]),
    .b(i_exu_op1[8]),
    .c(i_exu_op2[0]),
    .o(_al_u1327_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u1328 (
    .a(_al_u1284_o),
    .b(_al_u1327_o),
    .c(i_exu_op2[2]),
    .d(i_exu_op2[1]),
    .o(_al_u1328_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(~D*C))"),
    .INIT(16'h2202))
    _al_u1329 (
    .a(_al_u1324_o),
    .b(_al_u1195_o),
    .c(_al_u1326_o),
    .d(_al_u1328_o),
    .o(_al_u1329_o));
  AL_MAP_LUT5 #(
    .EQN("(D*~(A*~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)))"),
    .INIT(32'hdd00f500))
    _al_u1330 (
    .a(_al_u1159_o),
    .b(_al_u1048_o),
    .c(_al_u1049_o),
    .d(i_exu_op2[4]),
    .e(i_exu_op2[1]),
    .o(_al_u1330_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)))"),
    .INIT(32'h88aaa0aa))
    _al_u1331 (
    .a(_al_u1330_o),
    .b(_al_u1124_o),
    .c(_al_u1185_o),
    .d(_al_u954_o),
    .e(i_exu_op2[2]),
    .o(_al_u1331_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(B)*~(A)+(D*C)*B*~(A)+~((D*C))*B*A+(D*C)*B*A))"),
    .INIT(32'h00002777))
    _al_u1332 (
    .a(bju_rdwen),
    .b(bju_rdwdata[4]),
    .c(i_csr_rdata[4]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1332_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(A*~(D*~C*~B)))"),
    .INIT(32'h00005755))
    _al_u1333 (
    .a(_al_u1320_o),
    .b(_al_u1329_o),
    .c(_al_u1331_o),
    .d(\u_EXU_ALU/n281_neg_lutinv ),
    .e(_al_u1332_o),
    .o(o_rdwdata0[4]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1334 (
    .a(_al_u1181_o),
    .b(\u_EXU_ALU/n281_neg_lutinv ),
    .c(i_exu_op2[4]),
    .o(_al_u1334_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1335 (
    .a(_al_u1233_o),
    .b(_al_u1261_o),
    .c(_al_u1134_o),
    .d(i_exu_op2[2]),
    .o(_al_u1335_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*(~A*~(B)*~(E)+~A*B*~(E)+~(~A)*B*E+~A*B*E)))"),
    .INIT(32'h030f0a0f))
    _al_u1336 (
    .a(_al_u1102_o),
    .b(\u_EXU_ALU/n351_lutinv ),
    .c(_al_u1323_o),
    .d(_al_u1059_o),
    .e(i_exu_op2[2]),
    .o(_al_u1336_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~D*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)))"),
    .INIT(32'haa22aa0a))
    _al_u1337 (
    .a(_al_u954_o),
    .b(_al_u1267_o),
    .c(_al_u1268_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1337_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~A*~(C*~(E*D)))"),
    .INIT(32'h44040404))
    _al_u1338 (
    .a(_al_u1335_o),
    .b(_al_u1336_o),
    .c(_al_u1337_o),
    .d(_al_u1263_o),
    .e(i_exu_op2[2]),
    .o(_al_u1338_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u1339 (
    .a(\u_EXU_ALU/n33 [5]),
    .b(i_decinfo[1]),
    .c(i_decinfo_grp[0]),
    .o(_al_u1339_o));
  AL_MAP_LUT5 #(
    .EQN("(A*(~(B)*~(C)*~(D)*~(E)+B*~(C)*~(D)*~(E)+~(B)*C*~(D)*~(E)+B*C*~(D)*~(E)+~(B)*~(C)*D*~(E)+B*~(C)*D*~(E)+~(B)*~(C)*~(D)*E+B*~(C)*~(D)*E+~(B)*~(C)*D*E+~(B)*C*D*E))"),
    .INIT(32'h220a0aaa))
    _al_u1340 (
    .a(_al_u1339_o),
    .b(i_decinfo[6]),
    .c(i_decinfo[5]),
    .d(i_exu_op1[5]),
    .e(i_exu_op2[5]),
    .o(_al_u1340_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(~D*~B))"),
    .INIT(16'ha080))
    _al_u1341 (
    .a(_al_u1108_o),
    .b(_al_u1007_o),
    .c(i_exu_op2[4]),
    .d(i_exu_op2[2]),
    .o(_al_u1341_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~(~E*~D)*B)*~(C*A))"),
    .INIT(32'h1313135f))
    _al_u1342 (
    .a(\u_EXU_ALU/n0 [5]),
    .b(i_decinfo[7]),
    .c(i_decinfo_grp[5]),
    .d(i_exu_op1[5]),
    .e(i_exu_op2[5]),
    .o(_al_u1342_o));
  AL_MAP_LUT5 #(
    .EQN("(E*B*~(D*C*A))"),
    .INIT(32'h4ccc0000))
    _al_u1343 (
    .a(_al_u1065_o),
    .b(_al_u1340_o),
    .c(_al_u961_o),
    .d(_al_u1341_o),
    .e(_al_u1342_o),
    .o(_al_u1343_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(B)*~(A)+(D*C)*B*~(A)+~((D*C))*B*A+(D*C)*B*A))"),
    .INIT(32'h00002777))
    _al_u1344 (
    .a(bju_rdwen),
    .b(bju_rdwdata[5]),
    .c(i_csr_rdata[5]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1344_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(~B*A)))"),
    .INIT(16'h002f))
    _al_u1345 (
    .a(_al_u1334_o),
    .b(_al_u1338_o),
    .c(_al_u1343_o),
    .d(_al_u1344_o),
    .o(o_rdwdata0[5]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1346 (
    .a(_al_u1163_o),
    .b(\u_EXU_ALU/n281_neg_lutinv ),
    .c(i_exu_op2[4]),
    .o(_al_u1346_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(16'h50c0))
    _al_u1347 (
    .a(_al_u1217_o),
    .b(\u_EXU_ALU/n127_lutinv ),
    .c(_al_u1134_o),
    .d(i_exu_op2[2]),
    .o(_al_u1347_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'h0c0f0a0f))
    _al_u1348 (
    .a(_al_u1088_o),
    .b(_al_u970_o),
    .c(_al_u1323_o),
    .d(_al_u1059_o),
    .e(i_exu_op2[2]),
    .o(_al_u1348_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~D*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)))"),
    .INIT(32'haa22aa0a))
    _al_u1349 (
    .a(_al_u954_o),
    .b(_al_u1327_o),
    .c(_al_u1287_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1349_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~A*~(C*~(E*D)))"),
    .INIT(32'h44040404))
    _al_u1350 (
    .a(_al_u1347_o),
    .b(_al_u1348_o),
    .c(_al_u1349_o),
    .d(_al_u1285_o),
    .e(i_exu_op2[2]),
    .o(_al_u1350_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1351 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[6]),
    .d(i_exu_op2[6]),
    .o(_al_u1351_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1352 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[6]),
    .c(i_exu_op2[6]),
    .o(\u_EXU_ALU/alu_and [6]));
  AL_MAP_LUT5 #(
    .EQN("(~C*~B*~A*~(E*D))"),
    .INIT(32'h00010101))
    _al_u1353 (
    .a(alu2lsu_result[6]),
    .b(_al_u1351_o),
    .c(\u_EXU_ALU/alu_and [6]),
    .d(\u_EXU_ALU/n33 [6]),
    .e(i_decinfo[1]),
    .o(_al_u1353_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u1354 (
    .a(_al_u1108_o),
    .b(_al_u948_o),
    .c(i_exu_op2[4]),
    .o(_al_u1354_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*A))"),
    .INIT(16'h4ccc))
    _al_u1355 (
    .a(_al_u1065_o),
    .b(_al_u1353_o),
    .c(_al_u961_o),
    .d(_al_u1354_o),
    .o(_al_u1355_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(B)*~(A)+(D*C)*B*~(A)+~((D*C))*B*A+(D*C)*B*A)"),
    .INIT(16'h2777))
    _al_u1356 (
    .a(bju_rdwen),
    .b(bju_rdwdata[6]),
    .c(i_csr_rdata[6]),
    .d(i_decinfo_grp[4]),
    .o(_al_u1356_o));
  AL_MAP_LUT5 #(
    .EQN("~(D*~((C*~(~B*A)))*~(E)+D*(C*~(~B*A))*~(E)+~(D)*(C*~(~B*A))*E+D*(C*~(~B*A))*E)"),
    .INIT(32'h2f2f00ff))
    _al_u1357 (
    .a(_al_u1346_o),
    .b(_al_u1350_o),
    .c(_al_u1355_o),
    .d(_al_u1356_o),
    .e(i_decinfo_grp[0]),
    .o(o_rdwdata0[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u1358 (
    .a(_al_u1136_o),
    .b(\u_EXU_ALU/n281_neg_lutinv ),
    .c(i_exu_op2[4]),
    .o(_al_u1358_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)))"),
    .INIT(32'h44555055))
    _al_u1359 (
    .a(_al_u1139_o),
    .b(_al_u1200_o),
    .c(_al_u1301_o),
    .d(_al_u1134_o),
    .e(i_exu_op2[2]),
    .o(_al_u1359_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D*B)*~(C*A))"),
    .INIT(32'h135f5f5f))
    _al_u1360 (
    .a(\u_EXU_ALU/n33 [7]),
    .b(i_decinfo[6]),
    .c(i_decinfo[1]),
    .d(i_exu_op1[7]),
    .e(i_exu_op2[7]),
    .o(_al_u1360_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1361 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[7]),
    .d(i_exu_op2[7]),
    .o(_al_u1361_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~B*A*~(D*C))"),
    .INIT(32'h02220000))
    _al_u1362 (
    .a(_al_u1360_o),
    .b(_al_u1361_o),
    .c(\u_EXU_ALU/n0 [7]),
    .d(i_decinfo_grp[5]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1362_o));
  AL_MAP_LUT5 #(
    .EQN("(D*C*B*~(~E*A))"),
    .INIT(32'hc0004000))
    _al_u1363 (
    .a(_al_u948_o),
    .b(i_exu_op1[31]),
    .c(i_exu_op2[4]),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[0]),
    .o(_al_u1363_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*A))"),
    .INIT(16'h4ccc))
    _al_u1364 (
    .a(_al_u1065_o),
    .b(_al_u1362_o),
    .c(_al_u961_o),
    .d(_al_u1363_o),
    .o(_al_u1364_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(C*~(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)))"),
    .INIT(32'h00cf00af))
    _al_u1365 (
    .a(_al_u1304_o),
    .b(_al_u1302_o),
    .c(_al_u954_o),
    .d(_al_u1323_o),
    .e(i_exu_op2[2]),
    .o(_al_u1365_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(B)*~(A)+(D*C)*B*~(A)+~((D*C))*B*A+(D*C)*B*A))"),
    .INIT(32'h00002777))
    _al_u1366 (
    .a(bju_rdwen),
    .b(bju_rdwdata[7]),
    .c(i_csr_rdata[7]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1366_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*~(A*~(D*B))))"),
    .INIT(32'h00002faf))
    _al_u1367 (
    .a(_al_u1358_o),
    .b(_al_u1359_o),
    .c(_al_u1364_o),
    .d(_al_u1365_o),
    .e(_al_u1366_o),
    .o(o_rdwdata0[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1368 (
    .a(_al_u1048_o),
    .b(_al_u1049_o),
    .c(i_exu_op2[1]),
    .o(_al_u1368_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~(~B*~A))"),
    .INIT(16'h00e0))
    _al_u1369 (
    .a(i_decinfo[4]),
    .b(i_decinfo[3]),
    .c(i_exu_op2[4]),
    .d(i_exu_op2[3]),
    .o(_al_u1369_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1370 (
    .a(_al_u1368_o),
    .b(_al_u1124_o),
    .c(_al_u1369_o),
    .d(i_exu_op2[2]),
    .o(_al_u1370_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u1371 (
    .a(_al_u1117_o),
    .b(_al_u1370_o),
    .c(_al_u1026_o),
    .o(_al_u1371_o));
  AL_MAP_LUT3 #(
    .EQN("~(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'h3a))
    _al_u1372 (
    .a(\u_EXU_ALU/n125_lutinv ),
    .b(_al_u1185_o),
    .c(i_exu_op2[2]),
    .o(\u_EXU_ALU/n92_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'h5533550f))
    _al_u1373 (
    .a(_al_u1322_o),
    .b(_al_u1284_o),
    .c(_al_u1327_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(\u_EXU_ALU/n101_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u1374 (
    .a(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .b(i_exu_op2[4]),
    .o(_al_u1374_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u1375 (
    .a(\u_EXU_ALU/n92_lutinv ),
    .b(\u_EXU_ALU/n101_lutinv ),
    .c(_al_u1374_o),
    .d(i_exu_op2[3]),
    .o(_al_u1375_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D*B)*~(C*A))"),
    .INIT(32'h135f5f5f))
    _al_u1376 (
    .a(\u_EXU_ALU/n33 [8]),
    .b(i_decinfo[6]),
    .c(i_decinfo[1]),
    .d(i_exu_op1[8]),
    .e(i_exu_op2[8]),
    .o(_al_u1376_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1377 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[8]),
    .d(i_exu_op2[8]),
    .o(_al_u1377_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~B*A*~(D*C))"),
    .INIT(32'h02220000))
    _al_u1378 (
    .a(_al_u1376_o),
    .b(_al_u1377_o),
    .c(\u_EXU_ALU/n0 [8]),
    .d(i_decinfo_grp[5]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1378_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(E*D*C*A))"),
    .INIT(32'h4ccccccc))
    _al_u1379 (
    .a(_al_u1065_o),
    .b(_al_u1378_o),
    .c(_al_u961_o),
    .d(_al_u1193_o),
    .e(i_exu_op2[3]),
    .o(_al_u1379_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(B)*~(A)+(D*C)*B*~(A)+~((D*C))*B*A+(D*C)*B*A))"),
    .INIT(32'h00002777))
    _al_u1380 (
    .a(bju_rdwen),
    .b(bju_rdwdata[8]),
    .c(i_csr_rdata[8]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1380_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*~(D*~(~B*A))))"),
    .INIT(32'h0000df0f))
    _al_u1381 (
    .a(_al_u1371_o),
    .b(_al_u1375_o),
    .c(_al_u1379_o),
    .d(\u_EXU_ALU/n281_neg_lutinv ),
    .e(_al_u1380_o),
    .o(o_rdwdata0[8]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1382 (
    .a(_al_u1261_o),
    .b(_al_u1263_o),
    .c(_al_u954_o),
    .d(i_exu_op2[2]),
    .o(_al_u1382_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1383 (
    .a(_al_u1179_o),
    .b(_al_u1233_o),
    .c(_al_u1134_o),
    .d(i_exu_op2[2]),
    .o(_al_u1383_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u1384 (
    .a(_al_u1103_o),
    .b(_al_u1382_o),
    .c(_al_u1383_o),
    .d(i_exu_op2[4]),
    .o(_al_u1384_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*(~(B)*~(C)*~(D)*~(E)+B*~(C)*~(D)*~(E)+~(B)*C*~(D)*~(E)+B*C*~(D)*~(E)+~(B)*~(C)*D*~(E)+~(B)*~(C)*~(D)*E+~(B)*~(C)*D*E+~(B)*C*D*E))"),
    .INIT(32'h11010155))
    _al_u1385 (
    .a(alu2lsu_result[9]),
    .b(i_decinfo[7]),
    .c(i_decinfo[5]),
    .d(i_exu_op1[9]),
    .e(i_exu_op2[9]),
    .o(_al_u1385_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1386 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[9]),
    .c(i_exu_op2[9]),
    .o(\u_EXU_ALU/alu_and [9]));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u1387 (
    .a(\u_EXU_ALU/alu_and [9]),
    .b(\u_EXU_ALU/n33 [9]),
    .c(i_decinfo[1]),
    .d(i_decinfo_grp[0]),
    .o(_al_u1387_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*~(E*~D*A))"),
    .INIT(32'hc040c0c0))
    _al_u1388 (
    .a(_al_u1006_o),
    .b(_al_u1385_o),
    .c(_al_u1387_o),
    .d(_al_u1109_o),
    .e(_al_u1319_o),
    .o(_al_u1388_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(C*B)))"),
    .INIT(16'h80aa))
    _al_u1389 (
    .a(\u_EXU_ALU/n281_neg_lutinv ),
    .b(\u_EXU_ALU/n83_lutinv ),
    .c(_al_u954_o),
    .d(i_exu_op2[4]),
    .o(_al_u1389_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(B)*~(A)+(D*C)*B*~(A)+~((D*C))*B*A+(D*C)*B*A))"),
    .INIT(32'h00002777))
    _al_u1390 (
    .a(bju_rdwen),
    .b(bju_rdwdata[9]),
    .c(i_csr_rdata[9]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1390_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(C*~A)))"),
    .INIT(16'h0073))
    _al_u1391 (
    .a(_al_u1384_o),
    .b(_al_u1388_o),
    .c(_al_u1389_o),
    .d(_al_u1390_o),
    .o(o_rdwdata0[9]));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u1392 (
    .a(_al_u911_o),
    .b(_al_u917_o),
    .c(_al_u951_o),
    .d(_al_u912_o),
    .e(_al_u1323_o),
    .o(_al_u1392_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u1393 (
    .a(\u_EXU_ALU/n33 [10]),
    .b(i_decinfo[1]),
    .c(i_decinfo_grp[0]),
    .o(_al_u1393_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h155f))
    _al_u1394 (
    .a(i_decinfo[7]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[10]),
    .d(i_exu_op2[10]),
    .o(_al_u1394_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u1395 (
    .a(i_decinfo[5]),
    .b(i_exu_op1[10]),
    .c(i_exu_op2[10]),
    .o(\u_EXU_ALU/alu_xor [10]));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*A*~(E*D))"),
    .INIT(32'h00080808))
    _al_u1396 (
    .a(_al_u1393_o),
    .b(_al_u1394_o),
    .c(\u_EXU_ALU/alu_xor [10]),
    .d(\u_EXU_ALU/n0 [10]),
    .e(i_decinfo_grp[5]),
    .o(_al_u1396_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(D*B)))"),
    .INIT(16'he0a0))
    _al_u1397 (
    .a(_al_u1108_o),
    .b(_al_u1277_o),
    .c(_al_u1319_o),
    .d(i_exu_op2[1]),
    .o(_al_u1397_o));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C*B)*~(E*A))"),
    .INIT(32'h15003f00))
    _al_u1398 (
    .a(\u_EXU_ALU/n179_neg_lutinv ),
    .b(_al_u1392_o),
    .c(\u_EXU_ALU/n49_lutinv ),
    .d(_al_u1396_o),
    .e(_al_u1397_o),
    .o(_al_u1398_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1399 (
    .a(_al_u1089_o),
    .b(i_decinfo[2]),
    .o(_al_u1399_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1400 (
    .a(_al_u1162_o),
    .b(_al_u1217_o),
    .c(_al_u1134_o),
    .d(i_exu_op2[2]),
    .o(_al_u1400_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E)))"),
    .INIT(32'h11555055))
    _al_u1401 (
    .a(_al_u1400_o),
    .b(\u_EXU_ALU/n127_lutinv ),
    .c(_al_u1285_o),
    .d(_al_u954_o),
    .e(i_exu_op2[2]),
    .o(_al_u1401_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(B)*~(A)+(D*C)*B*~(A)+~((D*C))*B*A+(D*C)*B*A))"),
    .INIT(32'h00002777))
    _al_u1402 (
    .a(bju_rdwen),
    .b(bju_rdwdata[10]),
    .c(i_csr_rdata[10]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1402_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(A*~(D*~(C*~B))))"),
    .INIT(32'h0000df55))
    _al_u1403 (
    .a(_al_u1398_o),
    .b(_al_u1399_o),
    .c(_al_u1401_o),
    .d(\u_EXU_ALU/u1029_sel_is_0_o ),
    .e(_al_u1402_o),
    .o(o_rdwdata0[10]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1404 (
    .a(_al_u1133_o),
    .b(_al_u1200_o),
    .c(_al_u1134_o),
    .d(i_exu_op2[2]),
    .o(_al_u1404_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u1405 (
    .a(_al_u1060_o),
    .b(\u_EXU_ALU/n97_lutinv ),
    .c(_al_u1404_o),
    .d(_al_u954_o),
    .o(_al_u1405_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h155f))
    _al_u1406 (
    .a(i_decinfo[7]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[11]),
    .d(i_exu_op2[11]),
    .o(_al_u1406_o));
  AL_MAP_LUT5 #(
    .EQN("(E*B*~A*~(D*C))"),
    .INIT(32'h04440000))
    _al_u1407 (
    .a(alu2lsu_result[11]),
    .b(_al_u1406_o),
    .c(\u_EXU_ALU/n33 [11]),
    .d(i_decinfo[1]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1407_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u1408 (
    .a(\u_EXU_ALU/n256_lutinv ),
    .b(_al_u1108_o),
    .c(_al_u1319_o),
    .o(_al_u1408_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u1409 (
    .a(i_decinfo[5]),
    .b(i_exu_op1[11]),
    .c(i_exu_op2[11]),
    .o(\u_EXU_ALU/alu_xor [11]));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(C*A))"),
    .INIT(16'h004c))
    _al_u1410 (
    .a(_al_u1006_o),
    .b(_al_u1407_o),
    .c(_al_u1408_o),
    .d(\u_EXU_ALU/alu_xor [11]),
    .o(_al_u1410_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u1411 (
    .a(\u_EXU_ALU/n281_neg_lutinv ),
    .b(_al_u1063_o),
    .c(i_exu_op2[4]),
    .o(_al_u1411_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1412 (
    .a(bju_rdwdata[11]),
    .b(bju_rdwen),
    .c(i_csr_rdata[11]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1412_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(B*~(C*~(~E*A))))"),
    .INIT(32'h00f30073))
    _al_u1413 (
    .a(_al_u1405_o),
    .b(_al_u1410_o),
    .c(_al_u1411_o),
    .d(_al_u1412_o),
    .e(i_exu_op2[4]),
    .o(o_rdwdata0[11]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u1414 (
    .a(_al_u1124_o),
    .b(_al_u1185_o),
    .c(i_exu_op2[2]),
    .o(\u_EXU_ALU/n88_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'ha3))
    _al_u1415 (
    .a(\u_EXU_ALU/n125_lutinv ),
    .b(_al_u1322_o),
    .c(i_exu_op2[2]),
    .o(\u_EXU_ALU/n96_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u1416 (
    .a(\u_EXU_ALU/n88_lutinv ),
    .b(\u_EXU_ALU/n96_lutinv ),
    .c(_al_u1374_o),
    .d(i_exu_op2[3]),
    .o(_al_u1416_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*A*~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))"),
    .INIT(32'h0022000a))
    _al_u1417 (
    .a(_al_u1369_o),
    .b(_al_u1048_o),
    .c(_al_u1049_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u1417_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(D*~(~A*~(C)*~(E)+~A*C*~(E)+~(~A)*C*E+~A*C*E)))"),
    .INIT(32'h30331133))
    _al_u1418 (
    .a(\u_EXU_ALU/n372_lutinv ),
    .b(_al_u1417_o),
    .c(_al_u1045_o),
    .d(_al_u1026_o),
    .e(i_exu_op2[3]),
    .o(_al_u1418_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D*B)*~(C*A))"),
    .INIT(32'h135f5f5f))
    _al_u1419 (
    .a(\u_EXU_ALU/n33 [12]),
    .b(i_decinfo[6]),
    .c(i_decinfo[1]),
    .d(i_exu_op1[12]),
    .e(i_exu_op2[12]),
    .o(_al_u1419_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1420 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[12]),
    .d(i_exu_op2[12]),
    .o(_al_u1420_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~B*A*~(D*C))"),
    .INIT(32'h02220000))
    _al_u1421 (
    .a(_al_u1419_o),
    .b(_al_u1420_o),
    .c(\u_EXU_ALU/n0 [12]),
    .d(i_decinfo_grp[5]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1421_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1422 (
    .a(_al_u965_o),
    .b(i_exu_op1[31]),
    .o(\u_EXU_ALU/n249_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*D*C*B))"),
    .INIT(32'h2aaaaaaa))
    _al_u1423 (
    .a(_al_u1421_o),
    .b(_al_u1065_o),
    .c(_al_u961_o),
    .d(\u_EXU_ALU/n249_lutinv ),
    .e(i_exu_op2[4]),
    .o(_al_u1423_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1424 (
    .a(bju_rdwdata[12]),
    .b(bju_rdwen),
    .c(i_csr_rdata[12]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1424_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*~(D*~(B*~A))))"),
    .INIT(32'h0000bf0f))
    _al_u1425 (
    .a(_al_u1416_o),
    .b(_al_u1418_o),
    .c(_al_u1423_o),
    .d(\u_EXU_ALU/n281_neg_lutinv ),
    .e(_al_u1424_o),
    .o(o_rdwdata0[12]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1426 (
    .a(_al_u1233_o),
    .b(_al_u1261_o),
    .c(_al_u954_o),
    .d(i_exu_op2[2]),
    .o(_al_u1426_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)))"),
    .INIT(32'h50554455))
    _al_u1427 (
    .a(_al_u1426_o),
    .b(_al_u1179_o),
    .c(_al_u1180_o),
    .d(_al_u1134_o),
    .e(i_exu_op2[2]),
    .o(_al_u1427_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(~A*~(C)*~(D)+~A*C*~(D)+~(~A)*C*D+~A*C*D))"),
    .INIT(16'hc044))
    _al_u1428 (
    .a(_al_u1427_o),
    .b(\u_EXU_ALU/n281_neg_lutinv ),
    .c(\u_EXU_ALU/n46_lutinv ),
    .d(_al_u1323_o),
    .o(_al_u1428_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D*B)*~(C*A))"),
    .INIT(32'h135f5f5f))
    _al_u1429 (
    .a(\u_EXU_ALU/n33 [13]),
    .b(i_decinfo[6]),
    .c(i_decinfo[1]),
    .d(i_exu_op1[13]),
    .e(i_exu_op2[13]),
    .o(_al_u1429_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1430 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[13]),
    .d(i_exu_op2[13]),
    .o(_al_u1430_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*~A)"),
    .INIT(8'h04))
    _al_u1431 (
    .a(alu2lsu_result[13]),
    .b(_al_u1429_o),
    .c(_al_u1430_o),
    .o(_al_u1431_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(B*~A))"),
    .INIT(16'hb000))
    _al_u1432 (
    .a(_al_u1007_o),
    .b(_al_u965_o),
    .c(i_exu_op1[31]),
    .d(i_exu_op2[4]),
    .o(_al_u1432_o));
  AL_MAP_LUT4 #(
    .EQN("(D*B*~(C*A))"),
    .INIT(16'h4c00))
    _al_u1433 (
    .a(_al_u1066_o),
    .b(_al_u1431_o),
    .c(_al_u1432_o),
    .d(i_decinfo_grp[0]),
    .o(_al_u1433_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1434 (
    .a(bju_rdwdata[13]),
    .b(bju_rdwen),
    .c(i_csr_rdata[13]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1434_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(B*~A*~(D*~C)))"),
    .INIT(32'h0000bfbb))
    _al_u1435 (
    .a(_al_u1428_o),
    .b(_al_u1433_o),
    .c(_al_u1015_o),
    .d(_al_u1027_o),
    .e(_al_u1434_o),
    .o(o_rdwdata0[13]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(16'h50c0))
    _al_u1436 (
    .a(_al_u1217_o),
    .b(\u_EXU_ALU/n127_lutinv ),
    .c(_al_u954_o),
    .d(i_exu_op2[2]),
    .o(_al_u1436_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E)))"),
    .INIT(32'h11555055))
    _al_u1437 (
    .a(_al_u1436_o),
    .b(\u_EXU_ALU/n115_lutinv ),
    .c(_al_u1162_o),
    .d(_al_u1134_o),
    .e(i_exu_op2[2]),
    .o(_al_u1437_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(A*~(C*B)))"),
    .INIT(16'h00d5))
    _al_u1438 (
    .a(_al_u1437_o),
    .b(\u_EXU_ALU/n402_lutinv ),
    .c(i_decinfo[2]),
    .d(i_exu_op2[4]),
    .o(_al_u1438_o));
  AL_MAP_LUT5 #(
    .EQN("(D*B*A*~(~E*C))"),
    .INIT(32'h88000800))
    _al_u1439 (
    .a(\u_EXU_ALU/n179_neg_lutinv ),
    .b(_al_u1193_o),
    .c(_al_u965_o),
    .d(i_decinfo[4]),
    .e(i_exu_op2[1]),
    .o(_al_u1439_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D*B)*~(C*A))"),
    .INIT(32'h135f5f5f))
    _al_u1440 (
    .a(\u_EXU_ALU/n33 [14]),
    .b(i_decinfo[6]),
    .c(i_decinfo[1]),
    .d(i_exu_op1[14]),
    .e(i_exu_op2[14]),
    .o(_al_u1440_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u1441 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[14]),
    .d(i_exu_op2[14]),
    .o(_al_u1441_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u1442 (
    .a(alu2lsu_result[14]),
    .b(_al_u1440_o),
    .c(_al_u1441_o),
    .d(i_decinfo_grp[0]),
    .o(_al_u1442_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*A))"),
    .INIT(16'h4ccc))
    _al_u1443 (
    .a(\u_EXU_ALU/n281_neg_lutinv ),
    .b(_al_u1442_o),
    .c(\u_EXU_ALU/n45_lutinv ),
    .d(_al_u1323_o),
    .o(_al_u1443_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1444 (
    .a(bju_rdwdata[14]),
    .b(bju_rdwen),
    .c(i_csr_rdata[14]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1444_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*~B*~(D*A)))"),
    .INIT(32'h0000efcf))
    _al_u1445 (
    .a(_al_u1438_o),
    .b(_al_u1439_o),
    .c(_al_u1443_o),
    .d(\u_EXU_ALU/n281_neg_lutinv ),
    .e(_al_u1444_o),
    .o(o_rdwdata0[14]));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u1446 (
    .a(_al_u1200_o),
    .b(_al_u1301_o),
    .c(_al_u954_o),
    .d(i_exu_op2[2]),
    .o(_al_u1446_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)))"),
    .INIT(32'h50554455))
    _al_u1447 (
    .a(_al_u1446_o),
    .b(_al_u1133_o),
    .c(_al_u1061_o),
    .d(_al_u1134_o),
    .e(i_exu_op2[2]),
    .o(_al_u1447_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1448 (
    .a(\u_EXU_ALU/n77_lutinv ),
    .b(_al_u1369_o),
    .o(_al_u1448_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~E*~(A*~(D*~B))))"),
    .INIT(32'h0f0f080a))
    _al_u1449 (
    .a(_al_u1447_o),
    .b(_al_u907_o),
    .c(_al_u1448_o),
    .d(i_decinfo[2]),
    .e(i_exu_op2[4]),
    .o(_al_u1449_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u1450 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[15]),
    .c(i_exu_op2[15]),
    .o(\u_EXU_ALU/alu_and [15]));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(C*A))"),
    .INIT(16'h1300))
    _al_u1451 (
    .a(\u_EXU_ALU/n33 [15]),
    .b(\u_EXU_ALU/alu_and [15]),
    .c(i_decinfo[1]),
    .d(i_decinfo_grp[0]),
    .o(_al_u1451_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B*(D@C)))"),
    .INIT(16'ha22a))
    _al_u1452 (
    .a(_al_u1451_o),
    .b(i_decinfo[5]),
    .c(i_exu_op1[15]),
    .d(i_exu_op2[15]),
    .o(_al_u1452_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(B*~(~D*~C)))"),
    .INIT(16'h1115))
    _al_u1453 (
    .a(alu2lsu_result[15]),
    .b(i_decinfo[7]),
    .c(i_exu_op1[15]),
    .d(i_exu_op2[15]),
    .o(_al_u1453_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*~(~E*~D*A))"),
    .INIT(32'hc0c0c040))
    _al_u1454 (
    .a(_al_u948_o),
    .b(i_exu_op1[31]),
    .c(i_exu_op2[4]),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[0]),
    .o(_al_u1454_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*A))"),
    .INIT(16'h40c0))
    _al_u1455 (
    .a(_al_u1066_o),
    .b(_al_u1452_o),
    .c(_al_u1453_o),
    .d(_al_u1454_o),
    .o(_al_u1455_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u1456 (
    .a(bju_rdwdata[15]),
    .b(bju_rdwen),
    .c(i_csr_rdata[15]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u1456_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(C*~A)))"),
    .INIT(16'h0073))
    _al_u1457 (
    .a(_al_u1449_o),
    .b(_al_u1455_o),
    .c(\u_EXU_ALU/n281_neg_lutinv ),
    .d(_al_u1456_o),
    .o(o_rdwdata0[15]));
  AL_MAP_LUT5 #(
    .EQN("(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~(~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+~(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haa33aa0f))
    _al_u1458 (
    .a(_al_u1287_o),
    .b(i_exu_op1[5]),
    .c(i_exu_op1[4]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1458_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hffccaaf0))
    _al_u1459 (
    .a(i_exu_op1[2]),
    .b(i_exu_op1[1]),
    .c(i_exu_op1[0]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u1459_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(~D*C))*~(A)*~(E)+~(B*~(~D*C))*A*~(E)+~(~(B*~(~D*C)))*A*E+~(B*~(~D*C))*A*E)"),
    .INIT(32'h5555cc0c))
    _al_u1460 (
    .a(_al_u1458_o),
    .b(_al_u1459_o),
    .c(_al_u1007_o),
    .d(i_exu_op1[3]),
    .e(i_exu_op2[2]),
    .o(\u_EXU_ALU/n109_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~D*A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))"),
    .INIT(32'h008800a0))
    _al_u1461 (
    .a(\u_EXU_ALU/u1029_sel_is_0_o ),
    .b(\u_EXU_ALU/n101_lutinv ),
    .c(\u_EXU_ALU/n109_lutinv ),
    .d(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .e(i_exu_op2[3]),
    .o(_al_u1461_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u1462 (
    .a(\u_EXU_ALU/n253 ),
    .b(\u_EXU_ALU/n33 [0]),
    .c(i_decinfo[8]),
    .d(i_decinfo[1]),
    .o(_al_u1462_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(C*A))"),
    .INIT(16'h1300))
    _al_u1463 (
    .a(\u_EXU_ALU/n261 ),
    .b(alu2lsu_result[0]),
    .c(i_decinfo[9]),
    .d(i_decinfo_grp[0]),
    .o(_al_u1463_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u1464 (
    .a(\u_EXU_ALU/n352_lutinv ),
    .b(_al_u965_o),
    .o(\u_EXU_ALU/n416_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'heefafa00))
    _al_u1465 (
    .a(i_decinfo[7]),
    .b(i_decinfo[6]),
    .c(i_decinfo[5]),
    .d(i_exu_op1[0]),
    .e(i_exu_op2[0]),
    .o(_al_u1465_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*B*A*~(E*C))"),
    .INIT(32'h00080088))
    _al_u1466 (
    .a(_al_u1462_o),
    .b(_al_u1463_o),
    .c(\u_EXU_ALU/n416_lutinv ),
    .d(_al_u1465_o),
    .e(_al_u1027_o),
    .o(_al_u1466_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~((C*B)*~(E)*~(A)+(C*B)*E*~(A)+~((C*B))*E*A+(C*B)*E*A))"),
    .INIT(32'h001500bf))
    _al_u1467 (
    .a(bju_rdwen),
    .b(i_csr_rdata[0]),
    .c(i_decinfo_grp[4]),
    .d(i_decinfo_grp[0]),
    .e(i_iaddr[0]),
    .o(_al_u1467_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(B*~A*~(D*~C)))"),
    .INIT(32'h0000bfbb))
    _al_u1468 (
    .a(_al_u1461_o),
    .b(_al_u1466_o),
    .c(_al_u1249_o),
    .d(_al_u1392_o),
    .e(_al_u1467_o),
    .o(o_rdwdata0[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u386 (
    .a(i_decinfo[7]),
    .b(i_decinfo_grp[4]),
    .o(o_csr_wen));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u387 (
    .a(\u_EXU_ALU/n0 [0]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u388 (
    .a(\u_EXU_ALU/n0 [1]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u389 (
    .a(\u_EXU_BJU/bxx_nxtpc [0]),
    .b(i_decinfo[8]),
    .c(i_iaddr[0]),
    .o(o_exu_jaddr[0]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u390 (
    .a(\u_EXU_BJU/bxx_nxtpc [1]),
    .b(i_decinfo[8]),
    .c(i_iaddr[1]),
    .o(o_exu_jaddr[1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u391 (
    .a(\u_EXU_BJU/bxx_nxtpc [2]),
    .b(bju_rdwdata[2]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[2]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u392 (
    .a(\u_EXU_BJU/bxx_nxtpc [3]),
    .b(bju_rdwdata[3]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[3]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u393 (
    .a(\u_EXU_BJU/bxx_nxtpc [12]),
    .b(bju_rdwdata[12]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[12]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u394 (
    .a(\u_EXU_BJU/bxx_nxtpc [13]),
    .b(bju_rdwdata[13]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[13]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u395 (
    .a(\u_EXU_BJU/bxx_nxtpc [14]),
    .b(bju_rdwdata[14]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[14]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u396 (
    .a(\u_EXU_BJU/bxx_nxtpc [15]),
    .b(bju_rdwdata[15]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[15]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u397 (
    .a(\u_EXU_BJU/bxx_nxtpc [16]),
    .b(bju_rdwdata[16]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[16]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u398 (
    .a(\u_EXU_BJU/bxx_nxtpc [17]),
    .b(bju_rdwdata[17]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[17]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u399 (
    .a(\u_EXU_BJU/bxx_nxtpc [18]),
    .b(bju_rdwdata[18]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[18]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u400 (
    .a(\u_EXU_BJU/bxx_nxtpc [19]),
    .b(bju_rdwdata[19]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[19]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u401 (
    .a(\u_EXU_BJU/bxx_nxtpc [20]),
    .b(bju_rdwdata[20]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[20]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u402 (
    .a(\u_EXU_BJU/bxx_nxtpc [21]),
    .b(bju_rdwdata[21]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[21]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u403 (
    .a(\u_EXU_BJU/bxx_nxtpc [4]),
    .b(bju_rdwdata[4]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[4]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u404 (
    .a(\u_EXU_BJU/bxx_nxtpc [22]),
    .b(bju_rdwdata[22]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[22]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u405 (
    .a(\u_EXU_BJU/bxx_nxtpc [23]),
    .b(bju_rdwdata[23]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[23]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u406 (
    .a(\u_EXU_BJU/bxx_nxtpc [24]),
    .b(bju_rdwdata[24]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[24]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u407 (
    .a(\u_EXU_BJU/bxx_nxtpc [25]),
    .b(bju_rdwdata[25]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[25]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u408 (
    .a(\u_EXU_BJU/bxx_nxtpc [26]),
    .b(bju_rdwdata[26]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[26]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u409 (
    .a(\u_EXU_BJU/bxx_nxtpc [27]),
    .b(bju_rdwdata[27]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[27]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u410 (
    .a(\u_EXU_BJU/bxx_nxtpc [28]),
    .b(bju_rdwdata[28]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[28]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u411 (
    .a(\u_EXU_BJU/bxx_nxtpc [29]),
    .b(bju_rdwdata[29]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[29]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u412 (
    .a(\u_EXU_BJU/bxx_nxtpc [30]),
    .b(bju_rdwdata[30]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[30]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u413 (
    .a(\u_EXU_BJU/bxx_nxtpc [31]),
    .b(bju_rdwdata[31]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[31]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u414 (
    .a(\u_EXU_BJU/bxx_nxtpc [5]),
    .b(bju_rdwdata[5]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[5]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u415 (
    .a(\u_EXU_BJU/bxx_nxtpc [6]),
    .b(bju_rdwdata[6]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u416 (
    .a(\u_EXU_BJU/bxx_nxtpc [7]),
    .b(bju_rdwdata[7]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u417 (
    .a(\u_EXU_BJU/bxx_nxtpc [8]),
    .b(bju_rdwdata[8]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[8]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u418 (
    .a(\u_EXU_BJU/bxx_nxtpc [9]),
    .b(bju_rdwdata[9]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[9]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u419 (
    .a(\u_EXU_BJU/bxx_nxtpc [10]),
    .b(bju_rdwdata[10]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[10]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u420 (
    .a(\u_EXU_BJU/bxx_nxtpc [11]),
    .b(bju_rdwdata[11]),
    .c(i_decinfo[8]),
    .o(o_exu_jaddr[11]));
  AL_MAP_LUT2 #(
    .EQN("~(B*~A)"),
    .INIT(4'hb))
    _al_u421 (
    .a(i_ribm_rsp),
    .b(\u_EXU_LSU/handshake_rdy_last ),
    .o(\u_EXU_LSU/n1 ));
  AL_MAP_LUT4 #(
    .EQN("(D*A*~(C*~B))"),
    .INIT(16'h8a00))
    _al_u422 (
    .a(i_ribm_rsp),
    .b(\u_EXU_LSU/access2_once ),
    .c(\u_EXU_LSU/access2_vld ),
    .d(\u_EXU_LSU/handshake_rdy_last ),
    .o(_al_u422_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u423 (
    .a(_al_u422_o),
    .b(\u_EXU_LSU/access2_vld ),
    .c(o_exu_rdwen2),
    .o(o_rdwen2));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u424 (
    .a(i_decinfo[1]),
    .b(i_decinfo_grp[2]),
    .o(bju_rdwen));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*~A))"),
    .INIT(16'hfe00))
    _al_u425 (
    .a(bju_rdwen),
    .b(i_decinfo_grp[4]),
    .c(i_decinfo_grp[0]),
    .d(o_exu_rdwen0),
    .o(o_rdwen0));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55ff330f))
    _al_u426 (
    .a(i_ribm_rdata[26]),
    .b(i_ribm_rdata[10]),
    .c(i_ribm_rdata[2]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u426_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u427 (
    .a(\u_EXU_LSU/lsuinfo [2]),
    .b(\u_EXU_LSU/lsuinfo [3]),
    .o(\u_EXU_LSU/mux32_b0_sel_is_0_o ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u428 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u428_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u429 (
    .a(i_ribm_rdata[18]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(_al_u428_o),
    .o(_al_u429_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u430 (
    .a(i_ribm_rdata[2]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(_al_u430_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hea62))
    _al_u431 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/overleft_buffer [18]),
    .d(\u_EXU_LSU/overleft_buffer [26]),
    .o(_al_u431_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u432 (
    .a(\u_EXU_LSU/access2_vld ),
    .b(\u_EXU_LSU/lsuinfo [3]),
    .c(\u_EXU_LSU/lsuinfo [4]),
    .o(_al_u432_o));
  AL_MAP_LUT5 #(
    .EQN("(B*(A*C*~(D)*~(E)+A*~(C)*D*~(E)+A*C*D*~(E)+~(A)*~(C)*~(D)*E+A*C*~(D)*E+~(A)*~(C)*D*E+A*~(C)*D*E+A*C*D*E))"),
    .INIT(32'h8c848880))
    _al_u433 (
    .a(_al_u431_o),
    .b(_al_u432_o),
    .c(\u_EXU_LSU/align_mode_reg [1]),
    .d(\u_EXU_LSU/overleft_buffer [10]),
    .e(\u_EXU_LSU/overleft_buffer [2]),
    .o(_al_u433_o));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~(~E*~C*~(B*A)))"),
    .INIT(32'hff00ff07))
    _al_u434 (
    .a(_al_u426_o),
    .b(_al_u429_o),
    .c(_al_u430_o),
    .d(_al_u433_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[2]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55ff330f))
    _al_u435 (
    .a(i_ribm_rdata[27]),
    .b(i_ribm_rdata[11]),
    .c(i_ribm_rdata[3]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u435_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u436 (
    .a(i_ribm_rdata[19]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(_al_u428_o),
    .o(_al_u436_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u437 (
    .a(i_ribm_rdata[3]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(_al_u437_o));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hccb8))
    _al_u438 (
    .a(\u_EXU_LSU/overleft_buffer [19]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/overleft_buffer [3]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u438_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u439 (
    .a(\u_EXU_LSU/overleft_buffer [11]),
    .b(\u_EXU_LSU/overleft_buffer [27]),
    .c(_al_u438_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u439_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u440 (
    .a(_al_u439_o),
    .b(_al_u432_o),
    .o(_al_u440_o));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~(~E*~C*~(B*A)))"),
    .INIT(32'hff00ff07))
    _al_u441 (
    .a(_al_u435_o),
    .b(_al_u436_o),
    .c(_al_u437_o),
    .d(_al_u440_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[3]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55ff330f))
    _al_u442 (
    .a(i_ribm_rdata[28]),
    .b(i_ribm_rdata[12]),
    .c(i_ribm_rdata[4]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u442_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u443 (
    .a(i_ribm_rdata[20]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(_al_u428_o),
    .o(_al_u443_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u444 (
    .a(i_ribm_rdata[4]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(_al_u444_o));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hccb8))
    _al_u445 (
    .a(\u_EXU_LSU/overleft_buffer [20]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/overleft_buffer [4]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u445_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u446 (
    .a(\u_EXU_LSU/overleft_buffer [12]),
    .b(\u_EXU_LSU/overleft_buffer [28]),
    .c(_al_u445_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u446_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u447 (
    .a(_al_u446_o),
    .b(_al_u432_o),
    .o(_al_u447_o));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~(~E*~C*~(B*A)))"),
    .INIT(32'hff00ff07))
    _al_u448 (
    .a(_al_u442_o),
    .b(_al_u443_o),
    .c(_al_u444_o),
    .d(_al_u447_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[4]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55ff330f))
    _al_u449 (
    .a(i_ribm_rdata[29]),
    .b(i_ribm_rdata[13]),
    .c(i_ribm_rdata[5]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u449_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u450 (
    .a(i_ribm_rdata[21]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(_al_u428_o),
    .o(_al_u450_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u451 (
    .a(i_ribm_rdata[5]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u451_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~C*~(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)))"),
    .INIT(32'haaa2a8a0))
    _al_u452 (
    .a(_al_u432_o),
    .b(\u_EXU_LSU/align_mode_reg [0]),
    .c(\u_EXU_LSU/align_mode_reg [1]),
    .d(\u_EXU_LSU/overleft_buffer [13]),
    .e(\u_EXU_LSU/overleft_buffer [5]),
    .o(_al_u452_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u453 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/overleft_buffer [21]),
    .d(\u_EXU_LSU/overleft_buffer [29]),
    .o(_al_u453_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(~E*D)*~(C*~(B*A)))"),
    .INIT(32'h7070ff70))
    _al_u454 (
    .a(_al_u449_o),
    .b(_al_u450_o),
    .c(_al_u451_o),
    .d(_al_u452_o),
    .e(_al_u453_o),
    .o(o_rdwdata2[5]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55ff330f))
    _al_u455 (
    .a(i_ribm_rdata[30]),
    .b(i_ribm_rdata[14]),
    .c(i_ribm_rdata[6]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u455_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u456 (
    .a(i_ribm_rdata[22]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(_al_u428_o),
    .o(_al_u456_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u457 (
    .a(i_ribm_rdata[6]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(_al_u457_o));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hccb8))
    _al_u458 (
    .a(\u_EXU_LSU/overleft_buffer [22]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/overleft_buffer [6]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u458_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u459 (
    .a(\u_EXU_LSU/overleft_buffer [14]),
    .b(\u_EXU_LSU/overleft_buffer [30]),
    .c(_al_u458_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u459_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u460 (
    .a(_al_u459_o),
    .b(_al_u432_o),
    .o(_al_u460_o));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~(~E*~C*~(B*A)))"),
    .INIT(32'hff00ff07))
    _al_u461 (
    .a(_al_u455_o),
    .b(_al_u456_o),
    .c(_al_u457_o),
    .d(_al_u460_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[6]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haaffccf0))
    _al_u462 (
    .a(i_ribm_rdata[31]),
    .b(i_ribm_rdata[15]),
    .c(i_ribm_rdata[7]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u462_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u463 (
    .a(i_ribm_rdata[23]),
    .b(_al_u428_o),
    .o(_al_u463_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u464 (
    .a(i_ribm_rdata[7]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u464_o));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hccb8))
    _al_u465 (
    .a(\u_EXU_LSU/overleft_buffer [23]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/overleft_buffer [7]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u465_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u466 (
    .a(\u_EXU_LSU/overleft_buffer [15]),
    .b(\u_EXU_LSU/overleft_buffer [31]),
    .c(_al_u465_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u466_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u467 (
    .a(_al_u466_o),
    .b(_al_u432_o),
    .o(_al_u467_o));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~(C*~(~E*~(~B*A))))"),
    .INIT(32'hfff0ff20))
    _al_u468 (
    .a(_al_u462_o),
    .b(_al_u463_o),
    .c(_al_u464_o),
    .d(_al_u467_o),
    .e(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(o_rdwdata2[7]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55ff330f))
    _al_u469 (
    .a(i_ribm_rdata[24]),
    .b(i_ribm_rdata[8]),
    .c(i_ribm_rdata[0]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u469_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u470 (
    .a(i_ribm_rdata[16]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(_al_u428_o),
    .o(_al_u470_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u471 (
    .a(i_ribm_rdata[0]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(_al_u471_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'he6c4))
    _al_u472 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/overleft_buffer [24]),
    .d(\u_EXU_LSU/overleft_buffer [8]),
    .o(_al_u472_o));
  AL_MAP_LUT5 #(
    .EQN("(B*(A*C*~(D)*~(E)+~(A)*~(C)*D*~(E)+A*C*D*~(E)+A*~(C)*~(D)*E+A*C*~(D)*E+~(A)*~(C)*D*E+A*~(C)*D*E+A*C*D*E))"),
    .INIT(32'h8c888480))
    _al_u473 (
    .a(_al_u472_o),
    .b(_al_u432_o),
    .c(\u_EXU_LSU/align_mode_reg [0]),
    .d(\u_EXU_LSU/overleft_buffer [0]),
    .e(\u_EXU_LSU/overleft_buffer [16]),
    .o(_al_u473_o));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~(~E*~C*~(B*A)))"),
    .INIT(32'hff00ff07))
    _al_u474 (
    .a(_al_u469_o),
    .b(_al_u470_o),
    .c(_al_u471_o),
    .d(_al_u473_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[0]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55ff330f))
    _al_u475 (
    .a(i_ribm_rdata[25]),
    .b(i_ribm_rdata[9]),
    .c(i_ribm_rdata[1]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u475_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u476 (
    .a(i_ribm_rdata[17]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(_al_u428_o),
    .o(_al_u476_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u477 (
    .a(i_ribm_rdata[1]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(_al_u477_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'he6c4))
    _al_u478 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/overleft_buffer [25]),
    .d(\u_EXU_LSU/overleft_buffer [9]),
    .o(_al_u478_o));
  AL_MAP_LUT5 #(
    .EQN("(B*(A*C*~(D)*~(E)+~(A)*~(C)*D*~(E)+A*C*D*~(E)+A*~(C)*~(D)*E+A*C*~(D)*E+~(A)*~(C)*D*E+A*~(C)*D*E+A*C*D*E))"),
    .INIT(32'h8c888480))
    _al_u479 (
    .a(_al_u478_o),
    .b(_al_u432_o),
    .c(\u_EXU_LSU/align_mode_reg [0]),
    .d(\u_EXU_LSU/overleft_buffer [1]),
    .e(\u_EXU_LSU/overleft_buffer [17]),
    .o(_al_u479_o));
  AL_MAP_LUT5 #(
    .EQN("~(~D*~(~E*~C*~(B*A)))"),
    .INIT(32'hff00ff07))
    _al_u480 (
    .a(_al_u475_o),
    .b(_al_u476_o),
    .c(_al_u477_o),
    .d(_al_u479_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[1]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u481 (
    .a(i_decinfo[5]),
    .b(i_decinfo[4]),
    .o(_al_u481_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u482 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[31]),
    .c(i_csr_zimm[31]),
    .o(_al_u482_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u483 (
    .a(i_decinfo[4]),
    .b(i_decinfo[3]),
    .o(\u_EXU_LSU/mux14_b1_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(C)*~(B)+~(D*~A)*C*~(B)+~(~(D*~A))*C*B+~(D*~A)*C*B)"),
    .INIT(16'h1d0c))
    _al_u484 (
    .a(_al_u481_o),
    .b(_al_u482_o),
    .c(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .d(i_csr_rdata[31]),
    .o(o_csr_wdata[31]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u485 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[30]),
    .c(i_csr_zimm[30]),
    .o(_al_u485_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u486 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u485_o),
    .d(i_csr_rdata[30]),
    .o(o_csr_wdata[30]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u487 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[29]),
    .c(i_csr_zimm[29]),
    .o(_al_u487_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u488 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u487_o),
    .d(i_csr_rdata[29]),
    .o(o_csr_wdata[29]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u489 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[28]),
    .c(i_csr_zimm[28]),
    .o(_al_u489_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u490 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u489_o),
    .d(i_csr_rdata[28]),
    .o(o_csr_wdata[28]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u491 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[27]),
    .c(i_csr_zimm[27]),
    .o(_al_u491_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u492 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u491_o),
    .d(i_csr_rdata[27]),
    .o(o_csr_wdata[27]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u493 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[26]),
    .c(i_csr_zimm[26]),
    .o(_al_u493_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u494 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u493_o),
    .d(i_csr_rdata[26]),
    .o(o_csr_wdata[26]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u495 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[25]),
    .c(i_csr_zimm[25]),
    .o(_al_u495_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u496 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u495_o),
    .d(i_csr_rdata[25]),
    .o(o_csr_wdata[25]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u497 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[24]),
    .c(i_csr_zimm[24]),
    .o(_al_u497_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u498 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u497_o),
    .d(i_csr_rdata[24]),
    .o(o_csr_wdata[24]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u499 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[23]),
    .c(i_csr_zimm[23]),
    .o(_al_u499_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u500 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u499_o),
    .d(i_csr_rdata[23]),
    .o(o_csr_wdata[23]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u501 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[22]),
    .c(i_csr_zimm[22]),
    .o(_al_u501_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u502 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u501_o),
    .d(i_csr_rdata[22]),
    .o(o_csr_wdata[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u503 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[21]),
    .c(i_csr_zimm[21]),
    .o(_al_u503_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u504 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u503_o),
    .d(i_csr_rdata[21]),
    .o(o_csr_wdata[21]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u505 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[20]),
    .c(i_csr_zimm[20]),
    .o(_al_u505_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u506 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u505_o),
    .d(i_csr_rdata[20]),
    .o(o_csr_wdata[20]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u507 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[19]),
    .c(i_csr_zimm[19]),
    .o(_al_u507_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u508 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u507_o),
    .d(i_csr_rdata[19]),
    .o(o_csr_wdata[19]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u509 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[18]),
    .c(i_csr_zimm[18]),
    .o(_al_u509_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u510 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u509_o),
    .d(i_csr_rdata[18]),
    .o(o_csr_wdata[18]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u511 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[17]),
    .c(i_csr_zimm[17]),
    .o(_al_u511_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u512 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u511_o),
    .d(i_csr_rdata[17]),
    .o(o_csr_wdata[17]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u513 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[16]),
    .c(i_csr_zimm[16]),
    .o(_al_u513_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u514 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u513_o),
    .d(i_csr_rdata[16]),
    .o(o_csr_wdata[16]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u515 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[15]),
    .c(i_csr_zimm[15]),
    .o(_al_u515_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u516 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u515_o),
    .d(i_csr_rdata[15]),
    .o(o_csr_wdata[15]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u517 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[14]),
    .c(i_csr_zimm[14]),
    .o(_al_u517_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u518 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u517_o),
    .d(i_csr_rdata[14]),
    .o(o_csr_wdata[14]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u519 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[13]),
    .c(i_csr_zimm[13]),
    .o(_al_u519_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u520 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u519_o),
    .d(i_csr_rdata[13]),
    .o(o_csr_wdata[13]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u521 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[12]),
    .c(i_csr_zimm[12]),
    .o(_al_u521_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u522 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u521_o),
    .d(i_csr_rdata[12]),
    .o(o_csr_wdata[12]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u523 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[11]),
    .c(i_csr_zimm[11]),
    .o(_al_u523_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u524 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u523_o),
    .d(i_csr_rdata[11]),
    .o(o_csr_wdata[11]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u525 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[10]),
    .c(i_csr_zimm[10]),
    .o(_al_u525_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u526 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u525_o),
    .d(i_csr_rdata[10]),
    .o(o_csr_wdata[10]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u527 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[9]),
    .c(i_csr_zimm[9]),
    .o(_al_u527_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u528 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u527_o),
    .d(i_csr_rdata[9]),
    .o(o_csr_wdata[9]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u529 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[8]),
    .c(i_csr_zimm[8]),
    .o(_al_u529_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u530 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u529_o),
    .d(i_csr_rdata[8]),
    .o(o_csr_wdata[8]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u531 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[7]),
    .c(i_csr_zimm[7]),
    .o(_al_u531_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u532 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u531_o),
    .d(i_csr_rdata[7]),
    .o(o_csr_wdata[7]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u533 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[6]),
    .c(i_csr_zimm[6]),
    .o(_al_u533_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u534 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u533_o),
    .d(i_csr_rdata[6]),
    .o(o_csr_wdata[6]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u535 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[5]),
    .c(i_csr_zimm[5]),
    .o(_al_u535_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~A)*~(B)*~(C)+~(D*~A)*B*~(C)+~(~(D*~A))*B*C+~(D*~A)*B*C)"),
    .INIT(16'h3530))
    _al_u536 (
    .a(_al_u481_o),
    .b(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .c(_al_u535_o),
    .d(i_csr_rdata[5]),
    .o(o_csr_wdata[5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u537 (
    .a(i_csr_zimm[4]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[4]),
    .o(_al_u537_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~B)*~(C)*~(A)+~(D*~B)*C*~(A)+~(~(D*~B))*C*A+~(D*~B)*C*A)"),
    .INIT(16'h1b0a))
    _al_u538 (
    .a(_al_u537_o),
    .b(_al_u481_o),
    .c(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .d(i_csr_rdata[4]),
    .o(o_csr_wdata[4]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u539 (
    .a(i_csr_zimm[3]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[3]),
    .o(_al_u539_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~B)*~(C)*~(A)+~(D*~B)*C*~(A)+~(~(D*~B))*C*A+~(D*~B)*C*A)"),
    .INIT(16'h1b0a))
    _al_u540 (
    .a(_al_u539_o),
    .b(_al_u481_o),
    .c(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .d(i_csr_rdata[3]),
    .o(o_csr_wdata[3]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u541 (
    .a(i_csr_zimm[2]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[2]),
    .o(_al_u541_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~B)*~(C)*~(A)+~(D*~B)*C*~(A)+~(~(D*~B))*C*A+~(D*~B)*C*A)"),
    .INIT(16'h1b0a))
    _al_u542 (
    .a(_al_u541_o),
    .b(_al_u481_o),
    .c(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .d(i_csr_rdata[2]),
    .o(o_csr_wdata[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u543 (
    .a(i_csr_zimm[1]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[1]),
    .o(_al_u543_o));
  AL_MAP_LUT4 #(
    .EQN("~(~(D*~B)*~(C)*~(A)+~(D*~B)*C*~(A)+~(~(D*~B))*C*A+~(D*~B)*C*A)"),
    .INIT(16'h1b0a))
    _al_u544 (
    .a(_al_u543_o),
    .b(_al_u481_o),
    .c(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .d(i_csr_rdata[1]),
    .o(o_csr_wdata[1]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'h47))
    _al_u545 (
    .a(i_csr_zimm[0]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[0]),
    .o(\u_EXU_SCU/n0 [0]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~((D*~B))*~(A)+~C*(D*~B)*~(A)+~(~C)*(D*~B)*A+~C*(D*~B)*A)"),
    .INIT(16'h2705))
    _al_u546 (
    .a(\u_EXU_SCU/n0 [0]),
    .b(_al_u481_o),
    .c(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .d(i_csr_rdata[0]),
    .o(o_csr_wdata[0]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D*A*~(C*~B)))"),
    .INIT(32'h75ff0000))
    _al_u547 (
    .a(i_ribm_rsp),
    .b(\u_EXU_LSU/access2_once ),
    .c(\u_EXU_LSU/access2_vld ),
    .d(\u_EXU_LSU/handshake_rdy_last ),
    .e(\u_EXU_LSU/working ),
    .o(o_lsu_working));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff55330f))
    _al_u548 (
    .a(i_ribm_rdata[25]),
    .b(i_ribm_rdata[17]),
    .c(i_ribm_rdata[9]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u548_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(A)*~(D)+~(~C*B)*A*~(D)+~(~(~C*B))*A*D+~(~C*B)*A*D)"),
    .INIT(16'haaf3))
    _al_u549 (
    .a(_al_u548_o),
    .b(i_ribm_rdata[9]),
    .c(\u_EXU_LSU/lsuinfo [2]),
    .d(\u_EXU_LSU/lsuinfo [3]),
    .o(_al_u549_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u550 (
    .a(i_ribm_rdata[15]),
    .b(i_ribm_rdata[7]),
    .c(\u_EXU_LSU/align_mode_reg [0]),
    .d(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u550_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u551 (
    .a(\u_EXU_LSU/lsuinfo [2]),
    .b(\u_EXU_LSU/lsuinfo [3]),
    .c(\u_EXU_LSU/lsuinfo [5]),
    .o(_al_u551_o));
  AL_MAP_LUT5 #(
    .EQN("(D*(A*~(B)*~(C)*~(E)+A*B*~(C)*~(E)+A*~(B)*C*~(E)+A*B*C*~(E)+A*B*~(C)*E+~(A)*~(B)*C*E+~(A)*B*C*E+A*B*C*E))"),
    .INIT(32'hd800aa00))
    _al_u552 (
    .a(_al_u550_o),
    .b(i_ribm_rdata[31]),
    .c(i_ribm_rdata[23]),
    .d(_al_u551_o),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u552_o));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haad8))
    _al_u553 (
    .a(\u_EXU_LSU/align_mode_reg [1]),
    .b(\u_EXU_LSU/overleft_buffer [25]),
    .c(\u_EXU_LSU/overleft_buffer [9]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u553_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u554 (
    .a(i_ribm_rdata[1]),
    .b(\u_EXU_LSU/overleft_buffer [17]),
    .c(_al_u553_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/access2_data [9]));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*C)*~(~E*~(~B*A)))"),
    .INIT(32'hf000fddd))
    _al_u555 (
    .a(_al_u549_o),
    .b(_al_u552_o),
    .c(\u_EXU_LSU/access2_data [9]),
    .d(_al_u432_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[9]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff55330f))
    _al_u556 (
    .a(i_ribm_rdata[24]),
    .b(i_ribm_rdata[16]),
    .c(i_ribm_rdata[8]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u556_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(A)*~(D)+~(~C*B)*A*~(D)+~(~(~C*B))*A*D+~(~C*B)*A*D)"),
    .INIT(16'haaf3))
    _al_u557 (
    .a(_al_u556_o),
    .b(i_ribm_rdata[8]),
    .c(\u_EXU_LSU/lsuinfo [2]),
    .d(\u_EXU_LSU/lsuinfo [3]),
    .o(_al_u557_o));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haad8))
    _al_u558 (
    .a(\u_EXU_LSU/align_mode_reg [1]),
    .b(\u_EXU_LSU/overleft_buffer [24]),
    .c(\u_EXU_LSU/overleft_buffer [8]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u558_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u559 (
    .a(i_ribm_rdata[0]),
    .b(\u_EXU_LSU/overleft_buffer [16]),
    .c(_al_u558_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/access2_data [8]));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*C)*~(~E*~(~B*A)))"),
    .INIT(32'hf000fddd))
    _al_u560 (
    .a(_al_u557_o),
    .b(_al_u552_o),
    .c(\u_EXU_LSU/access2_data [8]),
    .d(_al_u432_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u561 (
    .a(\u_EXU_LSU/align_mode_reg [1]),
    .b(\u_EXU_LSU/lsuinfo [4]),
    .o(_al_u561_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u562 (
    .a(i_ribm_rdata[23]),
    .b(i_ribm_rdata[15]),
    .c(_al_u561_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u562_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u563 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/overleft_buffer [15]),
    .c(\u_EXU_LSU/overleft_buffer [23]),
    .o(_al_u563_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~((E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C))*~(D)+~B*(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*~(D)+~(~B)*(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*D+~B*(E*~(A)*~(C)+E*A*~(C)+~(E)*A*C+E*A*C)*D)"),
    .INIT(32'haf33a033))
    _al_u564 (
    .a(i_ribm_rdata[7]),
    .b(_al_u563_o),
    .c(\u_EXU_LSU/align_mode_reg [0]),
    .d(\u_EXU_LSU/align_mode_reg [1]),
    .e(\u_EXU_LSU/overleft_buffer [31]),
    .o(\u_EXU_LSU/access2_data [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u565 (
    .a(\u_EXU_LSU/align_mode_reg [1]),
    .b(\u_EXU_LSU/lsuinfo [4]),
    .o(_al_u565_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u566 (
    .a(i_ribm_rdata[7]),
    .b(_al_u565_o),
    .c(\u_EXU_LSU/align_mode_reg [0]),
    .d(\u_EXU_LSU/overleft_buffer [31]),
    .o(_al_u566_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u567 (
    .a(\u_EXU_LSU/lsuinfo [3]),
    .b(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/mux16_b3_sel_is_2_o ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u568 (
    .a(\u_EXU_LSU/mux16_b3_sel_is_2_o ),
    .b(\u_EXU_LSU/lsuinfo [5]),
    .o(_al_u568_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~C*~A*~(D*B))"),
    .INIT(32'h01050000))
    _al_u569 (
    .a(_al_u562_o),
    .b(\u_EXU_LSU/access2_data [15]),
    .c(_al_u566_o),
    .d(_al_u568_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(_al_u569_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff55330f))
    _al_u570 (
    .a(i_ribm_rdata[31]),
    .b(i_ribm_rdata[23]),
    .c(i_ribm_rdata[15]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u570_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u571 (
    .a(i_ribm_rdata[31]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u571_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u572 (
    .a(\u_EXU_LSU/lsuinfo [3]),
    .b(\u_EXU_LSU/lsuinfo [5]),
    .o(\u_EXU_LSU/mux27_b16_sel_is_1_o ));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~B*~(E*~C)))"),
    .INIT(32'h45554455))
    _al_u573 (
    .a(_al_u569_o),
    .b(_al_u552_o),
    .c(_al_u570_o),
    .d(_al_u571_o),
    .e(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .o(o_rdwdata2[31]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'h5f003f00))
    _al_u574 (
    .a(i_ribm_rdata[22]),
    .b(i_ribm_rdata[14]),
    .c(_al_u561_o),
    .d(\u_EXU_LSU/access2_vld ),
    .e(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u574_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u575 (
    .a(i_ribm_rdata[6]),
    .b(_al_u565_o),
    .c(\u_EXU_LSU/align_mode_reg [0]),
    .d(\u_EXU_LSU/overleft_buffer [30]),
    .o(_al_u575_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u576 (
    .a(_al_u574_o),
    .b(\u_EXU_LSU/access2_data [15]),
    .c(_al_u575_o),
    .d(_al_u568_o),
    .o(_al_u576_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u577 (
    .a(i_ribm_rdata[30]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u577_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~B*~(E*~C)))"),
    .INIT(32'h45554455))
    _al_u578 (
    .a(_al_u576_o),
    .b(_al_u552_o),
    .c(_al_u570_o),
    .d(_al_u577_o),
    .e(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .o(o_rdwdata2[30]));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u579 (
    .a(i_ribm_rdata[21]),
    .b(i_ribm_rdata[13]),
    .c(_al_u561_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u579_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u580 (
    .a(i_ribm_rdata[5]),
    .b(_al_u565_o),
    .c(\u_EXU_LSU/align_mode_reg [0]),
    .d(\u_EXU_LSU/overleft_buffer [29]),
    .o(_al_u580_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~C*~A*~(D*B))"),
    .INIT(32'h01050000))
    _al_u581 (
    .a(_al_u579_o),
    .b(\u_EXU_LSU/access2_data [15]),
    .c(_al_u580_o),
    .d(_al_u568_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(_al_u581_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u582 (
    .a(i_ribm_rdata[29]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u582_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~B*~(E*~C)))"),
    .INIT(32'h45554455))
    _al_u583 (
    .a(_al_u581_o),
    .b(_al_u552_o),
    .c(_al_u570_o),
    .d(_al_u582_o),
    .e(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .o(o_rdwdata2[29]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'h5f003f00))
    _al_u584 (
    .a(i_ribm_rdata[20]),
    .b(i_ribm_rdata[12]),
    .c(_al_u561_o),
    .d(\u_EXU_LSU/access2_vld ),
    .e(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u584_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u585 (
    .a(i_ribm_rdata[4]),
    .b(_al_u565_o),
    .c(\u_EXU_LSU/align_mode_reg [0]),
    .d(\u_EXU_LSU/overleft_buffer [28]),
    .o(_al_u585_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u586 (
    .a(_al_u584_o),
    .b(\u_EXU_LSU/access2_data [15]),
    .c(_al_u585_o),
    .d(_al_u568_o),
    .o(_al_u586_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u587 (
    .a(i_ribm_rdata[28]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u587_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~B*~(E*~C)))"),
    .INIT(32'h45554455))
    _al_u588 (
    .a(_al_u586_o),
    .b(_al_u552_o),
    .c(_al_u570_o),
    .d(_al_u587_o),
    .e(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .o(o_rdwdata2[28]));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u589 (
    .a(i_ribm_rdata[19]),
    .b(i_ribm_rdata[11]),
    .c(_al_u561_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u589_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u590 (
    .a(i_ribm_rdata[3]),
    .b(_al_u565_o),
    .c(\u_EXU_LSU/align_mode_reg [0]),
    .d(\u_EXU_LSU/overleft_buffer [27]),
    .o(_al_u590_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~C*~A*~(D*B))"),
    .INIT(32'h01050000))
    _al_u591 (
    .a(_al_u589_o),
    .b(\u_EXU_LSU/access2_data [15]),
    .c(_al_u590_o),
    .d(_al_u568_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(_al_u591_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u592 (
    .a(i_ribm_rdata[27]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u592_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~B*~(E*~C)))"),
    .INIT(32'h45554455))
    _al_u593 (
    .a(_al_u591_o),
    .b(_al_u552_o),
    .c(_al_u570_o),
    .d(_al_u592_o),
    .e(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .o(o_rdwdata2[27]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(C*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'h5f003f00))
    _al_u594 (
    .a(i_ribm_rdata[18]),
    .b(i_ribm_rdata[10]),
    .c(_al_u561_o),
    .d(\u_EXU_LSU/access2_vld ),
    .e(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u594_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u595 (
    .a(i_ribm_rdata[2]),
    .b(_al_u565_o),
    .c(\u_EXU_LSU/align_mode_reg [0]),
    .d(\u_EXU_LSU/overleft_buffer [26]),
    .o(_al_u595_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u596 (
    .a(_al_u594_o),
    .b(\u_EXU_LSU/access2_data [15]),
    .c(_al_u595_o),
    .d(_al_u568_o),
    .o(_al_u596_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u597 (
    .a(i_ribm_rdata[26]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u597_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~B*~(E*~C)))"),
    .INIT(32'h45554455))
    _al_u598 (
    .a(_al_u596_o),
    .b(_al_u552_o),
    .c(_al_u570_o),
    .d(_al_u597_o),
    .e(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .o(o_rdwdata2[26]));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u599 (
    .a(i_ribm_rdata[17]),
    .b(i_ribm_rdata[9]),
    .c(_al_u561_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u599_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u600 (
    .a(i_ribm_rdata[1]),
    .b(_al_u565_o),
    .c(\u_EXU_LSU/align_mode_reg [0]),
    .d(\u_EXU_LSU/overleft_buffer [25]),
    .o(_al_u600_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~C*~A*~(D*B))"),
    .INIT(32'h01050000))
    _al_u601 (
    .a(_al_u599_o),
    .b(\u_EXU_LSU/access2_data [15]),
    .c(_al_u600_o),
    .d(_al_u568_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(_al_u601_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u602 (
    .a(i_ribm_rdata[25]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u602_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~B*~(E*~C)))"),
    .INIT(32'h45554455))
    _al_u603 (
    .a(_al_u601_o),
    .b(_al_u552_o),
    .c(_al_u570_o),
    .d(_al_u602_o),
    .e(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .o(o_rdwdata2[25]));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u604 (
    .a(i_ribm_rdata[16]),
    .b(i_ribm_rdata[8]),
    .c(_al_u561_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u604_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u605 (
    .a(i_ribm_rdata[0]),
    .b(_al_u565_o),
    .c(\u_EXU_LSU/align_mode_reg [0]),
    .d(\u_EXU_LSU/overleft_buffer [24]),
    .o(_al_u605_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~C*~A*~(D*B))"),
    .INIT(32'h01050000))
    _al_u606 (
    .a(_al_u604_o),
    .b(\u_EXU_LSU/access2_data [15]),
    .c(_al_u605_o),
    .d(_al_u568_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(_al_u606_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u607 (
    .a(i_ribm_rdata[24]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u607_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*~B*~(E*~C)))"),
    .INIT(32'h45554455))
    _al_u608 (
    .a(_al_u606_o),
    .b(_al_u552_o),
    .c(_al_u570_o),
    .d(_al_u607_o),
    .e(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .o(o_rdwdata2[24]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u609 (
    .a(_al_u570_o),
    .b(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u609_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u610 (
    .a(\u_EXU_LSU/access2_data [15]),
    .b(_al_u568_o),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u610_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u611 (
    .a(_al_u565_o),
    .b(\u_EXU_LSU/align_mode_reg [0]),
    .c(\u_EXU_LSU/overleft_buffer [23]),
    .d(\u_EXU_LSU/overleft_buffer [31]),
    .o(_al_u611_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'h050f030f))
    _al_u612 (
    .a(i_ribm_rdata[15]),
    .b(i_ribm_rdata[7]),
    .c(_al_u611_o),
    .d(_al_u561_o),
    .e(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u612_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u613 (
    .a(i_ribm_rdata[23]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(_al_u613_o));
  AL_MAP_LUT5 #(
    .EQN("(~(D*C)*~(~E*~B*A))"),
    .INIT(32'h0fff0ddd))
    _al_u614 (
    .a(_al_u609_o),
    .b(_al_u552_o),
    .c(_al_u610_o),
    .d(_al_u612_o),
    .e(_al_u613_o),
    .o(o_rdwdata2[23]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u615 (
    .a(_al_u565_o),
    .b(\u_EXU_LSU/align_mode_reg [0]),
    .c(\u_EXU_LSU/overleft_buffer [22]),
    .d(\u_EXU_LSU/overleft_buffer [30]),
    .o(_al_u615_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'h050f030f))
    _al_u616 (
    .a(i_ribm_rdata[14]),
    .b(i_ribm_rdata[6]),
    .c(_al_u615_o),
    .d(_al_u561_o),
    .e(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u616_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u617 (
    .a(i_ribm_rdata[22]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(_al_u617_o));
  AL_MAP_LUT5 #(
    .EQN("(~(D*C)*~(~E*~B*A))"),
    .INIT(32'h0fff0ddd))
    _al_u618 (
    .a(_al_u609_o),
    .b(_al_u552_o),
    .c(_al_u610_o),
    .d(_al_u616_o),
    .e(_al_u617_o),
    .o(o_rdwdata2[22]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*B)*~(D*~A))"),
    .INIT(32'h00002a3f))
    _al_u619 (
    .a(_al_u570_o),
    .b(i_ribm_rdata[21]),
    .c(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .d(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .e(\u_EXU_LSU/access2_vld ),
    .o(_al_u619_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haae4))
    _al_u620 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/overleft_buffer [21]),
    .c(\u_EXU_LSU/overleft_buffer [29]),
    .d(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u620_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u621 (
    .a(i_ribm_rdata[13]),
    .b(i_ribm_rdata[5]),
    .c(_al_u620_o),
    .d(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/access2_data [21]));
  AL_MAP_LUT5 #(
    .EQN("(~(~(E*D)*C)*~(~B*A))"),
    .INIT(32'hdd0d0d0d))
    _al_u622 (
    .a(_al_u619_o),
    .b(_al_u552_o),
    .c(_al_u610_o),
    .d(\u_EXU_LSU/access2_data [21]),
    .e(\u_EXU_LSU/lsuinfo [4]),
    .o(o_rdwdata2[21]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u623 (
    .a(_al_u565_o),
    .b(\u_EXU_LSU/align_mode_reg [0]),
    .c(\u_EXU_LSU/overleft_buffer [20]),
    .d(\u_EXU_LSU/overleft_buffer [28]),
    .o(_al_u623_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'h050f030f))
    _al_u624 (
    .a(i_ribm_rdata[12]),
    .b(i_ribm_rdata[4]),
    .c(_al_u623_o),
    .d(_al_u561_o),
    .e(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u624_o));
  AL_MAP_LUT4 #(
    .EQN("(D*A*~(C*B))"),
    .INIT(16'h2a00))
    _al_u625 (
    .a(_al_u624_o),
    .b(\u_EXU_LSU/access2_data [15]),
    .c(_al_u568_o),
    .d(\u_EXU_LSU/access2_vld ),
    .o(_al_u625_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u626 (
    .a(i_ribm_rdata[20]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u626_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(D*~A*~(E*~C)))"),
    .INIT(32'h23332233))
    _al_u627 (
    .a(_al_u552_o),
    .b(_al_u625_o),
    .c(_al_u570_o),
    .d(_al_u626_o),
    .e(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .o(o_rdwdata2[20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u628 (
    .a(_al_u565_o),
    .b(\u_EXU_LSU/align_mode_reg [0]),
    .c(\u_EXU_LSU/overleft_buffer [19]),
    .d(\u_EXU_LSU/overleft_buffer [27]),
    .o(_al_u628_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'h050f030f))
    _al_u629 (
    .a(i_ribm_rdata[11]),
    .b(i_ribm_rdata[3]),
    .c(_al_u628_o),
    .d(_al_u561_o),
    .e(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u629_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u630 (
    .a(i_ribm_rdata[19]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(_al_u630_o));
  AL_MAP_LUT5 #(
    .EQN("(~(D*C)*~(~E*~B*A))"),
    .INIT(32'h0fff0ddd))
    _al_u631 (
    .a(_al_u609_o),
    .b(_al_u552_o),
    .c(_al_u610_o),
    .d(_al_u629_o),
    .e(_al_u630_o),
    .o(o_rdwdata2[19]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u632 (
    .a(_al_u565_o),
    .b(\u_EXU_LSU/align_mode_reg [0]),
    .c(\u_EXU_LSU/overleft_buffer [18]),
    .d(\u_EXU_LSU/overleft_buffer [26]),
    .o(_al_u632_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'h050f030f))
    _al_u633 (
    .a(i_ribm_rdata[10]),
    .b(i_ribm_rdata[2]),
    .c(_al_u632_o),
    .d(_al_u561_o),
    .e(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u633_o));
  AL_MAP_LUT4 #(
    .EQN("(D*A*~(C*B))"),
    .INIT(16'h2a00))
    _al_u634 (
    .a(_al_u633_o),
    .b(\u_EXU_LSU/access2_data [15]),
    .c(_al_u568_o),
    .d(\u_EXU_LSU/access2_vld ),
    .o(_al_u634_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u635 (
    .a(i_ribm_rdata[18]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u635_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(D*~A*~(E*~C)))"),
    .INIT(32'h23332233))
    _al_u636 (
    .a(_al_u552_o),
    .b(_al_u634_o),
    .c(_al_u570_o),
    .d(_al_u635_o),
    .e(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .o(o_rdwdata2[18]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u637 (
    .a(_al_u565_o),
    .b(\u_EXU_LSU/align_mode_reg [0]),
    .c(\u_EXU_LSU/overleft_buffer [17]),
    .d(\u_EXU_LSU/overleft_buffer [25]),
    .o(_al_u637_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'h050f030f))
    _al_u638 (
    .a(i_ribm_rdata[9]),
    .b(i_ribm_rdata[1]),
    .c(_al_u637_o),
    .d(_al_u561_o),
    .e(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u638_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u639 (
    .a(i_ribm_rdata[17]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .o(_al_u639_o));
  AL_MAP_LUT5 #(
    .EQN("(~(D*C)*~(~E*~B*A))"),
    .INIT(32'h0fff0ddd))
    _al_u640 (
    .a(_al_u609_o),
    .b(_al_u552_o),
    .c(_al_u610_o),
    .d(_al_u638_o),
    .e(_al_u639_o),
    .o(o_rdwdata2[17]));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u641 (
    .a(_al_u565_o),
    .b(\u_EXU_LSU/align_mode_reg [0]),
    .c(\u_EXU_LSU/overleft_buffer [16]),
    .d(\u_EXU_LSU/overleft_buffer [24]),
    .o(_al_u641_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*(B*~(A)*~(E)+B*A*~(E)+~(B)*A*E+B*A*E)))"),
    .INIT(32'h050f030f))
    _al_u642 (
    .a(i_ribm_rdata[8]),
    .b(i_ribm_rdata[0]),
    .c(_al_u641_o),
    .d(_al_u561_o),
    .e(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u642_o));
  AL_MAP_LUT4 #(
    .EQN("(D*A*~(C*B))"),
    .INIT(16'h2a00))
    _al_u643 (
    .a(_al_u642_o),
    .b(\u_EXU_LSU/access2_data [15]),
    .c(_al_u568_o),
    .d(\u_EXU_LSU/access2_vld ),
    .o(_al_u643_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u644 (
    .a(i_ribm_rdata[16]),
    .b(\u_EXU_LSU/mux32_b0_sel_is_0_o ),
    .c(\u_EXU_LSU/access2_vld ),
    .o(_al_u644_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(D*~A*~(E*~C)))"),
    .INIT(32'h23332233))
    _al_u645 (
    .a(_al_u552_o),
    .b(_al_u643_o),
    .c(_al_u570_o),
    .d(_al_u644_o),
    .e(\u_EXU_LSU/mux27_b16_sel_is_1_o ),
    .o(o_rdwdata2[16]));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(A)*~(D)+~(~C*B)*A*~(D)+~(~(~C*B))*A*D+~(~C*B)*A*D)"),
    .INIT(16'haaf3))
    _al_u646 (
    .a(_al_u570_o),
    .b(i_ribm_rdata[15]),
    .c(\u_EXU_LSU/lsuinfo [2]),
    .d(\u_EXU_LSU/lsuinfo [3]),
    .o(_al_u646_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*C)*~(~E*~(~B*A)))"),
    .INIT(32'hf000fddd))
    _al_u647 (
    .a(_al_u646_o),
    .b(_al_u552_o),
    .c(\u_EXU_LSU/access2_data [15]),
    .d(_al_u432_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[15]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff55330f))
    _al_u648 (
    .a(i_ribm_rdata[30]),
    .b(i_ribm_rdata[22]),
    .c(i_ribm_rdata[14]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u648_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(A)*~(D)+~(~C*B)*A*~(D)+~(~(~C*B))*A*D+~(~C*B)*A*D)"),
    .INIT(16'haaf3))
    _al_u649 (
    .a(_al_u648_o),
    .b(i_ribm_rdata[14]),
    .c(\u_EXU_LSU/lsuinfo [2]),
    .d(\u_EXU_LSU/lsuinfo [3]),
    .o(_al_u649_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcce2))
    _al_u650 (
    .a(\u_EXU_LSU/overleft_buffer [14]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/overleft_buffer [30]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u650_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u651 (
    .a(i_ribm_rdata[6]),
    .b(\u_EXU_LSU/overleft_buffer [22]),
    .c(_al_u650_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/access2_data [14]));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*C)*~(~E*~(~B*A)))"),
    .INIT(32'hf000fddd))
    _al_u652 (
    .a(_al_u649_o),
    .b(_al_u552_o),
    .c(\u_EXU_LSU/access2_data [14]),
    .d(_al_u432_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[14]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff55330f))
    _al_u653 (
    .a(i_ribm_rdata[29]),
    .b(i_ribm_rdata[21]),
    .c(i_ribm_rdata[13]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u653_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(A)*~(D)+~(~C*B)*A*~(D)+~(~(~C*B))*A*D+~(~C*B)*A*D)"),
    .INIT(16'haaf3))
    _al_u654 (
    .a(_al_u653_o),
    .b(i_ribm_rdata[13]),
    .c(\u_EXU_LSU/lsuinfo [2]),
    .d(\u_EXU_LSU/lsuinfo [3]),
    .o(_al_u654_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u655 (
    .a(i_ribm_rdata[5]),
    .b(\u_EXU_LSU/align_mode_reg [0]),
    .c(\u_EXU_LSU/overleft_buffer [29]),
    .o(\u_EXU_LSU/n155_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u656 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/overleft_buffer [13]),
    .c(\u_EXU_LSU/overleft_buffer [21]),
    .o(_al_u656_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .INIT(16'h880c))
    _al_u657 (
    .a(\u_EXU_LSU/n155_lutinv ),
    .b(_al_u432_o),
    .c(_al_u656_o),
    .d(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u657_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(~D*~(~B*A)))"),
    .INIT(16'hf0fd))
    _al_u658 (
    .a(_al_u654_o),
    .b(_al_u552_o),
    .c(_al_u657_o),
    .d(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[13]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff55330f))
    _al_u659 (
    .a(i_ribm_rdata[28]),
    .b(i_ribm_rdata[20]),
    .c(i_ribm_rdata[12]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u659_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(A)*~(D)+~(~C*B)*A*~(D)+~(~(~C*B))*A*D+~(~C*B)*A*D)"),
    .INIT(16'haaf3))
    _al_u660 (
    .a(_al_u659_o),
    .b(i_ribm_rdata[12]),
    .c(\u_EXU_LSU/lsuinfo [2]),
    .d(\u_EXU_LSU/lsuinfo [3]),
    .o(_al_u660_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcce2))
    _al_u661 (
    .a(\u_EXU_LSU/overleft_buffer [12]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/overleft_buffer [28]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u661_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u662 (
    .a(i_ribm_rdata[4]),
    .b(\u_EXU_LSU/overleft_buffer [20]),
    .c(_al_u661_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(\u_EXU_LSU/access2_data [12]));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*C)*~(~E*~(~B*A)))"),
    .INIT(32'hf000fddd))
    _al_u663 (
    .a(_al_u660_o),
    .b(_al_u552_o),
    .c(\u_EXU_LSU/access2_data [12]),
    .d(_al_u432_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[12]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff55330f))
    _al_u664 (
    .a(i_ribm_rdata[27]),
    .b(i_ribm_rdata[19]),
    .c(i_ribm_rdata[11]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u664_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(A)*~(D)+~(~C*B)*A*~(D)+~(~(~C*B))*A*D+~(~C*B)*A*D)"),
    .INIT(16'haaf3))
    _al_u665 (
    .a(_al_u664_o),
    .b(i_ribm_rdata[11]),
    .c(\u_EXU_LSU/lsuinfo [2]),
    .d(\u_EXU_LSU/lsuinfo [3]),
    .o(_al_u665_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'hb8))
    _al_u666 (
    .a(i_ribm_rdata[3]),
    .b(\u_EXU_LSU/align_mode_reg [0]),
    .c(\u_EXU_LSU/overleft_buffer [27]),
    .o(\u_EXU_LSU/n157_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u667 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/overleft_buffer [11]),
    .c(\u_EXU_LSU/overleft_buffer [19]),
    .o(_al_u667_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(~C*~(A)*~(D)+~C*A*~(D)+~(~C)*A*D+~C*A*D))"),
    .INIT(16'h880c))
    _al_u668 (
    .a(\u_EXU_LSU/n157_lutinv ),
    .b(_al_u432_o),
    .c(_al_u667_o),
    .d(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u668_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(~D*~(~B*A)))"),
    .INIT(16'hf0fd))
    _al_u669 (
    .a(_al_u665_o),
    .b(_al_u552_o),
    .c(_al_u668_o),
    .d(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[11]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff55330f))
    _al_u670 (
    .a(i_ribm_rdata[26]),
    .b(i_ribm_rdata[18]),
    .c(i_ribm_rdata[10]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .e(\u_EXU_LSU/align_mode_reg [1]),
    .o(_al_u670_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(A)*~(D)+~(~C*B)*A*~(D)+~(~(~C*B))*A*D+~(~C*B)*A*D)"),
    .INIT(16'haaf3))
    _al_u671 (
    .a(_al_u670_o),
    .b(i_ribm_rdata[10]),
    .c(\u_EXU_LSU/lsuinfo [2]),
    .d(\u_EXU_LSU/lsuinfo [3]),
    .o(_al_u671_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcce2))
    _al_u672 (
    .a(\u_EXU_LSU/overleft_buffer [10]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/overleft_buffer [26]),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u672_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h530f))
    _al_u673 (
    .a(i_ribm_rdata[2]),
    .b(\u_EXU_LSU/overleft_buffer [18]),
    .c(_al_u672_o),
    .d(\u_EXU_LSU/align_mode_reg [0]),
    .o(_al_u673_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(D*~C)*~(~E*~(~B*A)))"),
    .INIT(32'h0f00dfdd))
    _al_u674 (
    .a(_al_u671_o),
    .b(_al_u552_o),
    .c(_al_u673_o),
    .d(_al_u432_o),
    .e(\u_EXU_LSU/access2_vld ),
    .o(o_rdwdata2[10]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u675 (
    .a(o_rdidx0[4]),
    .b(o_rdidx0[3]),
    .c(o_exu_rdidx1[4]),
    .d(o_exu_rdidx1[3]),
    .o(_al_u675_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u676 (
    .a(o_rdidx0[1]),
    .b(o_rdidx0[0]),
    .c(o_exu_rdidx1[1]),
    .d(o_exu_rdidx1[0]),
    .o(_al_u676_o));
  AL_MAP_LUT4 #(
    .EQN("(D*B*~(C@A))"),
    .INIT(16'h8400))
    _al_u677 (
    .a(o_rdidx0[2]),
    .b(o_exu_rdwen0),
    .c(o_exu_rdidx1[2]),
    .d(o_exu_rdwen1),
    .o(_al_u677_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u678 (
    .a(_al_u675_o),
    .b(_al_u676_o),
    .c(_al_u677_o),
    .o(mdu_flush));
  AL_MAP_LUT4 #(
    .EQN("~(~(C*B)*~(D*A))"),
    .INIT(16'heac0))
    _al_u679 (
    .a(o_lsu_working),
    .b(o_mdu_working),
    .c(i_decinfo_grp[3]),
    .d(i_decinfo_grp[1]),
    .o(o_exu_resource_match));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u680 (
    .a(i_vld),
    .b(o_lsu_working),
    .c(i_decinfo_grp[1]),
    .o(_al_u680_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*C*~(D)+~(A)*~(C)*D+~(A)*C*D))"),
    .INIT(16'h1120))
    _al_u681 (
    .a(i_ribm_gnt),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/access2_vld ),
    .d(\u_EXU_LSU/handshake_once ),
    .o(\u_EXU_LSU/n80 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u682 (
    .a(_al_u422_o),
    .b(\u_EXU_LSU/access2_vld ),
    .o(\u_EXU_LSU/n20_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h171f))
    _al_u683 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_decinfo[4]),
    .d(i_decinfo[3]),
    .o(_al_u683_o));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(C)*~((E*~D*A))+~B*C*~((E*~D*A))+~(~B)*C*(E*~D*A)+~B*C*(E*~D*A))"),
    .INIT(32'hcc4ecccc))
    _al_u684 (
    .a(i_vld),
    .b(\u_EXU_LSU/n20_lutinv ),
    .c(_al_u683_o),
    .d(o_lsu_working),
    .e(i_decinfo_grp[1]),
    .o(\u_EXU_LSU/n26 ));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    _al_u685 (
    .a(i_vld),
    .b(o_lsu_working),
    .c(i_decinfo_grp[1]),
    .o(\u_EXU_LSU/n25 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u686 (
    .a(\u_EXU_LSU/access2_vld ),
    .b(\u_EXU_LSU/handshake_once ),
    .o(\u_EXU_LSU/n57 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u687 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n57 ),
    .o(_al_u687_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u688 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[9]),
    .d(i_rs2rdata[1]),
    .o(\u_EXU_LSU/n55 [9]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u689 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [17]),
    .d(\u_EXU_LSU/rs2rdata_reg [25]),
    .o(\u_EXU_LSU/n67 [9]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u690 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [9]),
    .d(\u_EXU_LSU/n67 [9]),
    .e(o_ribm_wdata[9]),
    .o(\u_EXU_LSU/n79 [9]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u691 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[8]),
    .d(i_rs2rdata[0]),
    .o(\u_EXU_LSU/n55 [8]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u692 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [16]),
    .d(\u_EXU_LSU/rs2rdata_reg [24]),
    .o(\u_EXU_LSU/n67 [8]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u693 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [8]),
    .d(\u_EXU_LSU/n67 [8]),
    .e(o_ribm_wdata[8]),
    .o(\u_EXU_LSU/n79 [8]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u694 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[7]),
    .o(\u_EXU_LSU/n55 [7]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E)"),
    .INIT(32'h195d3b7f))
    _al_u695 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [15]),
    .d(\u_EXU_LSU/rs2rdata_reg [23]),
    .e(\u_EXU_LSU/rs2rdata_reg [31]),
    .o(_al_u695_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*~(C)*~(B)+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*~(B)+~(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A))*C*B+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*B)"),
    .INIT(32'hd1f3c0e2))
    _al_u696 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [7]),
    .d(_al_u695_o),
    .e(o_ribm_wdata[7]),
    .o(\u_EXU_LSU/n79 [7]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u697 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[6]),
    .o(\u_EXU_LSU/n55 [6]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E)"),
    .INIT(32'h195d3b7f))
    _al_u698 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [14]),
    .d(\u_EXU_LSU/rs2rdata_reg [22]),
    .e(\u_EXU_LSU/rs2rdata_reg [30]),
    .o(_al_u698_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*~(C)*~(B)+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*~(B)+~(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A))*C*B+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*B)"),
    .INIT(32'hd1f3c0e2))
    _al_u699 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [6]),
    .d(_al_u698_o),
    .e(o_ribm_wdata[6]),
    .o(\u_EXU_LSU/n79 [6]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u700 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[5]),
    .o(\u_EXU_LSU/n55 [5]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E)"),
    .INIT(32'h195d3b7f))
    _al_u701 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [13]),
    .d(\u_EXU_LSU/rs2rdata_reg [21]),
    .e(\u_EXU_LSU/rs2rdata_reg [29]),
    .o(_al_u701_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*~(C)*~(B)+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*~(B)+~(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A))*C*B+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*B)"),
    .INIT(32'hd1f3c0e2))
    _al_u702 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [5]),
    .d(_al_u701_o),
    .e(o_ribm_wdata[5]),
    .o(\u_EXU_LSU/n79 [5]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u703 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[4]),
    .o(\u_EXU_LSU/n55 [4]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E)"),
    .INIT(32'h195d3b7f))
    _al_u704 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [12]),
    .d(\u_EXU_LSU/rs2rdata_reg [20]),
    .e(\u_EXU_LSU/rs2rdata_reg [28]),
    .o(_al_u704_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*~(C)*~(B)+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*~(B)+~(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A))*C*B+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*B)"),
    .INIT(32'hd1f3c0e2))
    _al_u705 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [4]),
    .d(_al_u704_o),
    .e(o_ribm_wdata[4]),
    .o(\u_EXU_LSU/n79 [4]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hd8aa))
    _al_u706 (
    .a(alu2lsu_result[0]),
    .b(i_rs2rdata[7]),
    .c(i_rs2rdata[15]),
    .d(alu2lsu_result[1]),
    .o(_al_u706_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u707 (
    .a(i_rs2rdata[31]),
    .b(i_rs2rdata[23]),
    .c(_al_u706_o),
    .d(alu2lsu_result[1]),
    .o(_al_u707_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D*A))*~(C)*~(B)+~(E*~(D*A))*C*~(B)+~(~(E*~(D*A)))*C*B+~(E*~(D*A))*C*B)"),
    .INIT(32'h1d3f0c0c))
    _al_u708 (
    .a(i_ribm_gnt),
    .b(_al_u680_o),
    .c(_al_u707_o),
    .d(\u_EXU_LSU/n57 ),
    .e(o_ribm_wdata[31]),
    .o(\u_EXU_LSU/n79 [31]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hd8aa))
    _al_u709 (
    .a(alu2lsu_result[0]),
    .b(i_rs2rdata[6]),
    .c(i_rs2rdata[14]),
    .d(alu2lsu_result[1]),
    .o(_al_u709_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u710 (
    .a(i_rs2rdata[30]),
    .b(i_rs2rdata[22]),
    .c(_al_u709_o),
    .d(alu2lsu_result[1]),
    .o(_al_u710_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D*A))*~(C)*~(B)+~(E*~(D*A))*C*~(B)+~(~(E*~(D*A)))*C*B+~(E*~(D*A))*C*B)"),
    .INIT(32'h1d3f0c0c))
    _al_u711 (
    .a(i_ribm_gnt),
    .b(_al_u680_o),
    .c(_al_u710_o),
    .d(\u_EXU_LSU/n57 ),
    .e(o_ribm_wdata[30]),
    .o(\u_EXU_LSU/n79 [30]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u712 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[3]),
    .o(\u_EXU_LSU/n55 [3]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E)"),
    .INIT(32'h195d3b7f))
    _al_u713 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [11]),
    .d(\u_EXU_LSU/rs2rdata_reg [19]),
    .e(\u_EXU_LSU/rs2rdata_reg [27]),
    .o(_al_u713_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*~(C)*~(B)+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*~(B)+~(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A))*C*B+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*B)"),
    .INIT(32'hd1f3c0e2))
    _al_u714 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [3]),
    .d(_al_u713_o),
    .e(o_ribm_wdata[3]),
    .o(\u_EXU_LSU/n79 [3]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hd8aa))
    _al_u715 (
    .a(alu2lsu_result[0]),
    .b(i_rs2rdata[5]),
    .c(i_rs2rdata[13]),
    .d(alu2lsu_result[1]),
    .o(_al_u715_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u716 (
    .a(i_rs2rdata[29]),
    .b(i_rs2rdata[21]),
    .c(_al_u715_o),
    .d(alu2lsu_result[1]),
    .o(_al_u716_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D*A))*~(C)*~(B)+~(E*~(D*A))*C*~(B)+~(~(E*~(D*A)))*C*B+~(E*~(D*A))*C*B)"),
    .INIT(32'h1d3f0c0c))
    _al_u717 (
    .a(i_ribm_gnt),
    .b(_al_u680_o),
    .c(_al_u716_o),
    .d(\u_EXU_LSU/n57 ),
    .e(o_ribm_wdata[29]),
    .o(\u_EXU_LSU/n79 [29]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hd8aa))
    _al_u718 (
    .a(alu2lsu_result[0]),
    .b(i_rs2rdata[4]),
    .c(i_rs2rdata[12]),
    .d(alu2lsu_result[1]),
    .o(_al_u718_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u719 (
    .a(i_rs2rdata[28]),
    .b(i_rs2rdata[20]),
    .c(_al_u718_o),
    .d(alu2lsu_result[1]),
    .o(_al_u719_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D*A))*~(C)*~(B)+~(E*~(D*A))*C*~(B)+~(~(E*~(D*A)))*C*B+~(E*~(D*A))*C*B)"),
    .INIT(32'h1d3f0c0c))
    _al_u720 (
    .a(i_ribm_gnt),
    .b(_al_u680_o),
    .c(_al_u719_o),
    .d(\u_EXU_LSU/n57 ),
    .e(o_ribm_wdata[28]),
    .o(\u_EXU_LSU/n79 [28]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hd8aa))
    _al_u721 (
    .a(alu2lsu_result[0]),
    .b(i_rs2rdata[3]),
    .c(i_rs2rdata[11]),
    .d(alu2lsu_result[1]),
    .o(_al_u721_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u722 (
    .a(i_rs2rdata[27]),
    .b(i_rs2rdata[19]),
    .c(_al_u721_o),
    .d(alu2lsu_result[1]),
    .o(_al_u722_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D*A))*~(C)*~(B)+~(E*~(D*A))*C*~(B)+~(~(E*~(D*A)))*C*B+~(E*~(D*A))*C*B)"),
    .INIT(32'h1d3f0c0c))
    _al_u723 (
    .a(i_ribm_gnt),
    .b(_al_u680_o),
    .c(_al_u722_o),
    .d(\u_EXU_LSU/n57 ),
    .e(o_ribm_wdata[27]),
    .o(\u_EXU_LSU/n79 [27]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hd8aa))
    _al_u724 (
    .a(alu2lsu_result[0]),
    .b(i_rs2rdata[2]),
    .c(i_rs2rdata[10]),
    .d(alu2lsu_result[1]),
    .o(_al_u724_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u725 (
    .a(i_rs2rdata[26]),
    .b(i_rs2rdata[18]),
    .c(_al_u724_o),
    .d(alu2lsu_result[1]),
    .o(_al_u725_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D*A))*~(C)*~(B)+~(E*~(D*A))*C*~(B)+~(~(E*~(D*A)))*C*B+~(E*~(D*A))*C*B)"),
    .INIT(32'h1d3f0c0c))
    _al_u726 (
    .a(i_ribm_gnt),
    .b(_al_u680_o),
    .c(_al_u725_o),
    .d(\u_EXU_LSU/n57 ),
    .e(o_ribm_wdata[26]),
    .o(\u_EXU_LSU/n79 [26]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hd8aa))
    _al_u727 (
    .a(alu2lsu_result[0]),
    .b(i_rs2rdata[1]),
    .c(i_rs2rdata[9]),
    .d(alu2lsu_result[1]),
    .o(_al_u727_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u728 (
    .a(i_rs2rdata[25]),
    .b(i_rs2rdata[17]),
    .c(_al_u727_o),
    .d(alu2lsu_result[1]),
    .o(_al_u728_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D*A))*~(C)*~(B)+~(E*~(D*A))*C*~(B)+~(~(E*~(D*A)))*C*B+~(E*~(D*A))*C*B)"),
    .INIT(32'h1d3f0c0c))
    _al_u729 (
    .a(i_ribm_gnt),
    .b(_al_u680_o),
    .c(_al_u728_o),
    .d(\u_EXU_LSU/n57 ),
    .e(o_ribm_wdata[25]),
    .o(\u_EXU_LSU/n79 [25]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hd8aa))
    _al_u730 (
    .a(alu2lsu_result[0]),
    .b(i_rs2rdata[0]),
    .c(i_rs2rdata[8]),
    .d(alu2lsu_result[1]),
    .o(_al_u730_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u731 (
    .a(i_rs2rdata[24]),
    .b(i_rs2rdata[16]),
    .c(_al_u730_o),
    .d(alu2lsu_result[1]),
    .o(_al_u731_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D*A))*~(C)*~(B)+~(E*~(D*A))*C*~(B)+~(~(E*~(D*A)))*C*B+~(E*~(D*A))*C*B)"),
    .INIT(32'h1d3f0c0c))
    _al_u732 (
    .a(i_ribm_gnt),
    .b(_al_u680_o),
    .c(_al_u731_o),
    .d(\u_EXU_LSU/n57 ),
    .e(o_ribm_wdata[24]),
    .o(\u_EXU_LSU/n79 [24]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h89cdabef))
    _al_u733 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[23]),
    .d(i_rs2rdata[15]),
    .e(i_rs2rdata[7]),
    .o(_al_u733_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u734 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [31]),
    .o(\u_EXU_LSU/n67 [23]));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'h3f1d2e0c))
    _al_u735 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(_al_u733_o),
    .d(\u_EXU_LSU/n67 [23]),
    .e(o_ribm_wdata[23]),
    .o(\u_EXU_LSU/n79 [23]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h89cdabef))
    _al_u736 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[22]),
    .d(i_rs2rdata[14]),
    .e(i_rs2rdata[6]),
    .o(_al_u736_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u737 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [30]),
    .o(\u_EXU_LSU/n67 [22]));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'h3f1d2e0c))
    _al_u738 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(_al_u736_o),
    .d(\u_EXU_LSU/n67 [22]),
    .e(o_ribm_wdata[22]),
    .o(\u_EXU_LSU/n79 [22]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h89cdabef))
    _al_u739 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[21]),
    .d(i_rs2rdata[13]),
    .e(i_rs2rdata[5]),
    .o(_al_u739_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u740 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [29]),
    .o(\u_EXU_LSU/n67 [21]));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'h3f1d2e0c))
    _al_u741 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(_al_u739_o),
    .d(\u_EXU_LSU/n67 [21]),
    .e(o_ribm_wdata[21]),
    .o(\u_EXU_LSU/n79 [21]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h89cdabef))
    _al_u742 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[20]),
    .d(i_rs2rdata[12]),
    .e(i_rs2rdata[4]),
    .o(_al_u742_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u743 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [28]),
    .o(\u_EXU_LSU/n67 [20]));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'h3f1d2e0c))
    _al_u744 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(_al_u742_o),
    .d(\u_EXU_LSU/n67 [20]),
    .e(o_ribm_wdata[20]),
    .o(\u_EXU_LSU/n79 [20]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u745 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[2]),
    .o(\u_EXU_LSU/n55 [2]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E)"),
    .INIT(32'h195d3b7f))
    _al_u746 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [10]),
    .d(\u_EXU_LSU/rs2rdata_reg [18]),
    .e(\u_EXU_LSU/rs2rdata_reg [26]),
    .o(_al_u746_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*~(C)*~(B)+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*~(B)+~(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A))*C*B+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*B)"),
    .INIT(32'hd1f3c0e2))
    _al_u747 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [2]),
    .d(_al_u746_o),
    .e(o_ribm_wdata[2]),
    .o(\u_EXU_LSU/n79 [2]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h89cdabef))
    _al_u748 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[19]),
    .d(i_rs2rdata[11]),
    .e(i_rs2rdata[3]),
    .o(_al_u748_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u749 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [27]),
    .o(\u_EXU_LSU/n67 [19]));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'h3f1d2e0c))
    _al_u750 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(_al_u748_o),
    .d(\u_EXU_LSU/n67 [19]),
    .e(o_ribm_wdata[19]),
    .o(\u_EXU_LSU/n79 [19]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h89cdabef))
    _al_u751 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[18]),
    .d(i_rs2rdata[10]),
    .e(i_rs2rdata[2]),
    .o(_al_u751_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u752 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [26]),
    .o(\u_EXU_LSU/n67 [18]));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'h3f1d2e0c))
    _al_u753 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(_al_u751_o),
    .d(\u_EXU_LSU/n67 [18]),
    .e(o_ribm_wdata[18]),
    .o(\u_EXU_LSU/n79 [18]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h89cdabef))
    _al_u754 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[17]),
    .d(i_rs2rdata[9]),
    .e(i_rs2rdata[1]),
    .o(_al_u754_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u755 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [25]),
    .o(\u_EXU_LSU/n67 [17]));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'h3f1d2e0c))
    _al_u756 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(_al_u754_o),
    .d(\u_EXU_LSU/n67 [17]),
    .e(o_ribm_wdata[17]),
    .o(\u_EXU_LSU/n79 [17]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h89cdabef))
    _al_u757 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[16]),
    .d(i_rs2rdata[8]),
    .e(i_rs2rdata[0]),
    .o(_al_u757_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u758 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [24]),
    .o(\u_EXU_LSU/n67 [16]));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~(~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'h3f1d2e0c))
    _al_u759 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(_al_u757_o),
    .d(\u_EXU_LSU/n67 [16]),
    .e(o_ribm_wdata[16]),
    .o(\u_EXU_LSU/n79 [16]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u760 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[15]),
    .d(i_rs2rdata[7]),
    .o(\u_EXU_LSU/n55 [15]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u761 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [23]),
    .d(\u_EXU_LSU/rs2rdata_reg [31]),
    .o(\u_EXU_LSU/n67 [15]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u762 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [15]),
    .d(\u_EXU_LSU/n67 [15]),
    .e(o_ribm_wdata[15]),
    .o(\u_EXU_LSU/n79 [15]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u763 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[14]),
    .d(i_rs2rdata[6]),
    .o(\u_EXU_LSU/n55 [14]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u764 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [22]),
    .d(\u_EXU_LSU/rs2rdata_reg [30]),
    .o(\u_EXU_LSU/n67 [14]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u765 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [14]),
    .d(\u_EXU_LSU/n67 [14]),
    .e(o_ribm_wdata[14]),
    .o(\u_EXU_LSU/n79 [14]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u766 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[13]),
    .d(i_rs2rdata[5]),
    .o(\u_EXU_LSU/n55 [13]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u767 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [21]),
    .d(\u_EXU_LSU/rs2rdata_reg [29]),
    .o(\u_EXU_LSU/n67 [13]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u768 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [13]),
    .d(\u_EXU_LSU/n67 [13]),
    .e(o_ribm_wdata[13]),
    .o(\u_EXU_LSU/n79 [13]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u769 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[12]),
    .d(i_rs2rdata[4]),
    .o(\u_EXU_LSU/n55 [12]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u770 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [20]),
    .d(\u_EXU_LSU/rs2rdata_reg [28]),
    .o(\u_EXU_LSU/n67 [12]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u771 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [12]),
    .d(\u_EXU_LSU/n67 [12]),
    .e(o_ribm_wdata[12]),
    .o(\u_EXU_LSU/n79 [12]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u772 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[11]),
    .d(i_rs2rdata[3]),
    .o(\u_EXU_LSU/n55 [11]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u773 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [19]),
    .d(\u_EXU_LSU/rs2rdata_reg [27]),
    .o(\u_EXU_LSU/n67 [11]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u774 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [11]),
    .d(\u_EXU_LSU/n67 [11]),
    .e(o_ribm_wdata[11]),
    .o(\u_EXU_LSU/n79 [11]));
  AL_MAP_LUT4 #(
    .EQN("(~A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h5410))
    _al_u775 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[10]),
    .d(i_rs2rdata[2]),
    .o(\u_EXU_LSU/n55 [10]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u776 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [18]),
    .d(\u_EXU_LSU/rs2rdata_reg [26]),
    .o(\u_EXU_LSU/n67 [10]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u777 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [10]),
    .d(\u_EXU_LSU/n67 [10]),
    .e(o_ribm_wdata[10]),
    .o(\u_EXU_LSU/n79 [10]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u778 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[1]),
    .o(\u_EXU_LSU/n55 [1]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E)"),
    .INIT(32'h15379dbf))
    _al_u779 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [17]),
    .d(\u_EXU_LSU/rs2rdata_reg [25]),
    .e(\u_EXU_LSU/rs2rdata_reg [9]),
    .o(_al_u779_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*~(C)*~(B)+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*~(B)+~(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A))*C*B+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*B)"),
    .INIT(32'hd1f3c0e2))
    _al_u780 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [1]),
    .d(_al_u779_o),
    .e(o_ribm_wdata[1]),
    .o(\u_EXU_LSU/n79 [1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u781 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_rs2rdata[0]),
    .o(\u_EXU_LSU/n55 [0]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E)"),
    .INIT(32'h15379dbf))
    _al_u782 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/rs2rdata_reg [16]),
    .d(\u_EXU_LSU/rs2rdata_reg [24]),
    .e(\u_EXU_LSU/rs2rdata_reg [8]),
    .o(_al_u782_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*~(C)*~(B)+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*~(B)+~(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A))*C*B+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*B)"),
    .INIT(32'hd1f3c0e2))
    _al_u783 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n55 [0]),
    .d(_al_u782_o),
    .e(o_ribm_wdata[0]),
    .o(\u_EXU_LSU/n79 [0]));
  AL_MAP_LUT5 #(
    .EQN("(~(~(E*B)*C)*~(~D*~A))"),
    .INIT(32'hcf8a0f0a))
    _al_u784 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .d(i_decinfo[4]),
    .e(i_decinfo[2]),
    .o(\u_EXU_LSU/n54 [3]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u785 (
    .a(\u_EXU_LSU/mux16_b3_sel_is_2_o ),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .o(\u_EXU_LSU/n65 [3]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u786 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n54 [3]),
    .d(\u_EXU_LSU/n65 [3]),
    .e(o_ribm_mask[3]),
    .o(\u_EXU_LSU/n78 [3]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h76727670))
    _al_u787 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(i_decinfo[4]),
    .d(i_decinfo[3]),
    .e(i_decinfo[2]),
    .o(\u_EXU_LSU/n54 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h776f))
    _al_u788 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/lsuinfo [3]),
    .d(\u_EXU_LSU/lsuinfo [4]),
    .o(_al_u788_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*~(C)*~(B)+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*~(B)+~(~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A))*C*B+~(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)*C*B)"),
    .INIT(32'hd1f3c0e2))
    _al_u789 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n54 [2]),
    .d(_al_u788_o),
    .e(o_ribm_mask[2]),
    .o(\u_EXU_LSU/n78 [2]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D*B)))"),
    .INIT(16'h4505))
    _al_u790 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .d(i_decinfo[2]),
    .o(\u_EXU_LSU/n54 [1]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u791 (
    .a(\u_EXU_LSU/align_mode_reg [1]),
    .b(\u_EXU_LSU/lsuinfo [3]),
    .c(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n65 [1]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u792 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n54 [1]),
    .d(\u_EXU_LSU/n65 [1]),
    .e(o_ribm_mask[1]),
    .o(\u_EXU_LSU/n78 [1]));
  AL_MAP_LUT4 #(
    .EQN("(~(~D*~C)*~(~B*~A))"),
    .INIT(16'heee0))
    _al_u793 (
    .a(\u_EXU_LSU/align_mode_reg [0]),
    .b(\u_EXU_LSU/align_mode_reg [1]),
    .c(\u_EXU_LSU/lsuinfo [3]),
    .d(\u_EXU_LSU/lsuinfo [4]),
    .o(\u_EXU_LSU/n65 [0]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u794 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n65 [0]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_mask[0]),
    .o(_al_u794_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*~(~D*C))"),
    .INIT(16'h1101))
    _al_u795 (
    .a(alu2lsu_result[1]),
    .b(alu2lsu_result[0]),
    .c(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .d(i_decinfo[2]),
    .o(\u_EXU_LSU/n54 [0]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u796 (
    .a(_al_u794_o),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n54 [0]),
    .o(\u_EXU_LSU/n78 [0]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u797 (
    .a(\u_EXU_ALU/n0 [9]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[9]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u798 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[9]),
    .d(\u_EXU_LSU/n59 [7]),
    .e(o_ribm_addr[9]),
    .o(\u_EXU_LSU/n76 [9]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u799 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [6]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[8]),
    .o(_al_u799_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u800 (
    .a(_al_u799_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [8]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [8]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u801 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [5]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[7]),
    .o(_al_u801_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u802 (
    .a(_al_u801_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [7]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u803 (
    .a(\u_EXU_ALU/n0 [6]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[6]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u804 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[6]),
    .d(\u_EXU_LSU/n59 [4]),
    .e(o_ribm_addr[6]),
    .o(\u_EXU_LSU/n76 [6]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u805 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [3]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[5]),
    .o(_al_u805_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u806 (
    .a(_al_u805_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [5]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [5]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u807 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [2]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[4]),
    .o(_al_u807_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u808 (
    .a(_al_u807_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [4]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [4]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u809 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [29]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[31]),
    .o(_al_u809_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u810 (
    .a(_al_u809_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [31]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [31]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u811 (
    .a(\u_EXU_ALU/n0 [30]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[30]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u812 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[30]),
    .d(\u_EXU_LSU/n59 [28]),
    .e(o_ribm_addr[30]),
    .o(\u_EXU_LSU/n76 [30]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u813 (
    .a(\u_EXU_ALU/n0 [3]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[3]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u814 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[3]),
    .d(\u_EXU_LSU/n59 [1]),
    .e(o_ribm_addr[3]),
    .o(\u_EXU_LSU/n76 [3]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u815 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [27]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[29]),
    .o(_al_u815_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u816 (
    .a(_al_u815_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [29]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [29]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u817 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [26]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[28]),
    .o(_al_u817_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u818 (
    .a(_al_u817_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [28]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [28]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u819 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [25]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[27]),
    .o(_al_u819_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u820 (
    .a(_al_u819_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [27]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [27]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u821 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [24]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[26]),
    .o(_al_u821_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u822 (
    .a(_al_u821_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [26]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [26]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u823 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [23]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[25]),
    .o(_al_u823_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u824 (
    .a(_al_u823_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [25]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [25]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u825 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [22]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[24]),
    .o(_al_u825_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u826 (
    .a(_al_u825_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [24]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [24]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u827 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [21]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[23]),
    .o(_al_u827_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u828 (
    .a(_al_u827_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [23]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [23]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u829 (
    .a(\u_EXU_ALU/n0 [22]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[22]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u830 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[22]),
    .d(\u_EXU_LSU/n59 [20]),
    .e(o_ribm_addr[22]),
    .o(\u_EXU_LSU/n76 [22]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u831 (
    .a(\u_EXU_ALU/n0 [21]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[21]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u832 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[21]),
    .d(\u_EXU_LSU/n59 [19]),
    .e(o_ribm_addr[21]),
    .o(\u_EXU_LSU/n76 [21]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u833 (
    .a(\u_EXU_ALU/n0 [20]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[20]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u834 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[20]),
    .d(\u_EXU_LSU/n59 [18]),
    .e(o_ribm_addr[20]),
    .o(\u_EXU_LSU/n76 [20]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u835 (
    .a(\u_EXU_ALU/n0 [2]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[2]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u836 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[2]),
    .d(\u_EXU_LSU/n59 [0]),
    .e(o_ribm_addr[2]),
    .o(\u_EXU_LSU/n76 [2]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u837 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [17]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[19]),
    .o(_al_u837_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u838 (
    .a(_al_u837_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [19]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [19]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u839 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [16]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[18]),
    .o(_al_u839_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u840 (
    .a(_al_u839_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [18]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [18]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u841 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [15]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[17]),
    .o(_al_u841_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u842 (
    .a(_al_u841_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [17]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [17]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u843 (
    .a(\u_EXU_ALU/n0 [16]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[16]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u844 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[16]),
    .d(\u_EXU_LSU/n59 [14]),
    .e(o_ribm_addr[16]),
    .o(\u_EXU_LSU/n76 [16]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u845 (
    .a(\u_EXU_ALU/n0 [15]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[15]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u846 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[15]),
    .d(\u_EXU_LSU/n59 [13]),
    .e(o_ribm_addr[15]),
    .o(\u_EXU_LSU/n76 [15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u847 (
    .a(\u_EXU_ALU/n0 [14]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[14]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u848 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[14]),
    .d(\u_EXU_LSU/n59 [12]),
    .e(o_ribm_addr[14]),
    .o(\u_EXU_LSU/n76 [14]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u849 (
    .a(\u_EXU_ALU/n0 [13]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[13]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u850 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[13]),
    .d(\u_EXU_LSU/n59 [11]),
    .e(o_ribm_addr[13]),
    .o(\u_EXU_LSU/n76 [13]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~(B)*~((C*A))+D*B*~((C*A))+~(D)*B*(C*A)+D*B*(C*A))"),
    .INIT(16'h207f))
    _al_u851 (
    .a(i_ribm_gnt),
    .b(\u_EXU_LSU/n59 [10]),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_addr[12]),
    .o(_al_u851_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*C))*~(B)+~A*(D*C)*~(B)+~(~A)*(D*C)*B+~A*(D*C)*B)"),
    .INIT(16'hd111))
    _al_u852 (
    .a(_al_u851_o),
    .b(_al_u680_o),
    .c(\u_EXU_ALU/n0 [12]),
    .d(i_decinfo_grp[5]),
    .o(\u_EXU_LSU/n76 [12]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u853 (
    .a(\u_EXU_ALU/n0 [11]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[11]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u854 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[11]),
    .d(\u_EXU_LSU/n59 [9]),
    .e(o_ribm_addr[11]),
    .o(\u_EXU_LSU/n76 [11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u855 (
    .a(\u_EXU_ALU/n0 [10]),
    .b(i_decinfo_grp[5]),
    .o(alu2lsu_result[10]));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*~(C)*~(B)+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*~(B)+~((E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A))*C*B+(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)*C*B)"),
    .INIT(32'hf3d1e2c0))
    _al_u856 (
    .a(_al_u687_o),
    .b(_al_u680_o),
    .c(alu2lsu_result[10]),
    .d(\u_EXU_LSU/n59 [8]),
    .e(o_ribm_addr[10]),
    .o(\u_EXU_LSU/n76 [10]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u857 (
    .a(i_vld),
    .b(o_lsu_working),
    .c(i_decinfo_grp[1]),
    .d(i_rstn),
    .o(\u_EXU_LSU/mux10_b2_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u858 (
    .a(i_exu_op1[7]),
    .b(i_exu_op1[6]),
    .c(i_exu_op2[7]),
    .d(i_exu_op2[6]),
    .o(_al_u858_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u859 (
    .a(_al_u858_o),
    .b(i_exu_op1[5]),
    .c(i_exu_op1[4]),
    .d(i_exu_op2[5]),
    .e(i_exu_op2[4]),
    .o(_al_u859_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u860 (
    .a(i_exu_op1[22]),
    .b(i_exu_op1[20]),
    .c(i_exu_op2[22]),
    .d(i_exu_op2[20]),
    .o(_al_u860_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u861 (
    .a(i_exu_op1[17]),
    .b(i_exu_op2[17]),
    .o(\u_EXU_ALU/n168 [17]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u862 (
    .a(i_exu_op1[23]),
    .b(i_exu_op2[23]),
    .o(\u_EXU_ALU/n168 [23]));
  AL_MAP_LUT5 #(
    .EQN("(~C*~B*A*~(E@D))"),
    .INIT(32'h02000002))
    _al_u863 (
    .a(_al_u860_o),
    .b(\u_EXU_ALU/n168 [17]),
    .c(\u_EXU_ALU/n168 [23]),
    .d(i_exu_op1[21]),
    .e(i_exu_op2[21]),
    .o(_al_u863_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u864 (
    .a(i_exu_op1[1]),
    .b(i_exu_op1[0]),
    .c(i_exu_op2[1]),
    .d(i_exu_op2[0]),
    .o(_al_u864_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u865 (
    .a(i_exu_op1[3]),
    .b(i_exu_op1[2]),
    .c(i_exu_op2[3]),
    .d(i_exu_op2[2]),
    .o(_al_u865_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u866 (
    .a(_al_u859_o),
    .b(_al_u863_o),
    .c(_al_u864_o),
    .d(_al_u865_o),
    .o(_al_u866_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u867 (
    .a(i_exu_op1[26]),
    .b(i_exu_op1[24]),
    .c(i_exu_op2[26]),
    .d(i_exu_op2[24]),
    .o(_al_u867_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u868 (
    .a(i_exu_op1[31]),
    .b(i_exu_op2[31]),
    .o(\u_EXU_ALU/n168 [31]));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D@C))"),
    .INIT(16'h2002))
    _al_u869 (
    .a(_al_u867_o),
    .b(\u_EXU_ALU/n168 [31]),
    .c(i_exu_op1[28]),
    .d(i_exu_op2[28]),
    .o(_al_u869_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u870 (
    .a(i_exu_op1[14]),
    .b(i_exu_op1[13]),
    .c(i_exu_op2[14]),
    .d(i_exu_op2[13]),
    .o(_al_u870_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u871 (
    .a(i_exu_op1[10]),
    .b(i_exu_op1[8]),
    .c(i_exu_op2[10]),
    .d(i_exu_op2[8]),
    .o(_al_u871_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u872 (
    .a(_al_u869_o),
    .b(_al_u870_o),
    .c(_al_u871_o),
    .o(_al_u872_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u873 (
    .a(i_exu_op1[11]),
    .b(i_exu_op1[9]),
    .c(i_exu_op2[11]),
    .d(i_exu_op2[9]),
    .o(_al_u873_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u874 (
    .a(_al_u873_o),
    .b(i_exu_op1[15]),
    .c(i_exu_op1[12]),
    .d(i_exu_op2[15]),
    .e(i_exu_op2[12]),
    .o(_al_u874_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u875 (
    .a(i_exu_op1[27]),
    .b(i_exu_op1[25]),
    .c(i_exu_op2[27]),
    .d(i_exu_op2[25]),
    .o(_al_u875_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u876 (
    .a(i_exu_op1[29]),
    .b(i_exu_op2[29]),
    .o(\u_EXU_ALU/n168 [29]));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*A*~(E@D))"),
    .INIT(32'h08000008))
    _al_u877 (
    .a(_al_u874_o),
    .b(_al_u875_o),
    .c(\u_EXU_ALU/n168 [29]),
    .d(i_exu_op1[30]),
    .e(i_exu_op2[30]),
    .o(_al_u877_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u878 (
    .a(i_exu_op1[19]),
    .b(i_exu_op1[18]),
    .c(i_exu_op2[19]),
    .d(i_exu_op2[18]),
    .o(_al_u878_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u879 (
    .a(_al_u878_o),
    .b(i_exu_op1[16]),
    .c(i_exu_op2[16]),
    .o(_al_u879_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u880 (
    .a(_al_u866_o),
    .b(_al_u872_o),
    .c(_al_u877_o),
    .d(_al_u879_o),
    .e(i_decinfo[2]),
    .o(\u_EXU_BJU/bxx_beq ));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D*C*B*A))"),
    .INIT(32'h7fff0000))
    _al_u881 (
    .a(_al_u866_o),
    .b(_al_u872_o),
    .c(_al_u877_o),
    .d(_al_u879_o),
    .e(i_decinfo[3]),
    .o(\u_EXU_BJU/bxx_bne ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u882 (
    .a(\u_EXU_ALU/n253 ),
    .b(i_decinfo[5]),
    .c(i_decinfo[4]),
    .o(_al_u882_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h0145))
    _al_u883 (
    .a(_al_u882_o),
    .b(\u_EXU_ALU/n261 ),
    .c(i_decinfo[7]),
    .d(i_decinfo[6]),
    .o(_al_u883_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D@(C*~B*~A)))"),
    .INIT(32'h10ef0000))
    _al_u884 (
    .a(\u_EXU_BJU/bxx_beq ),
    .b(\u_EXU_BJU/bxx_bne ),
    .c(_al_u883_o),
    .d(i_decinfo[8]),
    .e(i_decinfo_grp[2]),
    .o(o_exu_taken));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u885 (
    .a(i_ribm_rsp),
    .b(\u_EXU_LSU/access2_once ),
    .c(\u_EXU_LSU/handshake_rdy_last ),
    .o(_al_u885_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~B*~(~E*D*A))"),
    .INIT(32'h03030103))
    _al_u886 (
    .a(i_vld),
    .b(_al_u422_o),
    .c(_al_u885_o),
    .d(i_decinfo_grp[1]),
    .e(\u_EXU_LSU/working ),
    .o(\u_EXU_LSU/n30 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u887 (
    .a(i_ribm_rsp),
    .b(\u_EXU_LSU/handshake_rdy_last ),
    .c(i_rstn),
    .o(_al_u887_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*~(~E*D*A))"),
    .INIT(32'h30301030))
    _al_u888 (
    .a(i_vld),
    .b(_al_u422_o),
    .c(_al_u887_o),
    .d(i_decinfo_grp[1]),
    .e(\u_EXU_LSU/working ),
    .o(\u_EXU_LSU/mux11_b0_sel_is_2_o ));
  AL_MAP_LUT4 #(
    .EQN("~(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hfdec))
    _al_u889 (
    .a(i_ribm_gnt),
    .b(_al_u680_o),
    .c(\u_EXU_LSU/n57 ),
    .d(o_ribm_req),
    .o(\u_EXU_LSU/n75 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u890 (
    .a(i_ribm_rsp),
    .b(o_exu_rdwen0),
    .c(\u_EXU_LSU/handshake_rdy_last ),
    .o(_al_u890_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u891 (
    .a(o_rdidx0[4]),
    .b(o_rdidx0[3]),
    .c(o_rdidx2[3]),
    .d(o_rdidx2[4]),
    .o(_al_u891_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C@B)*~(D@A))"),
    .INIT(16'h8241))
    _al_u892 (
    .a(o_rdidx0[1]),
    .b(o_rdidx0[0]),
    .c(o_rdidx2[0]),
    .d(o_rdidx2[1]),
    .o(_al_u892_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u893 (
    .a(_al_u891_o),
    .b(_al_u892_o),
    .c(o_rdidx0[2]),
    .d(o_rdidx2[2]),
    .o(n7_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(D*~A*~(C*B))"),
    .INIT(16'h1500))
    _al_u894 (
    .a(_al_u422_o),
    .b(_al_u890_o),
    .c(n7_lutinv),
    .d(o_exu_rdwen2),
    .o(\u_EXU_LSU/n18_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u895 (
    .a(i_decinfo[1]),
    .b(o_exu_rdwen0),
    .o(\u_EXU_LSU/n8 ));
  AL_MAP_LUT5 #(
    .EQN("(B*~(D)*~((E*~C*A))+B*D*~((E*~C*A))+~(B)*D*(E*~C*A)+B*D*(E*~C*A))"),
    .INIT(32'hcec4cccc))
    _al_u896 (
    .a(i_vld),
    .b(\u_EXU_LSU/n18_lutinv ),
    .c(o_lsu_working),
    .d(\u_EXU_LSU/n8 ),
    .e(i_decinfo_grp[1]),
    .o(\u_EXU_LSU/n23 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u897 (
    .a(i_exu_op1[15]),
    .b(i_exu_op1[14]),
    .c(i_exu_op2[0]),
    .o(_al_u897_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*~(D)+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(D)+~(~A)*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D)"),
    .INIT(32'h0faa33aa))
    _al_u898 (
    .a(_al_u897_o),
    .b(i_exu_op1[13]),
    .c(i_exu_op1[12]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u898_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u899 (
    .a(i_exu_op1[9]),
    .b(i_exu_op1[8]),
    .c(i_exu_op2[0]),
    .o(_al_u899_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u900 (
    .a(i_exu_op1[11]),
    .b(i_exu_op1[10]),
    .c(i_exu_op2[0]),
    .o(_al_u900_o));
  AL_MAP_LUT5 #(
    .EQN("~(A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'h33550f55))
    _al_u901 (
    .a(_al_u898_o),
    .b(_al_u899_o),
    .c(_al_u900_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(\u_EXU_ALU/n369_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u902 (
    .a(i_exu_op1[1]),
    .b(i_exu_op1[0]),
    .c(i_exu_op2[0]),
    .o(_al_u902_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u903 (
    .a(i_exu_op1[3]),
    .b(i_exu_op1[2]),
    .c(i_exu_op2[0]),
    .o(_al_u903_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u904 (
    .a(_al_u902_o),
    .b(_al_u903_o),
    .c(i_exu_op2[1]),
    .o(_al_u904_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u905 (
    .a(i_exu_op1[5]),
    .b(i_exu_op1[4]),
    .c(i_exu_op2[0]),
    .o(_al_u905_o));
  AL_MAP_LUT5 #(
    .EQN("(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'haa0faa33))
    _al_u906 (
    .a(_al_u905_o),
    .b(i_exu_op1[7]),
    .c(i_exu_op1[6]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u906_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*~(D)+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(D)+~(~A)*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D+~A*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*D)"),
    .INIT(32'hcc55f055))
    _al_u907 (
    .a(\u_EXU_ALU/n369_lutinv ),
    .b(_al_u904_o),
    .c(_al_u906_o),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(_al_u907_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u908 (
    .a(i_exu_op2[13]),
    .b(i_exu_op2[12]),
    .o(_al_u908_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u909 (
    .a(i_exu_op2[6]),
    .b(i_exu_op2[5]),
    .o(_al_u909_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u910 (
    .a(_al_u909_o),
    .b(i_exu_op2[10]),
    .c(i_exu_op2[9]),
    .d(i_exu_op2[8]),
    .e(i_exu_op2[7]),
    .o(_al_u910_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*~B*A)"),
    .INIT(32'h00000200))
    _al_u911 (
    .a(_al_u908_o),
    .b(i_exu_op2[15]),
    .c(i_exu_op2[14]),
    .d(_al_u910_o),
    .e(i_exu_op2[11]),
    .o(_al_u911_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u912 (
    .a(i_exu_op2[30]),
    .b(i_exu_op2[29]),
    .c(i_exu_op2[22]),
    .d(i_exu_op2[21]),
    .o(_al_u912_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u913 (
    .a(i_exu_op2[31]),
    .b(i_exu_op2[28]),
    .o(_al_u913_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u914 (
    .a(i_exu_op2[27]),
    .b(i_exu_op2[26]),
    .c(i_exu_op2[25]),
    .o(_al_u914_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u915 (
    .a(_al_u912_o),
    .b(_al_u913_o),
    .c(i_exu_op2[24]),
    .d(_al_u914_o),
    .o(_al_u915_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u916 (
    .a(i_exu_op2[17]),
    .b(i_exu_op2[16]),
    .o(_al_u916_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u917 (
    .a(_al_u916_o),
    .b(i_exu_op2[23]),
    .c(i_exu_op2[20]),
    .d(i_exu_op2[19]),
    .e(i_exu_op2[18]),
    .o(_al_u917_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u918 (
    .a(_al_u911_o),
    .b(_al_u915_o),
    .c(_al_u917_o),
    .d(i_decinfo[2]),
    .o(_al_u918_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u919 (
    .a(i_exu_op1[25]),
    .b(i_exu_op1[24]),
    .c(i_exu_op2[0]),
    .o(_al_u919_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u920 (
    .a(i_exu_op1[27]),
    .b(i_exu_op1[26]),
    .c(i_exu_op2[0]),
    .o(_al_u920_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u921 (
    .a(_al_u919_o),
    .b(_al_u920_o),
    .c(i_exu_op2[1]),
    .o(_al_u921_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcaf0))
    _al_u922 (
    .a(i_exu_op1[29]),
    .b(i_exu_op1[28]),
    .c(i_exu_op2[0]),
    .d(i_exu_op2[1]),
    .o(_al_u922_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u923 (
    .a(i_exu_op1[31]),
    .b(i_exu_op1[30]),
    .c(_al_u922_o),
    .d(i_exu_op2[1]),
    .o(_al_u923_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u924 (
    .a(i_exu_op2[4]),
    .b(i_exu_op2[3]),
    .o(_al_u924_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u925 (
    .a(_al_u921_o),
    .b(_al_u923_o),
    .c(_al_u924_o),
    .d(i_exu_op2[2]),
    .o(_al_u925_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u926 (
    .a(i_exu_op1[17]),
    .b(i_exu_op1[16]),
    .c(i_exu_op2[0]),
    .o(_al_u926_o));
  AL_MAP_LUT5 #(
    .EQN("(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'haa0faa33))
    _al_u927 (
    .a(_al_u926_o),
    .b(i_exu_op1[19]),
    .c(i_exu_op1[18]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u927_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u928 (
    .a(i_exu_op1[23]),
    .b(i_exu_op1[22]),
    .c(i_exu_op2[0]),
    .o(_al_u928_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*~(D)+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(D)+~(~A)*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D)"),
    .INIT(32'h0faa33aa))
    _al_u929 (
    .a(_al_u928_o),
    .b(i_exu_op1[21]),
    .c(i_exu_op1[20]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u929_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u930 (
    .a(i_exu_op2[4]),
    .b(i_exu_op2[3]),
    .o(_al_u930_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u931 (
    .a(_al_u927_o),
    .b(_al_u929_o),
    .c(_al_u930_o),
    .d(i_exu_op2[2]),
    .o(_al_u931_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~D*~C*~(E*~A)))"),
    .INIT(32'hccc4ccc0))
    _al_u932 (
    .a(_al_u907_o),
    .b(_al_u918_o),
    .c(_al_u925_o),
    .d(_al_u931_o),
    .e(i_exu_op2[4]),
    .o(\u_EXU_ALU/alu_sll [31]));
  AL_MAP_LUT5 #(
    .EQN("(E*~(C*B)*~(D*A))"),
    .INIT(32'h153f0000))
    _al_u933 (
    .a(\u_EXU_ALU/n0 [31]),
    .b(\u_EXU_ALU/n33 [31]),
    .c(i_decinfo[1]),
    .d(i_decinfo_grp[5]),
    .e(i_decinfo_grp[0]),
    .o(_al_u933_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D)"),
    .INIT(16'h155f))
    _al_u934 (
    .a(i_decinfo[7]),
    .b(i_decinfo[6]),
    .c(i_exu_op1[31]),
    .d(i_exu_op2[31]),
    .o(_al_u934_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u935 (
    .a(_al_u933_o),
    .b(_al_u934_o),
    .c(\u_EXU_ALU/n168 [31]),
    .d(i_decinfo[5]),
    .o(_al_u935_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u936 (
    .a(i_exu_op2[15]),
    .b(i_exu_op2[12]),
    .o(_al_u936_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u937 (
    .a(_al_u936_o),
    .b(i_exu_op2[11]),
    .c(i_exu_op2[10]),
    .d(i_exu_op2[9]),
    .e(i_exu_op2[8]),
    .o(_al_u937_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u938 (
    .a(i_exu_op2[14]),
    .b(i_exu_op2[13]),
    .c(i_exu_op2[7]),
    .d(i_exu_op2[6]),
    .e(i_exu_op2[5]),
    .o(_al_u938_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u939 (
    .a(_al_u937_o),
    .b(_al_u938_o),
    .o(_al_u939_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u940 (
    .a(i_exu_op2[19]),
    .b(i_exu_op2[18]),
    .c(i_exu_op2[17]),
    .d(i_exu_op2[16]),
    .o(_al_u940_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u941 (
    .a(i_exu_op2[23]),
    .b(i_exu_op2[22]),
    .o(_al_u941_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u942 (
    .a(i_exu_op2[21]),
    .b(i_exu_op2[20]),
    .o(_al_u942_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u943 (
    .a(_al_u940_o),
    .b(_al_u941_o),
    .c(_al_u942_o),
    .o(_al_u943_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u944 (
    .a(i_exu_op2[29]),
    .b(i_exu_op2[28]),
    .o(_al_u944_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u945 (
    .a(_al_u944_o),
    .b(i_exu_op2[31]),
    .c(i_exu_op2[30]),
    .o(_al_u945_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u946 (
    .a(i_exu_op2[27]),
    .b(i_exu_op2[26]),
    .c(i_exu_op2[25]),
    .d(i_exu_op2[24]),
    .o(_al_u946_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u947 (
    .a(_al_u939_o),
    .b(_al_u943_o),
    .c(_al_u945_o),
    .d(_al_u946_o),
    .o(\u_EXU_ALU/n179_neg_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u948 (
    .a(i_exu_op2[2]),
    .b(i_exu_op2[1]),
    .o(_al_u948_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*B*A))"),
    .INIT(16'hf070))
    _al_u949 (
    .a(_al_u924_o),
    .b(_al_u948_o),
    .c(i_exu_op1[31]),
    .d(i_exu_op2[0]),
    .o(\u_EXU_ALU/n237_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*C*B))"),
    .INIT(16'h2aaa))
    _al_u950 (
    .a(_al_u935_o),
    .b(\u_EXU_ALU/n179_neg_lutinv ),
    .c(\u_EXU_ALU/n237_lutinv ),
    .d(i_decinfo[4]),
    .o(_al_u950_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u951 (
    .a(_al_u913_o),
    .b(i_exu_op2[27]),
    .c(i_exu_op2[26]),
    .d(i_exu_op2[25]),
    .e(i_exu_op2[24]),
    .o(_al_u951_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    _al_u952 (
    .a(_al_u911_o),
    .b(_al_u917_o),
    .c(_al_u951_o),
    .d(_al_u912_o),
    .e(i_exu_op2[4]),
    .o(\u_EXU_ALU/u1029_sel_is_0_o ));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u953 (
    .a(i_exu_op1[31]),
    .b(i_exu_op2[2]),
    .c(i_exu_op2[1]),
    .d(i_exu_op2[0]),
    .o(\u_EXU_ALU/n77_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(~B*~A))"),
    .INIT(8'h0e))
    _al_u954 (
    .a(i_decinfo[4]),
    .b(i_decinfo[3]),
    .c(i_exu_op2[3]),
    .o(_al_u954_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u955 (
    .a(\u_EXU_ALU/u1029_sel_is_0_o ),
    .b(\u_EXU_ALU/n77_lutinv ),
    .c(_al_u954_o),
    .o(_al_u955_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B))"),
    .INIT(32'h00004777))
    _al_u956 (
    .a(bju_rdwdata[31]),
    .b(bju_rdwen),
    .c(i_csr_rdata[31]),
    .d(i_decinfo_grp[4]),
    .e(i_decinfo_grp[0]),
    .o(_al_u956_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*B*~A))"),
    .INIT(16'h00fb))
    _al_u957 (
    .a(\u_EXU_ALU/alu_sll [31]),
    .b(_al_u950_o),
    .c(_al_u955_o),
    .d(_al_u956_o),
    .o(o_rdwdata0[31]));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u958 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[30]),
    .d(i_exu_op2[30]),
    .o(_al_u958_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u959 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[30]),
    .c(i_exu_op2[30]),
    .o(\u_EXU_ALU/alu_and [30]));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*~A*~(E*B))"),
    .INIT(32'h00010005))
    _al_u960 (
    .a(alu2lsu_result[30]),
    .b(\u_EXU_ALU/n33 [30]),
    .c(_al_u958_o),
    .d(\u_EXU_ALU/alu_and [30]),
    .e(i_decinfo[1]),
    .o(_al_u960_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u961 (
    .a(_al_u946_o),
    .b(_al_u944_o),
    .c(i_decinfo[4]),
    .d(i_exu_op2[31]),
    .e(i_exu_op2[30]),
    .o(_al_u961_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B*A))"),
    .INIT(8'h70))
    _al_u962 (
    .a(_al_u924_o),
    .b(_al_u948_o),
    .c(i_exu_op1[31]),
    .o(\u_EXU_ALU/n236_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u963 (
    .a(_al_u943_o),
    .b(_al_u961_o),
    .c(\u_EXU_ALU/n236_lutinv ),
    .d(_al_u937_o),
    .e(_al_u938_o),
    .o(_al_u963_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u964 (
    .a(i_exu_op1[31]),
    .b(i_exu_op1[30]),
    .c(i_exu_op2[1]),
    .d(i_exu_op2[0]),
    .o(\u_EXU_ALU/n111_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u965 (
    .a(i_exu_op2[3]),
    .b(i_exu_op2[2]),
    .o(_al_u965_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u966 (
    .a(\u_EXU_ALU/n111_lutinv ),
    .b(_al_u965_o),
    .o(\u_EXU_ALU/n45_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u967 (
    .a(\u_EXU_ALU/n45_lutinv ),
    .b(i_exu_op2[4]),
    .c(_al_u911_o),
    .d(_al_u916_o),
    .o(_al_u967_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u968 (
    .a(_al_u911_o),
    .b(_al_u917_o),
    .c(_al_u951_o),
    .d(_al_u912_o),
    .o(\u_EXU_ALU/n281_neg_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*~(E*~D*C))"),
    .INIT(32'h22022222))
    _al_u969 (
    .a(_al_u960_o),
    .b(_al_u963_o),
    .c(_al_u967_o),
    .d(\u_EXU_LSU/mux14_b1_sel_is_0_o ),
    .e(\u_EXU_ALU/n281_neg_lutinv ),
    .o(_al_u969_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff330f55))
    _al_u970 (
    .a(i_exu_op1[2]),
    .b(i_exu_op1[1]),
    .c(i_exu_op1[0]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u970_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u971 (
    .a(i_exu_op1[4]),
    .b(i_exu_op1[3]),
    .c(i_exu_op2[0]),
    .o(_al_u971_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u972 (
    .a(i_exu_op1[6]),
    .b(i_exu_op1[5]),
    .c(i_exu_op2[0]),
    .o(_al_u972_o));
  AL_MAP_LUT5 #(
    .EQN("((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'haaccaaf0))
    _al_u973 (
    .a(_al_u970_o),
    .b(_al_u971_o),
    .c(_al_u972_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u973_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u974 (
    .a(i_exu_op1[10]),
    .b(i_exu_op1[9]),
    .c(i_exu_op2[0]),
    .o(_al_u974_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*~(D)+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(D)+~(~A)*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D)"),
    .INIT(32'h0faa33aa))
    _al_u975 (
    .a(_al_u974_o),
    .b(i_exu_op1[8]),
    .c(i_exu_op1[7]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u975_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u976 (
    .a(i_exu_op1[12]),
    .b(i_exu_op1[11]),
    .c(i_exu_op2[0]),
    .o(_al_u976_o));
  AL_MAP_LUT5 #(
    .EQN("(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~(~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+~(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'haa0faa33))
    _al_u977 (
    .a(_al_u976_o),
    .b(i_exu_op1[14]),
    .c(i_exu_op1[13]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u977_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'h5533550f))
    _al_u978 (
    .a(_al_u973_o),
    .b(_al_u975_o),
    .c(_al_u977_o),
    .d(i_exu_op2[3]),
    .e(i_exu_op2[2]),
    .o(\u_EXU_ALU/n402_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u979 (
    .a(i_exu_op1[20]),
    .b(i_exu_op1[19]),
    .c(i_exu_op2[0]),
    .o(_al_u979_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u980 (
    .a(i_exu_op1[22]),
    .b(i_exu_op1[21]),
    .c(i_exu_op2[0]),
    .o(_al_u980_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u981 (
    .a(_al_u979_o),
    .b(_al_u980_o),
    .c(i_exu_op2[1]),
    .o(_al_u981_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u982 (
    .a(i_exu_op1[18]),
    .b(i_exu_op1[17]),
    .c(i_exu_op2[0]),
    .o(_al_u982_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*~(D)+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(D)+~(~A)*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D)"),
    .INIT(32'h0faa33aa))
    _al_u983 (
    .a(_al_u982_o),
    .b(i_exu_op1[16]),
    .c(i_exu_op1[15]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u983_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u984 (
    .a(_al_u981_o),
    .b(_al_u983_o),
    .c(i_exu_op2[2]),
    .o(\u_EXU_ALU/n362_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u985 (
    .a(i_exu_op1[26]),
    .b(i_exu_op1[25]),
    .c(i_exu_op2[0]),
    .o(_al_u985_o));
  AL_MAP_LUT5 #(
    .EQN("~(~A*~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*~(D)+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(D)+~(~A)*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D+~A*(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*D)"),
    .INIT(32'h0faa33aa))
    _al_u986 (
    .a(_al_u985_o),
    .b(i_exu_op1[24]),
    .c(i_exu_op1[23]),
    .d(i_exu_op2[1]),
    .e(i_exu_op2[0]),
    .o(_al_u986_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u987 (
    .a(i_exu_op1[30]),
    .b(i_exu_op1[29]),
    .c(i_exu_op2[0]),
    .o(_al_u987_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u988 (
    .a(i_exu_op1[28]),
    .b(i_exu_op1[27]),
    .c(i_exu_op2[0]),
    .o(_al_u988_o));
  AL_MAP_LUT5 #(
    .EQN("((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*~(A)*~(D)+(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*~(D)+~((B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E))*A*D+(B*~(C)*~(E)+B*C*~(E)+~(B)*C*E+B*C*E)*A*D)"),
    .INIT(32'haaf0aacc))
    _al_u989 (
    .a(_al_u986_o),
    .b(_al_u987_o),
    .c(_al_u988_o),
    .d(i_exu_op2[2]),
    .e(i_exu_op2[1]),
    .o(_al_u989_o));
  AL_MAP_LUT5 #(
    .EQN("~((~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E)*~(A)*~(D)+(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E)*A*~(D)+~((~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E))*A*D+(~C*~(B)*~(E)+~C*B*~(E)+~(~C)*B*E+~C*B*E)*A*D)"),
    .INIT(32'h553355f0))
    _al_u990 (
    .a(\u_EXU_ALU/n402_lutinv ),
    .b(\u_EXU_ALU/n362_lutinv ),
    .c(_al_u989_o),
    .d(i_exu_op2[4]),
    .e(i_exu_op2[3]),
    .o(_al_u990_o));
  AL_MAP_LUT4 #(
    .EQN("~((D*C)*~(A)*~(B)+(D*C)*A*~(B)+~((D*C))*A*B+(D*C)*A*B)"),
    .INIT(16'h4777))
    _al_u991 (
    .a(bju_rdwdata[30]),
    .b(bju_rdwen),
    .c(i_csr_rdata[30]),
    .d(i_decinfo_grp[4]),
    .o(_al_u991_o));
  AL_MAP_LUT5 #(
    .EQN("~(C*~((A*~(E*~B)))*~(D)+C*(A*~(E*~B))*~(D)+~(C)*(A*~(E*~B))*D+C*(A*~(E*~B))*D)"),
    .INIT(32'h770f550f))
    _al_u992 (
    .a(_al_u969_o),
    .b(_al_u990_o),
    .c(_al_u991_o),
    .d(i_decinfo_grp[0]),
    .e(_al_u918_o),
    .o(o_rdwdata0[30]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u993 (
    .a(i_decinfo[6]),
    .b(i_exu_op1[29]),
    .c(i_exu_op2[29]),
    .o(\u_EXU_ALU/alu_and [29]));
  AL_MAP_LUT4 #(
    .EQN("(D*~B*~(C*A))"),
    .INIT(16'h1300))
    _al_u994 (
    .a(\u_EXU_ALU/n33 [29]),
    .b(\u_EXU_ALU/alu_and [29]),
    .c(i_decinfo[1]),
    .d(i_decinfo_grp[0]),
    .o(_al_u994_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'haee0))
    _al_u995 (
    .a(i_decinfo[7]),
    .b(i_decinfo[5]),
    .c(i_exu_op1[29]),
    .d(i_exu_op2[29]),
    .o(_al_u995_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u996 (
    .a(_al_u994_o),
    .b(\u_EXU_ALU/n0 [29]),
    .c(_al_u995_o),
    .d(i_decinfo_grp[5]),
    .o(_al_u996_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u997 (
    .a(i_exu_op2[27]),
    .b(i_exu_op2[26]),
    .c(i_exu_op2[25]),
    .d(i_exu_op2[24]),
    .o(_al_u997_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u998 (
    .a(_al_u997_o),
    .b(_al_u912_o),
    .c(_al_u913_o),
    .d(i_exu_op2[4]),
    .o(_al_u998_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u999 (
    .a(i_exu_op1[30]),
    .b(i_exu_op1[29]),
    .c(i_exu_op2[0]),
    .o(_al_u999_o));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/add0/ucin_al_u1469"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/add0/u11_al_u1472  (
    .a({i_exu_op1[13],i_exu_op1[11]}),
    .b({i_exu_op1[14],i_exu_op1[12]}),
    .c(2'b00),
    .d({i_exu_op2[13],i_exu_op2[11]}),
    .e({i_exu_op2[14],i_exu_op2[12]}),
    .fci(\u_EXU_ALU/add0/c11 ),
    .f({\u_EXU_ALU/n0 [13],\u_EXU_ALU/n0 [11]}),
    .fco(\u_EXU_ALU/add0/c15 ),
    .fx({\u_EXU_ALU/n0 [14],\u_EXU_ALU/n0 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/add0/ucin_al_u1469"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/add0/u15_al_u1473  (
    .a({i_exu_op1[17],i_exu_op1[15]}),
    .b({i_exu_op1[18],i_exu_op1[16]}),
    .c(2'b00),
    .d({i_exu_op2[17],i_exu_op2[15]}),
    .e({i_exu_op2[18],i_exu_op2[16]}),
    .fci(\u_EXU_ALU/add0/c15 ),
    .f({\u_EXU_ALU/n0 [17],\u_EXU_ALU/n0 [15]}),
    .fco(\u_EXU_ALU/add0/c19 ),
    .fx({\u_EXU_ALU/n0 [18],\u_EXU_ALU/n0 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/add0/ucin_al_u1469"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/add0/u19_al_u1474  (
    .a({i_exu_op1[21],i_exu_op1[19]}),
    .b({i_exu_op1[22],i_exu_op1[20]}),
    .c(2'b00),
    .d({i_exu_op2[21],i_exu_op2[19]}),
    .e({i_exu_op2[22],i_exu_op2[20]}),
    .fci(\u_EXU_ALU/add0/c19 ),
    .f({\u_EXU_ALU/n0 [21],\u_EXU_ALU/n0 [19]}),
    .fco(\u_EXU_ALU/add0/c23 ),
    .fx({\u_EXU_ALU/n0 [22],\u_EXU_ALU/n0 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/add0/ucin_al_u1469"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/add0/u23_al_u1475  (
    .a({i_exu_op1[25],i_exu_op1[23]}),
    .b({i_exu_op1[26],i_exu_op1[24]}),
    .c(2'b00),
    .d({i_exu_op2[25],i_exu_op2[23]}),
    .e({i_exu_op2[26],i_exu_op2[24]}),
    .fci(\u_EXU_ALU/add0/c23 ),
    .f({\u_EXU_ALU/n0 [25],\u_EXU_ALU/n0 [23]}),
    .fco(\u_EXU_ALU/add0/c27 ),
    .fx({\u_EXU_ALU/n0 [26],\u_EXU_ALU/n0 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/add0/ucin_al_u1469"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/add0/u27_al_u1476  (
    .a({i_exu_op1[29],i_exu_op1[27]}),
    .b({i_exu_op1[30],i_exu_op1[28]}),
    .c(2'b00),
    .d({i_exu_op2[29],i_exu_op2[27]}),
    .e({i_exu_op2[30],i_exu_op2[28]}),
    .fci(\u_EXU_ALU/add0/c27 ),
    .f({\u_EXU_ALU/n0 [29],\u_EXU_ALU/n0 [27]}),
    .fco(\u_EXU_ALU/add0/c31 ),
    .fx({\u_EXU_ALU/n0 [30],\u_EXU_ALU/n0 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/add0/ucin_al_u1469"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/add0/u31_al_u1477  (
    .a({open_n90,i_exu_op1[31]}),
    .c(2'b00),
    .d({open_n95,i_exu_op2[31]}),
    .fci(\u_EXU_ALU/add0/c31 ),
    .f({open_n112,\u_EXU_ALU/n0 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/add0/ucin_al_u1469"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/add0/u3_al_u1470  (
    .a({i_exu_op1[5],i_exu_op1[3]}),
    .b({i_exu_op1[6],i_exu_op1[4]}),
    .c(2'b00),
    .d({i_exu_op2[5],i_exu_op2[3]}),
    .e({i_exu_op2[6],i_exu_op2[4]}),
    .fci(\u_EXU_ALU/add0/c3 ),
    .f({\u_EXU_ALU/n0 [5],\u_EXU_ALU/n0 [3]}),
    .fco(\u_EXU_ALU/add0/c7 ),
    .fx({\u_EXU_ALU/n0 [6],\u_EXU_ALU/n0 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/add0/ucin_al_u1469"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/add0/u7_al_u1471  (
    .a({i_exu_op1[9],i_exu_op1[7]}),
    .b({i_exu_op1[10],i_exu_op1[8]}),
    .c(2'b00),
    .d({i_exu_op2[9],i_exu_op2[7]}),
    .e({i_exu_op2[10],i_exu_op2[8]}),
    .fci(\u_EXU_ALU/add0/c7 ),
    .f({\u_EXU_ALU/n0 [9],\u_EXU_ALU/n0 [7]}),
    .fco(\u_EXU_ALU/add0/c11 ),
    .fx({\u_EXU_ALU/n0 [10],\u_EXU_ALU/n0 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/add0/ucin_al_u1469"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/add0/ucin_al_u1469  (
    .a({i_exu_op1[1],1'b0}),
    .b({i_exu_op1[2],i_exu_op1[0]}),
    .c(2'b00),
    .d({i_exu_op2[1],1'b1}),
    .e({i_exu_op2[2],i_exu_op2[0]}),
    .f({\u_EXU_ALU/n0 [1],open_n171}),
    .fco(\u_EXU_ALU/add0/c3 ),
    .fx({\u_EXU_ALU/n0 [2],\u_EXU_ALU/n0 [0]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin  (
    .a({i_exu_op1[0],1'b0}),
    .b({i_exu_op2[0],open_n174}),
    .fco(\u_EXU_ALU/lt0_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_10|u_EXU_ALU/lt0_9  (
    .a(i_exu_op1[10:9]),
    .b(i_exu_op2[10:9]),
    .fci(\u_EXU_ALU/lt0_c9 ),
    .fco(\u_EXU_ALU/lt0_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_12|u_EXU_ALU/lt0_11  (
    .a(i_exu_op1[12:11]),
    .b(i_exu_op2[12:11]),
    .fci(\u_EXU_ALU/lt0_c11 ),
    .fco(\u_EXU_ALU/lt0_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_14|u_EXU_ALU/lt0_13  (
    .a(i_exu_op1[14:13]),
    .b(i_exu_op2[14:13]),
    .fci(\u_EXU_ALU/lt0_c13 ),
    .fco(\u_EXU_ALU/lt0_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_16|u_EXU_ALU/lt0_15  (
    .a(i_exu_op1[16:15]),
    .b(i_exu_op2[16:15]),
    .fci(\u_EXU_ALU/lt0_c15 ),
    .fco(\u_EXU_ALU/lt0_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_18|u_EXU_ALU/lt0_17  (
    .a(i_exu_op1[18:17]),
    .b(i_exu_op2[18:17]),
    .fci(\u_EXU_ALU/lt0_c17 ),
    .fco(\u_EXU_ALU/lt0_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_20|u_EXU_ALU/lt0_19  (
    .a(i_exu_op1[20:19]),
    .b(i_exu_op2[20:19]),
    .fci(\u_EXU_ALU/lt0_c19 ),
    .fco(\u_EXU_ALU/lt0_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_22|u_EXU_ALU/lt0_21  (
    .a(i_exu_op1[22:21]),
    .b(i_exu_op2[22:21]),
    .fci(\u_EXU_ALU/lt0_c21 ),
    .fco(\u_EXU_ALU/lt0_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_24|u_EXU_ALU/lt0_23  (
    .a(i_exu_op1[24:23]),
    .b(i_exu_op2[24:23]),
    .fci(\u_EXU_ALU/lt0_c23 ),
    .fco(\u_EXU_ALU/lt0_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_26|u_EXU_ALU/lt0_25  (
    .a(i_exu_op1[26:25]),
    .b(i_exu_op2[26:25]),
    .fci(\u_EXU_ALU/lt0_c25 ),
    .fco(\u_EXU_ALU/lt0_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_28|u_EXU_ALU/lt0_27  (
    .a(i_exu_op1[28:27]),
    .b(i_exu_op2[28:27]),
    .fci(\u_EXU_ALU/lt0_c27 ),
    .fco(\u_EXU_ALU/lt0_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_2|u_EXU_ALU/lt0_1  (
    .a(i_exu_op1[2:1]),
    .b(i_exu_op2[2:1]),
    .fci(\u_EXU_ALU/lt0_c1 ),
    .fco(\u_EXU_ALU/lt0_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_30|u_EXU_ALU/lt0_29  (
    .a(i_exu_op1[30:29]),
    .b(i_exu_op2[30:29]),
    .fci(\u_EXU_ALU/lt0_c29 ),
    .fco(\u_EXU_ALU/lt0_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_4|u_EXU_ALU/lt0_3  (
    .a(i_exu_op1[4:3]),
    .b(i_exu_op2[4:3]),
    .fci(\u_EXU_ALU/lt0_c3 ),
    .fco(\u_EXU_ALU/lt0_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_6|u_EXU_ALU/lt0_5  (
    .a(i_exu_op1[6:5]),
    .b(i_exu_op2[6:5]),
    .fci(\u_EXU_ALU/lt0_c5 ),
    .fco(\u_EXU_ALU/lt0_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_8|u_EXU_ALU/lt0_7  (
    .a(i_exu_op1[8:7]),
    .b(i_exu_op2[8:7]),
    .fci(\u_EXU_ALU/lt0_c7 ),
    .fco(\u_EXU_ALU/lt0_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt0_0|u_EXU_ALU/lt0_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt0_cout|u_EXU_ALU/lt0_31  (
    .a({1'b0,i_exu_op2[31]}),
    .b({1'b1,i_exu_op1[31]}),
    .fci(\u_EXU_ALU/lt0_c31 ),
    .f({\u_EXU_ALU/n253 ,open_n578}));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin  (
    .a({i_exu_op1[0],1'b0}),
    .b({i_exu_op2[0],open_n584}),
    .fco(\u_EXU_ALU/lt1_c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_10|u_EXU_ALU/lt1_9  (
    .a(i_exu_op1[10:9]),
    .b(i_exu_op2[10:9]),
    .fci(\u_EXU_ALU/lt1_c9 ),
    .fco(\u_EXU_ALU/lt1_c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_12|u_EXU_ALU/lt1_11  (
    .a(i_exu_op1[12:11]),
    .b(i_exu_op2[12:11]),
    .fci(\u_EXU_ALU/lt1_c11 ),
    .fco(\u_EXU_ALU/lt1_c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_14|u_EXU_ALU/lt1_13  (
    .a(i_exu_op1[14:13]),
    .b(i_exu_op2[14:13]),
    .fci(\u_EXU_ALU/lt1_c13 ),
    .fco(\u_EXU_ALU/lt1_c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_16|u_EXU_ALU/lt1_15  (
    .a(i_exu_op1[16:15]),
    .b(i_exu_op2[16:15]),
    .fci(\u_EXU_ALU/lt1_c15 ),
    .fco(\u_EXU_ALU/lt1_c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_18|u_EXU_ALU/lt1_17  (
    .a(i_exu_op1[18:17]),
    .b(i_exu_op2[18:17]),
    .fci(\u_EXU_ALU/lt1_c17 ),
    .fco(\u_EXU_ALU/lt1_c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_20|u_EXU_ALU/lt1_19  (
    .a(i_exu_op1[20:19]),
    .b(i_exu_op2[20:19]),
    .fci(\u_EXU_ALU/lt1_c19 ),
    .fco(\u_EXU_ALU/lt1_c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_22|u_EXU_ALU/lt1_21  (
    .a(i_exu_op1[22:21]),
    .b(i_exu_op2[22:21]),
    .fci(\u_EXU_ALU/lt1_c21 ),
    .fco(\u_EXU_ALU/lt1_c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_24|u_EXU_ALU/lt1_23  (
    .a(i_exu_op1[24:23]),
    .b(i_exu_op2[24:23]),
    .fci(\u_EXU_ALU/lt1_c23 ),
    .fco(\u_EXU_ALU/lt1_c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_26|u_EXU_ALU/lt1_25  (
    .a(i_exu_op1[26:25]),
    .b(i_exu_op2[26:25]),
    .fci(\u_EXU_ALU/lt1_c25 ),
    .fco(\u_EXU_ALU/lt1_c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_28|u_EXU_ALU/lt1_27  (
    .a(i_exu_op1[28:27]),
    .b(i_exu_op2[28:27]),
    .fci(\u_EXU_ALU/lt1_c27 ),
    .fco(\u_EXU_ALU/lt1_c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_2|u_EXU_ALU/lt1_1  (
    .a(i_exu_op1[2:1]),
    .b(i_exu_op2[2:1]),
    .fci(\u_EXU_ALU/lt1_c1 ),
    .fco(\u_EXU_ALU/lt1_c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_30|u_EXU_ALU/lt1_29  (
    .a(i_exu_op1[30:29]),
    .b(i_exu_op2[30:29]),
    .fci(\u_EXU_ALU/lt1_c29 ),
    .fco(\u_EXU_ALU/lt1_c31 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_4|u_EXU_ALU/lt1_3  (
    .a(i_exu_op1[4:3]),
    .b(i_exu_op2[4:3]),
    .fci(\u_EXU_ALU/lt1_c3 ),
    .fco(\u_EXU_ALU/lt1_c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_6|u_EXU_ALU/lt1_5  (
    .a(i_exu_op1[6:5]),
    .b(i_exu_op2[6:5]),
    .fci(\u_EXU_ALU/lt1_c5 ),
    .fco(\u_EXU_ALU/lt1_c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_8|u_EXU_ALU/lt1_7  (
    .a(i_exu_op1[8:7]),
    .b(i_exu_op2[8:7]),
    .fci(\u_EXU_ALU/lt1_c7 ),
    .fco(\u_EXU_ALU/lt1_c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_ALU/lt1_0|u_EXU_ALU/lt1_cin"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_EXU_ALU/lt1_cout|u_EXU_ALU/lt1_31  (
    .a({1'b0,i_exu_op1[31]}),
    .b({1'b1,i_exu_op2[31]}),
    .fci(\u_EXU_ALU/lt1_c31 ),
    .f({\u_EXU_ALU/n261 ,open_n988}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/sub0/ucin_al_u1478"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/sub0/u11_al_u1481  (
    .a({i_exu_op1[13],i_exu_op1[11]}),
    .b({i_exu_op1[14],i_exu_op1[12]}),
    .c(2'b11),
    .d({i_exu_op2[13],i_exu_op2[11]}),
    .e({i_exu_op2[14],i_exu_op2[12]}),
    .fci(\u_EXU_ALU/sub0/c11 ),
    .f({\u_EXU_ALU/n33 [13],\u_EXU_ALU/n33 [11]}),
    .fco(\u_EXU_ALU/sub0/c15 ),
    .fx({\u_EXU_ALU/n33 [14],\u_EXU_ALU/n33 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/sub0/ucin_al_u1478"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/sub0/u15_al_u1482  (
    .a({i_exu_op1[17],i_exu_op1[15]}),
    .b({i_exu_op1[18],i_exu_op1[16]}),
    .c(2'b11),
    .d({i_exu_op2[17],i_exu_op2[15]}),
    .e({i_exu_op2[18],i_exu_op2[16]}),
    .fci(\u_EXU_ALU/sub0/c15 ),
    .f({\u_EXU_ALU/n33 [17],\u_EXU_ALU/n33 [15]}),
    .fco(\u_EXU_ALU/sub0/c19 ),
    .fx({\u_EXU_ALU/n33 [18],\u_EXU_ALU/n33 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/sub0/ucin_al_u1478"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/sub0/u19_al_u1483  (
    .a({i_exu_op1[21],i_exu_op1[19]}),
    .b({i_exu_op1[22],i_exu_op1[20]}),
    .c(2'b11),
    .d({i_exu_op2[21],i_exu_op2[19]}),
    .e({i_exu_op2[22],i_exu_op2[20]}),
    .fci(\u_EXU_ALU/sub0/c19 ),
    .f({\u_EXU_ALU/n33 [21],\u_EXU_ALU/n33 [19]}),
    .fco(\u_EXU_ALU/sub0/c23 ),
    .fx({\u_EXU_ALU/n33 [22],\u_EXU_ALU/n33 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/sub0/ucin_al_u1478"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/sub0/u23_al_u1484  (
    .a({i_exu_op1[25],i_exu_op1[23]}),
    .b({i_exu_op1[26],i_exu_op1[24]}),
    .c(2'b11),
    .d({i_exu_op2[25],i_exu_op2[23]}),
    .e({i_exu_op2[26],i_exu_op2[24]}),
    .fci(\u_EXU_ALU/sub0/c23 ),
    .f({\u_EXU_ALU/n33 [25],\u_EXU_ALU/n33 [23]}),
    .fco(\u_EXU_ALU/sub0/c27 ),
    .fx({\u_EXU_ALU/n33 [26],\u_EXU_ALU/n33 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/sub0/ucin_al_u1478"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/sub0/u27_al_u1485  (
    .a({i_exu_op1[29],i_exu_op1[27]}),
    .b({i_exu_op1[30],i_exu_op1[28]}),
    .c(2'b11),
    .d({i_exu_op2[29],i_exu_op2[27]}),
    .e({i_exu_op2[30],i_exu_op2[28]}),
    .fci(\u_EXU_ALU/sub0/c27 ),
    .f({\u_EXU_ALU/n33 [29],\u_EXU_ALU/n33 [27]}),
    .fco(\u_EXU_ALU/sub0/c31 ),
    .fx({\u_EXU_ALU/n33 [30],\u_EXU_ALU/n33 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/sub0/ucin_al_u1478"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/sub0/u31_al_u1486  (
    .a({open_n1084,i_exu_op1[31]}),
    .c(2'b11),
    .d({open_n1089,i_exu_op2[31]}),
    .fci(\u_EXU_ALU/sub0/c31 ),
    .f({open_n1106,\u_EXU_ALU/n33 [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/sub0/ucin_al_u1478"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/sub0/u3_al_u1479  (
    .a({i_exu_op1[5],i_exu_op1[3]}),
    .b({i_exu_op1[6],i_exu_op1[4]}),
    .c(2'b11),
    .d({i_exu_op2[5],i_exu_op2[3]}),
    .e({i_exu_op2[6],i_exu_op2[4]}),
    .fci(\u_EXU_ALU/sub0/c3 ),
    .f({\u_EXU_ALU/n33 [5],\u_EXU_ALU/n33 [3]}),
    .fco(\u_EXU_ALU/sub0/c7 ),
    .fx({\u_EXU_ALU/n33 [6],\u_EXU_ALU/n33 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/sub0/ucin_al_u1478"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/sub0/u7_al_u1480  (
    .a({i_exu_op1[9],i_exu_op1[7]}),
    .b({i_exu_op1[10],i_exu_op1[8]}),
    .c(2'b11),
    .d({i_exu_op2[9],i_exu_op2[7]}),
    .e({i_exu_op2[10],i_exu_op2[8]}),
    .fci(\u_EXU_ALU/sub0/c7 ),
    .f({\u_EXU_ALU/n33 [9],\u_EXU_ALU/n33 [7]}),
    .fco(\u_EXU_ALU/sub0/c11 ),
    .fx({\u_EXU_ALU/n33 [10],\u_EXU_ALU/n33 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_ALU/sub0/ucin_al_u1478"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_ALU/sub0/ucin_al_u1478  (
    .a({i_exu_op1[1],1'b0}),
    .b({i_exu_op1[2],i_exu_op1[0]}),
    .c(2'b11),
    .d({i_exu_op2[1],1'b1}),
    .e({i_exu_op2[2],i_exu_op2[0]}),
    .f({\u_EXU_ALU/n33 [1],open_n1165}),
    .fco(\u_EXU_ALU/sub0/c3 ),
    .fx({\u_EXU_ALU/n33 [2],\u_EXU_ALU/n33 [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add0/ucin_al_u1487"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add0/u11_al_u1490  (
    .a({i_iaddr[13],i_iaddr[11]}),
    .b({i_iaddr[14],i_iaddr[12]}),
    .c(2'b00),
    .d({i_imm[13],i_imm[11]}),
    .e({i_imm[14],i_imm[12]}),
    .fci(\u_EXU_BJU/add0/c11 ),
    .f({\u_EXU_BJU/bxx_nxtpc [13],\u_EXU_BJU/bxx_nxtpc [11]}),
    .fco(\u_EXU_BJU/add0/c15 ),
    .fx({\u_EXU_BJU/bxx_nxtpc [14],\u_EXU_BJU/bxx_nxtpc [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add0/ucin_al_u1487"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add0/u15_al_u1491  (
    .a({i_iaddr[17],i_iaddr[15]}),
    .b({i_iaddr[18],i_iaddr[16]}),
    .c(2'b00),
    .d({i_imm[17],i_imm[15]}),
    .e({i_imm[18],i_imm[16]}),
    .fci(\u_EXU_BJU/add0/c15 ),
    .f({\u_EXU_BJU/bxx_nxtpc [17],\u_EXU_BJU/bxx_nxtpc [15]}),
    .fco(\u_EXU_BJU/add0/c19 ),
    .fx({\u_EXU_BJU/bxx_nxtpc [18],\u_EXU_BJU/bxx_nxtpc [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add0/ucin_al_u1487"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add0/u19_al_u1492  (
    .a({i_iaddr[21],i_iaddr[19]}),
    .b({i_iaddr[22],i_iaddr[20]}),
    .c(2'b00),
    .d({i_imm[21],i_imm[19]}),
    .e({i_imm[22],i_imm[20]}),
    .fci(\u_EXU_BJU/add0/c19 ),
    .f({\u_EXU_BJU/bxx_nxtpc [21],\u_EXU_BJU/bxx_nxtpc [19]}),
    .fco(\u_EXU_BJU/add0/c23 ),
    .fx({\u_EXU_BJU/bxx_nxtpc [22],\u_EXU_BJU/bxx_nxtpc [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add0/ucin_al_u1487"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add0/u23_al_u1493  (
    .a({i_iaddr[25],i_iaddr[23]}),
    .b({i_iaddr[26],i_iaddr[24]}),
    .c(2'b00),
    .d({i_imm[25],i_imm[23]}),
    .e({i_imm[26],i_imm[24]}),
    .fci(\u_EXU_BJU/add0/c23 ),
    .f({\u_EXU_BJU/bxx_nxtpc [25],\u_EXU_BJU/bxx_nxtpc [23]}),
    .fco(\u_EXU_BJU/add0/c27 ),
    .fx({\u_EXU_BJU/bxx_nxtpc [26],\u_EXU_BJU/bxx_nxtpc [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add0/ucin_al_u1487"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add0/u27_al_u1494  (
    .a({i_iaddr[29],i_iaddr[27]}),
    .b({i_iaddr[30],i_iaddr[28]}),
    .c(2'b00),
    .d({i_imm[29],i_imm[27]}),
    .e({i_imm[30],i_imm[28]}),
    .fci(\u_EXU_BJU/add0/c27 ),
    .f({\u_EXU_BJU/bxx_nxtpc [29],\u_EXU_BJU/bxx_nxtpc [27]}),
    .fco(\u_EXU_BJU/add0/c31 ),
    .fx({\u_EXU_BJU/bxx_nxtpc [30],\u_EXU_BJU/bxx_nxtpc [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add0/ucin_al_u1487"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add0/u31_al_u1495  (
    .a({open_n1258,i_iaddr[31]}),
    .c(2'b00),
    .d({open_n1263,i_imm[31]}),
    .fci(\u_EXU_BJU/add0/c31 ),
    .f({open_n1280,\u_EXU_BJU/bxx_nxtpc [31]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add0/ucin_al_u1487"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add0/u3_al_u1488  (
    .a({i_iaddr[5],i_iaddr[3]}),
    .b({i_iaddr[6],i_iaddr[4]}),
    .c(2'b00),
    .d({i_imm[5],i_imm[3]}),
    .e({i_imm[6],i_imm[4]}),
    .fci(\u_EXU_BJU/add0/c3 ),
    .f({\u_EXU_BJU/bxx_nxtpc [5],\u_EXU_BJU/bxx_nxtpc [3]}),
    .fco(\u_EXU_BJU/add0/c7 ),
    .fx({\u_EXU_BJU/bxx_nxtpc [6],\u_EXU_BJU/bxx_nxtpc [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add0/ucin_al_u1487"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add0/u7_al_u1489  (
    .a({i_iaddr[9],i_iaddr[7]}),
    .b({i_iaddr[10],i_iaddr[8]}),
    .c(2'b00),
    .d({i_imm[9],i_imm[7]}),
    .e({i_imm[10],i_imm[8]}),
    .fci(\u_EXU_BJU/add0/c7 ),
    .f({\u_EXU_BJU/bxx_nxtpc [9],\u_EXU_BJU/bxx_nxtpc [7]}),
    .fco(\u_EXU_BJU/add0/c11 ),
    .fx({\u_EXU_BJU/bxx_nxtpc [10],\u_EXU_BJU/bxx_nxtpc [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add0/ucin_al_u1487"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add0/ucin_al_u1487  (
    .a({i_iaddr[1],1'b0}),
    .b({i_iaddr[2],i_iaddr[0]}),
    .c(2'b00),
    .d({i_imm[1],1'b1}),
    .e({i_imm[2],i_imm[0]}),
    .f({\u_EXU_BJU/bxx_nxtpc [1],open_n1339}),
    .fco(\u_EXU_BJU/add0/c3 ),
    .fx({\u_EXU_BJU/bxx_nxtpc [2],\u_EXU_BJU/bxx_nxtpc [0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add1/ucin_al_u1496"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add1/u11_al_u1499  (
    .a({i_iaddr[15],i_iaddr[13]}),
    .b({i_iaddr[16],i_iaddr[14]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_EXU_BJU/add1/c11 ),
    .f({bju_rdwdata[15],bju_rdwdata[13]}),
    .fco(\u_EXU_BJU/add1/c15 ),
    .fx({bju_rdwdata[16],bju_rdwdata[14]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add1/ucin_al_u1496"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add1/u15_al_u1500  (
    .a({i_iaddr[19],i_iaddr[17]}),
    .b({i_iaddr[20],i_iaddr[18]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_EXU_BJU/add1/c15 ),
    .f({bju_rdwdata[19],bju_rdwdata[17]}),
    .fco(\u_EXU_BJU/add1/c19 ),
    .fx({bju_rdwdata[20],bju_rdwdata[18]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add1/ucin_al_u1496"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add1/u19_al_u1501  (
    .a({i_iaddr[23],i_iaddr[21]}),
    .b({i_iaddr[24],i_iaddr[22]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_EXU_BJU/add1/c19 ),
    .f({bju_rdwdata[23],bju_rdwdata[21]}),
    .fco(\u_EXU_BJU/add1/c23 ),
    .fx({bju_rdwdata[24],bju_rdwdata[22]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add1/ucin_al_u1496"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add1/u23_al_u1502  (
    .a({i_iaddr[27],i_iaddr[25]}),
    .b({i_iaddr[28],i_iaddr[26]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_EXU_BJU/add1/c23 ),
    .f({bju_rdwdata[27],bju_rdwdata[25]}),
    .fco(\u_EXU_BJU/add1/c27 ),
    .fx({bju_rdwdata[28],bju_rdwdata[26]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add1/ucin_al_u1496"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add1/u27_al_u1503  (
    .a({i_iaddr[31],i_iaddr[29]}),
    .b({open_n1414,i_iaddr[30]}),
    .c(2'b00),
    .d(2'b00),
    .e({open_n1417,1'b0}),
    .fci(\u_EXU_BJU/add1/c27 ),
    .f({bju_rdwdata[31],bju_rdwdata[29]}),
    .fx({open_n1433,bju_rdwdata[30]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add1/ucin_al_u1496"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add1/u3_al_u1497  (
    .a({i_iaddr[7],i_iaddr[5]}),
    .b({i_iaddr[8],i_iaddr[6]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_EXU_BJU/add1/c3 ),
    .f({bju_rdwdata[7],bju_rdwdata[5]}),
    .fco(\u_EXU_BJU/add1/c7 ),
    .fx({bju_rdwdata[8],bju_rdwdata[6]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add1/ucin_al_u1496"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add1/u7_al_u1498  (
    .a({i_iaddr[11],i_iaddr[9]}),
    .b({i_iaddr[12],i_iaddr[10]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\u_EXU_BJU/add1/c7 ),
    .f({bju_rdwdata[11],bju_rdwdata[9]}),
    .fco(\u_EXU_BJU/add1/c11 ),
    .fx({bju_rdwdata[12],bju_rdwdata[10]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_EXU_BJU/add1/ucin_al_u1496"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_EXU_BJU/add1/ucin_al_u1496  (
    .a({i_iaddr[3],1'b0}),
    .b({i_iaddr[4],i_iaddr[2]}),
    .c(2'b00),
    .d(2'b01),
    .e(2'b01),
    .f({bju_rdwdata[3],open_n1489}),
    .fco(\u_EXU_BJU/add1/c3 ),
    .fx({bju_rdwdata[4],bju_rdwdata[2]}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_EXU_LSU/access2_once_reg  (
    .clk(i_clk),
    .d(\u_EXU_LSU/n30 ),
    .sr(i_rstn),
    .q(\u_EXU_LSU/access2_once ));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_EXU_LSU/access2_vld_reg  (
    .clk(i_clk),
    .d(\u_EXU_LSU/n26 ),
    .sr(i_rstn),
    .q(\u_EXU_LSU/access2_vld ));  // ../RTL/core/exu_lsu.v(105)
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin  (
    .a({o_ribm_addr[2],1'b0}),
    .b({1'b1,open_n1494}),
    .f({\u_EXU_LSU/n59 [0],open_n1514}),
    .fco(\u_EXU_LSU/add0/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u10|u_EXU_LSU/add0/u9  (
    .a(o_ribm_addr[12:11]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c9 ),
    .f(\u_EXU_LSU/n59 [10:9]),
    .fco(\u_EXU_LSU/add0/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u12|u_EXU_LSU/add0/u11  (
    .a(o_ribm_addr[14:13]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c11 ),
    .f(\u_EXU_LSU/n59 [12:11]),
    .fco(\u_EXU_LSU/add0/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u14|u_EXU_LSU/add0/u13  (
    .a(o_ribm_addr[16:15]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c13 ),
    .f(\u_EXU_LSU/n59 [14:13]),
    .fco(\u_EXU_LSU/add0/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u16|u_EXU_LSU/add0/u15  (
    .a(o_ribm_addr[18:17]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c15 ),
    .f(\u_EXU_LSU/n59 [16:15]),
    .fco(\u_EXU_LSU/add0/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u18|u_EXU_LSU/add0/u17  (
    .a(o_ribm_addr[20:19]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c17 ),
    .f(\u_EXU_LSU/n59 [18:17]),
    .fco(\u_EXU_LSU/add0/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u20|u_EXU_LSU/add0/u19  (
    .a(o_ribm_addr[22:21]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c19 ),
    .f(\u_EXU_LSU/n59 [20:19]),
    .fco(\u_EXU_LSU/add0/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u22|u_EXU_LSU/add0/u21  (
    .a(o_ribm_addr[24:23]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c21 ),
    .f(\u_EXU_LSU/n59 [22:21]),
    .fco(\u_EXU_LSU/add0/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u24|u_EXU_LSU/add0/u23  (
    .a(o_ribm_addr[26:25]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c23 ),
    .f(\u_EXU_LSU/n59 [24:23]),
    .fco(\u_EXU_LSU/add0/c25 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u26|u_EXU_LSU/add0/u25  (
    .a(o_ribm_addr[28:27]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c25 ),
    .f(\u_EXU_LSU/n59 [26:25]),
    .fco(\u_EXU_LSU/add0/c27 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u28|u_EXU_LSU/add0/u27  (
    .a(o_ribm_addr[30:29]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c27 ),
    .f(\u_EXU_LSU/n59 [28:27]),
    .fco(\u_EXU_LSU/add0/c29 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u29_al_u1504  (
    .a({open_n1739,o_ribm_addr[31]}),
    .b({open_n1740,1'b0}),
    .fci(\u_EXU_LSU/add0/c29 ),
    .f({open_n1759,\u_EXU_LSU/n59 [29]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u2|u_EXU_LSU/add0/u1  (
    .a(o_ribm_addr[4:3]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c1 ),
    .f(\u_EXU_LSU/n59 [2:1]),
    .fco(\u_EXU_LSU/add0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u4|u_EXU_LSU/add0/u3  (
    .a(o_ribm_addr[6:5]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c3 ),
    .f(\u_EXU_LSU/n59 [4:3]),
    .fco(\u_EXU_LSU/add0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u6|u_EXU_LSU/add0/u5  (
    .a(o_ribm_addr[8:7]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c5 ),
    .f(\u_EXU_LSU/n59 [6:5]),
    .fco(\u_EXU_LSU/add0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_EXU_LSU/add0/u0|u_EXU_LSU/add0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_EXU_LSU/add0/u8|u_EXU_LSU/add0/u7  (
    .a(o_ribm_addr[10:9]),
    .b(2'b00),
    .fci(\u_EXU_LSU/add0/c7 ),
    .f(\u_EXU_LSU/n59 [8:7]),
    .fco(\u_EXU_LSU/add0/c9 ));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_EXU_LSU/handshake_once_reg  (
    .clk(i_clk),
    .d(\u_EXU_LSU/n80 ),
    .sr(i_rstn),
    .q(\u_EXU_LSU/handshake_once ));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_EXU_LSU/handshake_rdy_last_reg  (
    .ce(\u_EXU_LSU/n1 ),
    .clk(i_clk),
    .d(i_ribm_gnt),
    .sr(i_rstn),
    .q(\u_EXU_LSU/handshake_rdy_last ));  // ../RTL/core/exu_lsu.v(73)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_EXU_LSU/o_ribm_req_reg  (
    .clk(i_clk),
    .d(\u_EXU_LSU/n75 ),
    .sr(i_rstn),
    .q(o_ribm_req));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/o_ribm_wrcs_reg  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_decinfo[1]),
    .q(o_ribm_wrcs));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_EXU_LSU/rdwen_reg  (
    .clk(i_clk),
    .d(\u_EXU_LSU/n23 ),
    .sr(i_rstn),
    .q(o_exu_rdwen2));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg0_b0  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(o_rdidx0[0]),
    .q(o_rdidx2[0]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg0_b1  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(o_rdidx0[1]),
    .q(o_rdidx2[1]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg0_b2  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(o_rdidx0[2]),
    .q(o_rdidx2[2]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg0_b3  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(o_rdidx0[3]),
    .q(o_rdidx2[3]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg0_b4  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(o_rdidx0[4]),
    .q(o_rdidx2[4]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg1_b0  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(alu2lsu_result[0]),
    .q(\u_EXU_LSU/align_mode_reg [0]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg1_b1  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(alu2lsu_result[1]),
    .q(\u_EXU_LSU/align_mode_reg [1]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b10  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[10]),
    .q(\u_EXU_LSU/rs2rdata_reg [10]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b11  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[11]),
    .q(\u_EXU_LSU/rs2rdata_reg [11]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b12  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[12]),
    .q(\u_EXU_LSU/rs2rdata_reg [12]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b13  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[13]),
    .q(\u_EXU_LSU/rs2rdata_reg [13]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b14  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[14]),
    .q(\u_EXU_LSU/rs2rdata_reg [14]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b15  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[15]),
    .q(\u_EXU_LSU/rs2rdata_reg [15]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b16  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[16]),
    .q(\u_EXU_LSU/rs2rdata_reg [16]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b17  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[17]),
    .q(\u_EXU_LSU/rs2rdata_reg [17]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b18  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[18]),
    .q(\u_EXU_LSU/rs2rdata_reg [18]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b19  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[19]),
    .q(\u_EXU_LSU/rs2rdata_reg [19]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b20  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[20]),
    .q(\u_EXU_LSU/rs2rdata_reg [20]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b21  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[21]),
    .q(\u_EXU_LSU/rs2rdata_reg [21]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b22  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[22]),
    .q(\u_EXU_LSU/rs2rdata_reg [22]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b23  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[23]),
    .q(\u_EXU_LSU/rs2rdata_reg [23]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b24  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[24]),
    .q(\u_EXU_LSU/rs2rdata_reg [24]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b25  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[25]),
    .q(\u_EXU_LSU/rs2rdata_reg [25]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b26  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[26]),
    .q(\u_EXU_LSU/rs2rdata_reg [26]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b27  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[27]),
    .q(\u_EXU_LSU/rs2rdata_reg [27]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b28  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[28]),
    .q(\u_EXU_LSU/rs2rdata_reg [28]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b29  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[29]),
    .q(\u_EXU_LSU/rs2rdata_reg [29]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b30  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[30]),
    .q(\u_EXU_LSU/rs2rdata_reg [30]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b31  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[31]),
    .q(\u_EXU_LSU/rs2rdata_reg [31]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b8  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[8]),
    .q(\u_EXU_LSU/rs2rdata_reg [8]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg2_b9  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_rs2rdata[9]),
    .q(\u_EXU_LSU/rs2rdata_reg [9]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg3_b2  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_decinfo[2]),
    .q(\u_EXU_LSU/lsuinfo [2]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg3_b3  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_decinfo[3]),
    .q(\u_EXU_LSU/lsuinfo [3]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg3_b4  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_decinfo[4]),
    .q(\u_EXU_LSU/lsuinfo [4]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg3_b5  (
    .ce(\u_EXU_LSU/mux10_b2_sel_is_2_o ),
    .clk(i_clk),
    .d(i_decinfo[5]),
    .q(\u_EXU_LSU/lsuinfo [5]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b0  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[0]),
    .q(\u_EXU_LSU/overleft_buffer [0]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b1  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[1]),
    .q(\u_EXU_LSU/overleft_buffer [1]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b10  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[10]),
    .q(\u_EXU_LSU/overleft_buffer [10]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b11  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[11]),
    .q(\u_EXU_LSU/overleft_buffer [11]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b12  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[12]),
    .q(\u_EXU_LSU/overleft_buffer [12]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b13  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[13]),
    .q(\u_EXU_LSU/overleft_buffer [13]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b14  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[14]),
    .q(\u_EXU_LSU/overleft_buffer [14]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b15  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[15]),
    .q(\u_EXU_LSU/overleft_buffer [15]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b16  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[16]),
    .q(\u_EXU_LSU/overleft_buffer [16]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b17  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[17]),
    .q(\u_EXU_LSU/overleft_buffer [17]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b18  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[18]),
    .q(\u_EXU_LSU/overleft_buffer [18]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b19  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[19]),
    .q(\u_EXU_LSU/overleft_buffer [19]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b2  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[2]),
    .q(\u_EXU_LSU/overleft_buffer [2]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b20  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[20]),
    .q(\u_EXU_LSU/overleft_buffer [20]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b21  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[21]),
    .q(\u_EXU_LSU/overleft_buffer [21]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b22  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[22]),
    .q(\u_EXU_LSU/overleft_buffer [22]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b23  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[23]),
    .q(\u_EXU_LSU/overleft_buffer [23]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b24  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[24]),
    .q(\u_EXU_LSU/overleft_buffer [24]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b25  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[25]),
    .q(\u_EXU_LSU/overleft_buffer [25]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b26  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[26]),
    .q(\u_EXU_LSU/overleft_buffer [26]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b27  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[27]),
    .q(\u_EXU_LSU/overleft_buffer [27]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b28  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[28]),
    .q(\u_EXU_LSU/overleft_buffer [28]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b29  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[29]),
    .q(\u_EXU_LSU/overleft_buffer [29]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b3  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[3]),
    .q(\u_EXU_LSU/overleft_buffer [3]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b30  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[30]),
    .q(\u_EXU_LSU/overleft_buffer [30]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b31  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[31]),
    .q(\u_EXU_LSU/overleft_buffer [31]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b4  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[4]),
    .q(\u_EXU_LSU/overleft_buffer [4]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b5  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[5]),
    .q(\u_EXU_LSU/overleft_buffer [5]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b6  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[6]),
    .q(\u_EXU_LSU/overleft_buffer [6]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b7  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[7]),
    .q(\u_EXU_LSU/overleft_buffer [7]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b8  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[8]),
    .q(\u_EXU_LSU/overleft_buffer [8]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg4_b9  (
    .ce(\u_EXU_LSU/mux11_b0_sel_is_2_o ),
    .clk(i_clk),
    .d(i_ribm_rdata[9]),
    .q(\u_EXU_LSU/overleft_buffer [9]));  // ../RTL/core/exu_lsu.v(105)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b10  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [10]),
    .q(o_ribm_addr[10]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b11  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [11]),
    .q(o_ribm_addr[11]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b12  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [12]),
    .q(o_ribm_addr[12]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b13  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [13]),
    .q(o_ribm_addr[13]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b14  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [14]),
    .q(o_ribm_addr[14]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b15  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [15]),
    .q(o_ribm_addr[15]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b16  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [16]),
    .q(o_ribm_addr[16]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b17  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [17]),
    .q(o_ribm_addr[17]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b18  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [18]),
    .q(o_ribm_addr[18]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b19  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [19]),
    .q(o_ribm_addr[19]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b2  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [2]),
    .q(o_ribm_addr[2]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b20  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [20]),
    .q(o_ribm_addr[20]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b21  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [21]),
    .q(o_ribm_addr[21]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b22  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [22]),
    .q(o_ribm_addr[22]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b23  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [23]),
    .q(o_ribm_addr[23]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b24  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [24]),
    .q(o_ribm_addr[24]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b25  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [25]),
    .q(o_ribm_addr[25]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b26  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [26]),
    .q(o_ribm_addr[26]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b27  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [27]),
    .q(o_ribm_addr[27]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b28  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [28]),
    .q(o_ribm_addr[28]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b29  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [29]),
    .q(o_ribm_addr[29]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b3  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [3]),
    .q(o_ribm_addr[3]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b30  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [30]),
    .q(o_ribm_addr[30]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b31  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [31]),
    .q(o_ribm_addr[31]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b4  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [4]),
    .q(o_ribm_addr[4]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b5  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [5]),
    .q(o_ribm_addr[5]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b6  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [6]),
    .q(o_ribm_addr[6]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b7  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [7]),
    .q(o_ribm_addr[7]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b8  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [8]),
    .q(o_ribm_addr[8]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg5_b9  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n76 [9]),
    .q(o_ribm_addr[9]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg6_b0  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n78 [0]),
    .q(o_ribm_mask[0]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg6_b1  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n78 [1]),
    .q(o_ribm_mask[1]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg6_b2  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n78 [2]),
    .q(o_ribm_mask[2]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg6_b3  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n78 [3]),
    .q(o_ribm_mask[3]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b0  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [0]),
    .q(o_ribm_wdata[0]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b1  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [1]),
    .q(o_ribm_wdata[1]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b10  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [10]),
    .q(o_ribm_wdata[10]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b11  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [11]),
    .q(o_ribm_wdata[11]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b12  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [12]),
    .q(o_ribm_wdata[12]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b13  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [13]),
    .q(o_ribm_wdata[13]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b14  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [14]),
    .q(o_ribm_wdata[14]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b15  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [15]),
    .q(o_ribm_wdata[15]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b16  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [16]),
    .q(o_ribm_wdata[16]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b17  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [17]),
    .q(o_ribm_wdata[17]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b18  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [18]),
    .q(o_ribm_wdata[18]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b19  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [19]),
    .q(o_ribm_wdata[19]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b2  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [2]),
    .q(o_ribm_wdata[2]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b20  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [20]),
    .q(o_ribm_wdata[20]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b21  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [21]),
    .q(o_ribm_wdata[21]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b22  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [22]),
    .q(o_ribm_wdata[22]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b23  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [23]),
    .q(o_ribm_wdata[23]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b24  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [24]),
    .q(o_ribm_wdata[24]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b25  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [25]),
    .q(o_ribm_wdata[25]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b26  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [26]),
    .q(o_ribm_wdata[26]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b27  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [27]),
    .q(o_ribm_wdata[27]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b28  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [28]),
    .q(o_ribm_wdata[28]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b29  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [29]),
    .q(o_ribm_wdata[29]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b3  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [3]),
    .q(o_ribm_wdata[3]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b30  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [30]),
    .q(o_ribm_wdata[30]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b31  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [31]),
    .q(o_ribm_wdata[31]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b4  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [4]),
    .q(o_ribm_wdata[4]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b5  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [5]),
    .q(o_ribm_wdata[5]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b6  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [6]),
    .q(o_ribm_wdata[6]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b7  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [7]),
    .q(o_ribm_wdata[7]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b8  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [8]),
    .q(o_ribm_wdata[8]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_EXU_LSU/reg7_b9  (
    .ce(i_rstn),
    .clk(i_clk),
    .d(\u_EXU_LSU/n79 [9]),
    .q(o_ribm_wdata[9]));  // ../RTL/core/exu_lsu.v(156)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_EXU_LSU/working_reg  (
    .clk(i_clk),
    .d(\u_EXU_LSU/n25 ),
    .sr(i_rstn),
    .q(\u_EXU_LSU/working ));  // ../RTL/core/exu_lsu.v(105)
  EXU_MDU u_EXU_MDU (
    .i_clk(i_clk),
    .i_decinfo_grp(i_decinfo_grp),
    .i_flush(mdu_flush),
    .i_mdu_op1(i_exu_op1),
    .i_mdu_op2(i_exu_op2),
    .i_mdu_rdidx(o_rdidx0),
    .i_mdu_rdwen(o_exu_rdwen0),
    .i_mduinfo({i_decinfo[9:1],1'b0}),
    .i_rstn(i_rstn),
    .i_vld(i_vld),
    .o_mdu_rdidx(o_rdidx1),
    .o_mdu_rdwdata(o_rdwdata1),
    .o_mdu_rdwen(o_rdwen1),
    .o_will_rdidx(o_exu_rdidx1),
    .o_will_rdwen(o_exu_rdwen1),
    .o_working(o_mdu_working));  // ../RTL/core/exu.v(176)

endmodule 

module REGFILE  // ../RTL/core/regfile.v(12)
  (
  i_clk,
  i_rd_wdata,
  i_rdidx,
  i_rdwen,
  i_rs1idx,
  i_rs1ren,
  i_rs2idx,
  i_rs2ren,
  i_rstn,
  o_rs1_rdata,
  o_rs2_rdata
  );

  input i_clk;  // ../RTL/core/regfile.v(13)
  input [31:0] i_rd_wdata;  // ../RTL/core/regfile.v(17)
  input [4:0] i_rdidx;  // ../RTL/core/regfile.v(16)
  input i_rdwen;  // ../RTL/core/regfile.v(15)
  input [4:0] i_rs1idx;  // ../RTL/core/regfile.v(19)
  input i_rs1ren;  // ../RTL/core/regfile.v(18)
  input [4:0] i_rs2idx;  // ../RTL/core/regfile.v(22)
  input i_rs2ren;  // ../RTL/core/regfile.v(21)
  input i_rstn;  // ../RTL/core/regfile.v(14)
  output [31:0] o_rs1_rdata;  // ../RTL/core/regfile.v(20)
  output [31:0] o_rs2_rdata;  // ../RTL/core/regfile.v(23)

  // localparam gen_regfile_rd[0].i = 0;
  // localparam gen_regfile_rd[10].i = 10;
  // localparam gen_regfile_rd[11].i = 11;
  // localparam gen_regfile_rd[12].i = 12;
  // localparam gen_regfile_rd[13].i = 13;
  // localparam gen_regfile_rd[14].i = 14;
  // localparam gen_regfile_rd[15].i = 15;
  // localparam gen_regfile_rd[16].i = 16;
  // localparam gen_regfile_rd[17].i = 17;
  // localparam gen_regfile_rd[18].i = 18;
  // localparam gen_regfile_rd[19].i = 19;
  // localparam gen_regfile_rd[1].i = 1;
  // localparam gen_regfile_rd[20].i = 20;
  // localparam gen_regfile_rd[21].i = 21;
  // localparam gen_regfile_rd[22].i = 22;
  // localparam gen_regfile_rd[23].i = 23;
  // localparam gen_regfile_rd[24].i = 24;
  // localparam gen_regfile_rd[25].i = 25;
  // localparam gen_regfile_rd[26].i = 26;
  // localparam gen_regfile_rd[27].i = 27;
  // localparam gen_regfile_rd[28].i = 28;
  // localparam gen_regfile_rd[29].i = 29;
  // localparam gen_regfile_rd[2].i = 2;
  // localparam gen_regfile_rd[30].i = 30;
  // localparam gen_regfile_rd[31].i = 31;
  // localparam gen_regfile_rd[3].i = 3;
  // localparam gen_regfile_rd[4].i = 4;
  // localparam gen_regfile_rd[5].i = 5;
  // localparam gen_regfile_rd[6].i = 6;
  // localparam gen_regfile_rd[7].i = 7;
  // localparam gen_regfile_rd[8].i = 8;
  // localparam gen_regfile_rd[9].i = 9;
  wire  \mux31_b0/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b0/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b0/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b0/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b0/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b0/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b0/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b0/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b1/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b10/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b11/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b12/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b12/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b12/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b12/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b12/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b12/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b12/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b12/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b13/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b13/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b13/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b13/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b13/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b13/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b13/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b13/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b14/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b14/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b14/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b14/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b14/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b14/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b14/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b14/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b15/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b15/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b15/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b15/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b15/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b15/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b15/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b15/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b16/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b16/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b16/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b16/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b16/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b16/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b16/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b16/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b17/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b19/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b2/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b2/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b2/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b20/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b21/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b22/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b23/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b23/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b23/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b23/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b23/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b23/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b23/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b23/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b24/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b24/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b24/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b24/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b24/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b24/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b24/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b24/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b26/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b26/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b26/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b26/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b26/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b26/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b26/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b26/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b28/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b28/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b28/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b28/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b28/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b28/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b28/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b28/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b29/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b29/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b29/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b29/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b29/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b29/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b29/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b29/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b3/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b30/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b30/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b30/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b30/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b30/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b30/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b30/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b30/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b31/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b31/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b31/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b31/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b31/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b31/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b4/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b4/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b4/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b4/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b4/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b4/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b4/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b4/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b5/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b6/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b7/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b7/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b7/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b8/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b8/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b8/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b8/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b8/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b8/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b8/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b8/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b9/B1_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b9/B1_2 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b9/B1_3 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b9/B1_4 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b9/B1_5 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b9/B1_6 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b9/B1_7 ;  // ../RTL/core/regfile.v(46)
  wire  \mux31_b9/B3_1 ;  // ../RTL/core/regfile.v(46)
  wire  \mux34_b0/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b0/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b0/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b0/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b0/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b0/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b0/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b1/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b10/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b10/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b10/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b11/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b11/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b11/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b12/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b12/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b12/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b12/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b12/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b12/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b12/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b12/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b13/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b13/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b13/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b13/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b13/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b13/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b13/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b13/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b14/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b14/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b14/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b14/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b14/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b14/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b14/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b14/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b15/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b15/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b15/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b15/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b15/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b15/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b15/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b15/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b16/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b17/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b17/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b17/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b17/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b17/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b17/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b17/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b17/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b18/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b18/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b18/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b18/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b18/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b18/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b18/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b18/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b19/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b19/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b19/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b2/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b20/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b21/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b22/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b22/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b22/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b22/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b22/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b22/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b22/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b22/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b23/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b23/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b23/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b23/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b23/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b23/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b24/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b24/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b24/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b24/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b24/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b24/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b24/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b24/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b25/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b25/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b25/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b25/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b25/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b25/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b25/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b25/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b26/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b26/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b26/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b27/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b27/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b27/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b27/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b27/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b27/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b27/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b27/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b28/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b28/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b28/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b28/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b28/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b28/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b28/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b28/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b29/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b29/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b29/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b29/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b29/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b29/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b3/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b3/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b3/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b30/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b30/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b30/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b30/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b30/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b30/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b30/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b30/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b31/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b31/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b31/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b31/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b31/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b31/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b31/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b31/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b4/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b5/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b5/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b5/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b5/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b5/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b5/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b6/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b6/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b6/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b6/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b6/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b6/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b6/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b6/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b7/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b7/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b7/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b7/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b7/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b7/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b7/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b7/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b8/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b8/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b8/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b8/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b8/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b8/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b9/B1_1 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b9/B1_2 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b9/B1_3 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b9/B1_4 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b9/B1_5 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b9/B1_6 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b9/B1_7 ;  // ../RTL/core/regfile.v(47)
  wire  \mux34_b9/B3_1 ;  // ../RTL/core/regfile.v(47)
  wire [31:0] \rfxs[10] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[11] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[12] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[13] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[14] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[15] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[16] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[17] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[18] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[19] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[1] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[20] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[21] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[22] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[23] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[24] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[25] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[26] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[27] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[28] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[29] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[2] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[30] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[31] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[3] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[4] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[5] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[6] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[7] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[8] ;  // ../RTL/core/regfile.v(27)
  wire [31:0] \rfxs[9] ;  // ../RTL/core/regfile.v(27)
  wire _al_u1001_o;
  wire _al_u1003_o;
  wire _al_u1005_o;
  wire _al_u1006_o;
  wire _al_u1008_o;
  wire _al_u1010_o;
  wire _al_u1012_o;
  wire _al_u1014_o;
  wire _al_u1016_o;
  wire _al_u1018_o;
  wire _al_u1019_o;
  wire _al_u1021_o;
  wire _al_u1022_o;
  wire _al_u1023_o;
  wire _al_u1024_o;
  wire _al_u1025_o;
  wire _al_u1026_o;
  wire _al_u1027_o;
  wire _al_u1028_o;
  wire _al_u1029_o;
  wire _al_u1030_o;
  wire _al_u1032_o;
  wire _al_u1033_o;
  wire _al_u1034_o;
  wire _al_u1035_o;
  wire _al_u1037_o;
  wire _al_u1039_o;
  wire _al_u1040_o;
  wire _al_u1042_o;
  wire _al_u1044_o;
  wire _al_u1046_o;
  wire _al_u1048_o;
  wire _al_u1050_o;
  wire _al_u1052_o;
  wire _al_u1053_o;
  wire _al_u1055_o;
  wire _al_u1056_o;
  wire _al_u1057_o;
  wire _al_u1058_o;
  wire _al_u1059_o;
  wire _al_u1061_o;
  wire _al_u1063_o;
  wire _al_u1065_o;
  wire _al_u1067_o;
  wire _al_u1069_o;
  wire _al_u1071_o;
  wire _al_u1072_o;
  wire _al_u1074_o;
  wire _al_u1076_o;
  wire _al_u1078_o;
  wire _al_u1080_o;
  wire _al_u1082_o;
  wire _al_u1084_o;
  wire _al_u1085_o;
  wire _al_u1087_o;
  wire _al_u1089_o;
  wire _al_u108_o;
  wire _al_u1091_o;
  wire _al_u1092_o;
  wire _al_u1093_o;
  wire _al_u1094_o;
  wire _al_u1095_o;
  wire _al_u1096_o;
  wire _al_u1098_o;
  wire _al_u1099_o;
  wire _al_u109_o;
  wire _al_u1100_o;
  wire _al_u1101_o;
  wire _al_u1102_o;
  wire _al_u1103_o;
  wire _al_u1104_o;
  wire _al_u1105_o;
  wire _al_u1106_o;
  wire _al_u1108_o;
  wire _al_u1110_o;
  wire _al_u1112_o;
  wire _al_u1114_o;
  wire _al_u1116_o;
  wire _al_u1118_o;
  wire _al_u1119_o;
  wire _al_u111_o;
  wire _al_u1121_o;
  wire _al_u1123_o;
  wire _al_u1125_o;
  wire _al_u1127_o;
  wire _al_u1129_o;
  wire _al_u112_o;
  wire _al_u1131_o;
  wire _al_u1132_o;
  wire _al_u1134_o;
  wire _al_u1136_o;
  wire _al_u1138_o;
  wire _al_u113_o;
  wire _al_u1140_o;
  wire _al_u1142_o;
  wire _al_u1144_o;
  wire _al_u1145_o;
  wire _al_u1147_o;
  wire _al_u1148_o;
  wire _al_u1149_o;
  wire _al_u114_o;
  wire _al_u1150_o;
  wire _al_u1151_o;
  wire _al_u1153_o;
  wire _al_u1155_o;
  wire _al_u1157_o;
  wire _al_u1159_o;
  wire _al_u115_o;
  wire _al_u1161_o;
  wire _al_u1163_o;
  wire _al_u1164_o;
  wire _al_u1166_o;
  wire _al_u1167_o;
  wire _al_u1168_o;
  wire _al_u1169_o;
  wire _al_u116_o;
  wire _al_u1170_o;
  wire _al_u1171_o;
  wire _al_u1172_o;
  wire _al_u1173_o;
  wire _al_u1174_o;
  wire _al_u1175_o;
  wire _al_u1177_o;
  wire _al_u1178_o;
  wire _al_u1179_o;
  wire _al_u117_o;
  wire _al_u1180_o;
  wire _al_u1181_o;
  wire _al_u1182_o;
  wire _al_u1183_o;
  wire _al_u1184_o;
  wire _al_u1185_o;
  wire _al_u1187_o;
  wire _al_u1188_o;
  wire _al_u1189_o;
  wire _al_u1190_o;
  wire _al_u1191_o;
  wire _al_u1192_o;
  wire _al_u1193_o;
  wire _al_u1194_o;
  wire _al_u1195_o;
  wire _al_u1196_o;
  wire _al_u1198_o;
  wire _al_u1199_o;
  wire _al_u119_o;
  wire _al_u1200_o;
  wire _al_u1201_o;
  wire _al_u1202_o;
  wire _al_u1203_o;
  wire _al_u1204_o;
  wire _al_u1205_o;
  wire _al_u1206_o;
  wire _al_u1208_o;
  wire _al_u1209_o;
  wire _al_u1210_o;
  wire _al_u1211_o;
  wire _al_u1212_o;
  wire _al_u1213_o;
  wire _al_u1214_o;
  wire _al_u1215_o;
  wire _al_u1216_o;
  wire _al_u1217_o;
  wire _al_u1219_o;
  wire _al_u121_o;
  wire _al_u1220_o;
  wire _al_u1221_o;
  wire _al_u1222_o;
  wire _al_u1223_o;
  wire _al_u1224_o;
  wire _al_u1225_o;
  wire _al_u1226_o;
  wire _al_u1227_o;
  wire _al_u1229_o;
  wire _al_u1230_o;
  wire _al_u1231_o;
  wire _al_u1232_o;
  wire _al_u1233_o;
  wire _al_u1234_o;
  wire _al_u1235_o;
  wire _al_u1236_o;
  wire _al_u1237_o;
  wire _al_u1238_o;
  wire _al_u123_o;
  wire _al_u1240_o;
  wire _al_u1241_o;
  wire _al_u1242_o;
  wire _al_u1243_o;
  wire _al_u1245_o;
  wire _al_u1247_o;
  wire _al_u1248_o;
  wire _al_u1250_o;
  wire _al_u1252_o;
  wire _al_u1254_o;
  wire _al_u1256_o;
  wire _al_u1258_o;
  wire _al_u125_o;
  wire _al_u1260_o;
  wire _al_u1261_o;
  wire _al_u1263_o;
  wire _al_u1265_o;
  wire _al_u1267_o;
  wire _al_u1269_o;
  wire _al_u126_o;
  wire _al_u1271_o;
  wire _al_u1273_o;
  wire _al_u1274_o;
  wire _al_u1276_o;
  wire _al_u1277_o;
  wire _al_u1278_o;
  wire _al_u1279_o;
  wire _al_u127_o;
  wire _al_u1280_o;
  wire _al_u1281_o;
  wire _al_u1282_o;
  wire _al_u1283_o;
  wire _al_u1284_o;
  wire _al_u1285_o;
  wire _al_u1287_o;
  wire _al_u1288_o;
  wire _al_u1289_o;
  wire _al_u1290_o;
  wire _al_u1291_o;
  wire _al_u1292_o;
  wire _al_u1293_o;
  wire _al_u1294_o;
  wire _al_u1295_o;
  wire _al_u1297_o;
  wire _al_u1299_o;
  wire _al_u129_o;
  wire _al_u1301_o;
  wire _al_u1303_o;
  wire _al_u1305_o;
  wire _al_u1307_o;
  wire _al_u1308_o;
  wire _al_u1310_o;
  wire _al_u1312_o;
  wire _al_u1314_o;
  wire _al_u1316_o;
  wire _al_u1318_o;
  wire _al_u131_o;
  wire _al_u1320_o;
  wire _al_u1321_o;
  wire _al_u1323_o;
  wire _al_u1325_o;
  wire _al_u1327_o;
  wire _al_u1329_o;
  wire _al_u1331_o;
  wire _al_u1333_o;
  wire _al_u1334_o;
  wire _al_u1336_o;
  wire _al_u1338_o;
  wire _al_u133_o;
  wire _al_u1340_o;
  wire _al_u1342_o;
  wire _al_u1344_o;
  wire _al_u1346_o;
  wire _al_u1347_o;
  wire _al_u1349_o;
  wire _al_u134_o;
  wire _al_u1351_o;
  wire _al_u1353_o;
  wire _al_u1354_o;
  wire _al_u1355_o;
  wire _al_u1356_o;
  wire _al_u1357_o;
  wire _al_u1358_o;
  wire _al_u1360_o;
  wire _al_u1361_o;
  wire _al_u1362_o;
  wire _al_u1363_o;
  wire _al_u1364_o;
  wire _al_u1365_o;
  wire _al_u1366_o;
  wire _al_u1367_o;
  wire _al_u1368_o;
  wire _al_u136_o;
  wire _al_u1370_o;
  wire _al_u1372_o;
  wire _al_u1374_o;
  wire _al_u1375_o;
  wire _al_u1376_o;
  wire _al_u1377_o;
  wire _al_u1378_o;
  wire _al_u1379_o;
  wire _al_u1381_o;
  wire _al_u1382_o;
  wire _al_u1383_o;
  wire _al_u1384_o;
  wire _al_u1385_o;
  wire _al_u1386_o;
  wire _al_u1387_o;
  wire _al_u1388_o;
  wire _al_u1389_o;
  wire _al_u138_o;
  wire _al_u1391_o;
  wire _al_u1392_o;
  wire _al_u1393_o;
  wire _al_u1394_o;
  wire _al_u1395_o;
  wire _al_u1396_o;
  wire _al_u1397_o;
  wire _al_u1398_o;
  wire _al_u1399_o;
  wire _al_u1401_o;
  wire _al_u1402_o;
  wire _al_u1403_o;
  wire _al_u1404_o;
  wire _al_u1405_o;
  wire _al_u1406_o;
  wire _al_u1407_o;
  wire _al_u1408_o;
  wire _al_u1409_o;
  wire _al_u140_o;
  wire _al_u1411_o;
  wire _al_u1413_o;
  wire _al_u1415_o;
  wire _al_u1417_o;
  wire _al_u1419_o;
  wire _al_u141_o;
  wire _al_u1420_o;
  wire _al_u1421_o;
  wire _al_u1422_o;
  wire _al_u1423_o;
  wire _al_u143_o;
  wire _al_u145_o;
  wire _al_u147_o;
  wire _al_u148_o;
  wire _al_u150_o;
  wire _al_u152_o;
  wire _al_u154_o;
  wire _al_u155_o;
  wire _al_u157_o;
  wire _al_u159_o;
  wire _al_u161_o;
  wire _al_u162_o;
  wire _al_u164_o;
  wire _al_u166_o;
  wire _al_u168_o;
  wire _al_u169_o;
  wire _al_u171_o;
  wire _al_u173_o;
  wire _al_u175_o;
  wire _al_u176_o;
  wire _al_u178_o;
  wire _al_u180_o;
  wire _al_u182_o;
  wire _al_u183_o;
  wire _al_u185_o;
  wire _al_u187_o;
  wire _al_u189_o;
  wire _al_u190_o;
  wire _al_u192_o;
  wire _al_u194_o;
  wire _al_u196_o;
  wire _al_u197_o;
  wire _al_u199_o;
  wire _al_u201_o;
  wire _al_u203_o;
  wire _al_u204_o;
  wire _al_u206_o;
  wire _al_u208_o;
  wire _al_u210_o;
  wire _al_u211_o;
  wire _al_u213_o;
  wire _al_u215_o;
  wire _al_u217_o;
  wire _al_u218_o;
  wire _al_u220_o;
  wire _al_u222_o;
  wire _al_u224_o;
  wire _al_u225_o;
  wire _al_u227_o;
  wire _al_u228_o;
  wire _al_u230_o;
  wire _al_u232_o;
  wire _al_u234_o;
  wire _al_u235_o;
  wire _al_u237_o;
  wire _al_u239_o;
  wire _al_u241_o;
  wire _al_u243_o;
  wire _al_u245_o;
  wire _al_u247_o;
  wire _al_u248_o;
  wire _al_u250_o;
  wire _al_u251_o;
  wire _al_u252_o;
  wire _al_u253_o;
  wire _al_u254_o;
  wire _al_u255_o;
  wire _al_u256_o;
  wire _al_u257_o;
  wire _al_u258_o;
  wire _al_u259_o;
  wire _al_u261_o;
  wire _al_u262_o;
  wire _al_u263_o;
  wire _al_u264_o;
  wire _al_u266_o;
  wire _al_u268_o;
  wire _al_u269_o;
  wire _al_u271_o;
  wire _al_u272_o;
  wire _al_u273_o;
  wire _al_u274_o;
  wire _al_u275_o;
  wire _al_u276_o;
  wire _al_u277_o;
  wire _al_u278_o;
  wire _al_u279_o;
  wire _al_u280_o;
  wire _al_u282_o;
  wire _al_u283_o;
  wire _al_u284_o;
  wire _al_u285_o;
  wire _al_u286_o;
  wire _al_u287_o;
  wire _al_u288_o;
  wire _al_u289_o;
  wire _al_u290_o;
  wire _al_u292_o;
  wire _al_u293_o;
  wire _al_u294_o;
  wire _al_u295_o;
  wire _al_u296_o;
  wire _al_u297_o;
  wire _al_u298_o;
  wire _al_u299_o;
  wire _al_u300_o;
  wire _al_u301_o;
  wire _al_u303_o;
  wire _al_u304_o;
  wire _al_u305_o;
  wire _al_u306_o;
  wire _al_u307_o;
  wire _al_u308_o;
  wire _al_u309_o;
  wire _al_u310_o;
  wire _al_u311_o;
  wire _al_u313_o;
  wire _al_u315_o;
  wire _al_u317_o;
  wire _al_u319_o;
  wire _al_u321_o;
  wire _al_u323_o;
  wire _al_u324_o;
  wire _al_u326_o;
  wire _al_u328_o;
  wire _al_u330_o;
  wire _al_u332_o;
  wire _al_u334_o;
  wire _al_u336_o;
  wire _al_u337_o;
  wire _al_u339_o;
  wire _al_u340_o;
  wire _al_u341_o;
  wire _al_u342_o;
  wire _al_u343_o;
  wire _al_u345_o;
  wire _al_u347_o;
  wire _al_u349_o;
  wire _al_u351_o;
  wire _al_u353_o;
  wire _al_u355_o;
  wire _al_u356_o;
  wire _al_u358_o;
  wire _al_u359_o;
  wire _al_u360_o;
  wire _al_u361_o;
  wire _al_u362_o;
  wire _al_u363_o;
  wire _al_u364_o;
  wire _al_u365_o;
  wire _al_u366_o;
  wire _al_u367_o;
  wire _al_u369_o;
  wire _al_u370_o;
  wire _al_u371_o;
  wire _al_u372_o;
  wire _al_u373_o;
  wire _al_u374_o;
  wire _al_u375_o;
  wire _al_u376_o;
  wire _al_u377_o;
  wire _al_u379_o;
  wire _al_u381_o;
  wire _al_u383_o;
  wire _al_u385_o;
  wire _al_u387_o;
  wire _al_u389_o;
  wire _al_u390_o;
  wire _al_u392_o;
  wire _al_u394_o;
  wire _al_u396_o;
  wire _al_u398_o;
  wire _al_u400_o;
  wire _al_u402_o;
  wire _al_u403_o;
  wire _al_u405_o;
  wire _al_u406_o;
  wire _al_u407_o;
  wire _al_u408_o;
  wire _al_u409_o;
  wire _al_u410_o;
  wire _al_u411_o;
  wire _al_u412_o;
  wire _al_u413_o;
  wire _al_u414_o;
  wire _al_u415_o;
  wire _al_u416_o;
  wire _al_u417_o;
  wire _al_u418_o;
  wire _al_u419_o;
  wire _al_u420_o;
  wire _al_u421_o;
  wire _al_u422_o;
  wire _al_u424_o;
  wire _al_u426_o;
  wire _al_u428_o;
  wire _al_u430_o;
  wire _al_u432_o;
  wire _al_u434_o;
  wire _al_u435_o;
  wire _al_u437_o;
  wire _al_u438_o;
  wire _al_u439_o;
  wire _al_u440_o;
  wire _al_u441_o;
  wire _al_u442_o;
  wire _al_u443_o;
  wire _al_u444_o;
  wire _al_u445_o;
  wire _al_u446_o;
  wire _al_u447_o;
  wire _al_u448_o;
  wire _al_u449_o;
  wire _al_u450_o;
  wire _al_u451_o;
  wire _al_u452_o;
  wire _al_u453_o;
  wire _al_u454_o;
  wire _al_u456_o;
  wire _al_u458_o;
  wire _al_u460_o;
  wire _al_u462_o;
  wire _al_u464_o;
  wire _al_u466_o;
  wire _al_u467_o;
  wire _al_u469_o;
  wire _al_u471_o;
  wire _al_u473_o;
  wire _al_u475_o;
  wire _al_u477_o;
  wire _al_u479_o;
  wire _al_u480_o;
  wire _al_u482_o;
  wire _al_u483_o;
  wire _al_u484_o;
  wire _al_u485_o;
  wire _al_u486_o;
  wire _al_u487_o;
  wire _al_u488_o;
  wire _al_u489_o;
  wire _al_u490_o;
  wire _al_u491_o;
  wire _al_u493_o;
  wire _al_u494_o;
  wire _al_u495_o;
  wire _al_u496_o;
  wire _al_u497_o;
  wire _al_u498_o;
  wire _al_u499_o;
  wire _al_u500_o;
  wire _al_u501_o;
  wire _al_u503_o;
  wire _al_u504_o;
  wire _al_u505_o;
  wire _al_u506_o;
  wire _al_u507_o;
  wire _al_u508_o;
  wire _al_u509_o;
  wire _al_u510_o;
  wire _al_u511_o;
  wire _al_u512_o;
  wire _al_u514_o;
  wire _al_u515_o;
  wire _al_u516_o;
  wire _al_u517_o;
  wire _al_u518_o;
  wire _al_u519_o;
  wire _al_u520_o;
  wire _al_u521_o;
  wire _al_u522_o;
  wire _al_u524_o;
  wire _al_u525_o;
  wire _al_u526_o;
  wire _al_u527_o;
  wire _al_u528_o;
  wire _al_u529_o;
  wire _al_u530_o;
  wire _al_u531_o;
  wire _al_u532_o;
  wire _al_u533_o;
  wire _al_u535_o;
  wire _al_u536_o;
  wire _al_u537_o;
  wire _al_u538_o;
  wire _al_u539_o;
  wire _al_u540_o;
  wire _al_u541_o;
  wire _al_u542_o;
  wire _al_u543_o;
  wire _al_u545_o;
  wire _al_u546_o;
  wire _al_u547_o;
  wire _al_u548_o;
  wire _al_u549_o;
  wire _al_u550_o;
  wire _al_u551_o;
  wire _al_u552_o;
  wire _al_u553_o;
  wire _al_u554_o;
  wire _al_u556_o;
  wire _al_u557_o;
  wire _al_u558_o;
  wire _al_u559_o;
  wire _al_u561_o;
  wire _al_u563_o;
  wire _al_u564_o;
  wire _al_u566_o;
  wire _al_u567_o;
  wire _al_u568_o;
  wire _al_u569_o;
  wire _al_u570_o;
  wire _al_u571_o;
  wire _al_u572_o;
  wire _al_u573_o;
  wire _al_u574_o;
  wire _al_u575_o;
  wire _al_u577_o;
  wire _al_u578_o;
  wire _al_u579_o;
  wire _al_u580_o;
  wire _al_u581_o;
  wire _al_u582_o;
  wire _al_u583_o;
  wire _al_u584_o;
  wire _al_u585_o;
  wire _al_u587_o;
  wire _al_u588_o;
  wire _al_u589_o;
  wire _al_u590_o;
  wire _al_u591_o;
  wire _al_u592_o;
  wire _al_u593_o;
  wire _al_u594_o;
  wire _al_u595_o;
  wire _al_u596_o;
  wire _al_u597_o;
  wire _al_u598_o;
  wire _al_u599_o;
  wire _al_u600_o;
  wire _al_u601_o;
  wire _al_u602_o;
  wire _al_u603_o;
  wire _al_u604_o;
  wire _al_u606_o;
  wire _al_u607_o;
  wire _al_u608_o;
  wire _al_u609_o;
  wire _al_u610_o;
  wire _al_u611_o;
  wire _al_u612_o;
  wire _al_u613_o;
  wire _al_u614_o;
  wire _al_u615_o;
  wire _al_u617_o;
  wire _al_u618_o;
  wire _al_u619_o;
  wire _al_u620_o;
  wire _al_u621_o;
  wire _al_u622_o;
  wire _al_u623_o;
  wire _al_u624_o;
  wire _al_u625_o;
  wire _al_u627_o;
  wire _al_u629_o;
  wire _al_u631_o;
  wire _al_u633_o;
  wire _al_u635_o;
  wire _al_u637_o;
  wire _al_u638_o;
  wire _al_u640_o;
  wire _al_u642_o;
  wire _al_u644_o;
  wire _al_u646_o;
  wire _al_u648_o;
  wire _al_u650_o;
  wire _al_u651_o;
  wire _al_u653_o;
  wire _al_u655_o;
  wire _al_u657_o;
  wire _al_u659_o;
  wire _al_u661_o;
  wire _al_u663_o;
  wire _al_u664_o;
  wire _al_u666_o;
  wire _al_u668_o;
  wire _al_u670_o;
  wire _al_u672_o;
  wire _al_u674_o;
  wire _al_u676_o;
  wire _al_u677_o;
  wire _al_u679_o;
  wire _al_u681_o;
  wire _al_u683_o;
  wire _al_u685_o;
  wire _al_u687_o;
  wire _al_u689_o;
  wire _al_u690_o;
  wire _al_u692_o;
  wire _al_u693_o;
  wire _al_u694_o;
  wire _al_u695_o;
  wire _al_u696_o;
  wire _al_u697_o;
  wire _al_u698_o;
  wire _al_u699_o;
  wire _al_u700_o;
  wire _al_u702_o;
  wire _al_u703_o;
  wire _al_u704_o;
  wire _al_u705_o;
  wire _al_u706_o;
  wire _al_u707_o;
  wire _al_u708_o;
  wire _al_u709_o;
  wire _al_u710_o;
  wire _al_u712_o;
  wire _al_u713_o;
  wire _al_u714_o;
  wire _al_u715_o;
  wire _al_u716_o;
  wire _al_u717_o;
  wire _al_u718_o;
  wire _al_u719_o;
  wire _al_u720_o;
  wire _al_u722_o;
  wire _al_u723_o;
  wire _al_u724_o;
  wire _al_u725_o;
  wire _al_u726_o;
  wire _al_u727_o;
  wire _al_u728_o;
  wire _al_u729_o;
  wire _al_u730_o;
  wire _al_u732_o;
  wire _al_u733_o;
  wire _al_u734_o;
  wire _al_u735_o;
  wire _al_u736_o;
  wire _al_u737_o;
  wire _al_u738_o;
  wire _al_u739_o;
  wire _al_u740_o;
  wire _al_u742_o;
  wire _al_u743_o;
  wire _al_u744_o;
  wire _al_u745_o;
  wire _al_u746_o;
  wire _al_u747_o;
  wire _al_u748_o;
  wire _al_u749_o;
  wire _al_u750_o;
  wire _al_u752_o;
  wire _al_u754_o;
  wire _al_u756_o;
  wire _al_u758_o;
  wire _al_u75_o;
  wire _al_u760_o;
  wire _al_u762_o;
  wire _al_u763_o;
  wire _al_u765_o;
  wire _al_u766_o;
  wire _al_u768_o;
  wire _al_u769_o;
  wire _al_u770_o;
  wire _al_u771_o;
  wire _al_u772_o;
  wire _al_u773_o;
  wire _al_u774_o;
  wire _al_u775_o;
  wire _al_u776_o;
  wire _al_u777_o;
  wire _al_u779_o;
  wire _al_u781_o;
  wire _al_u783_o;
  wire _al_u785_o;
  wire _al_u786_o;
  wire _al_u788_o;
  wire _al_u790_o;
  wire _al_u792_o;
  wire _al_u793_o;
  wire _al_u795_o;
  wire _al_u797_o;
  wire _al_u799_o;
  wire _al_u79_o;
  wire _al_u800_o;
  wire _al_u802_o;
  wire _al_u804_o;
  wire _al_u806_o;
  wire _al_u807_o;
  wire _al_u809_o;
  wire _al_u811_o;
  wire _al_u813_o;
  wire _al_u814_o;
  wire _al_u816_o;
  wire _al_u818_o;
  wire _al_u820_o;
  wire _al_u821_o;
  wire _al_u823_o;
  wire _al_u825_o;
  wire _al_u827_o;
  wire _al_u828_o;
  wire _al_u830_o;
  wire _al_u832_o;
  wire _al_u834_o;
  wire _al_u835_o;
  wire _al_u837_o;
  wire _al_u839_o;
  wire _al_u841_o;
  wire _al_u842_o;
  wire _al_u844_o;
  wire _al_u846_o;
  wire _al_u848_o;
  wire _al_u849_o;
  wire _al_u851_o;
  wire _al_u853_o;
  wire _al_u855_o;
  wire _al_u856_o;
  wire _al_u858_o;
  wire _al_u860_o;
  wire _al_u862_o;
  wire _al_u863_o;
  wire _al_u865_o;
  wire _al_u867_o;
  wire _al_u869_o;
  wire _al_u870_o;
  wire _al_u872_o;
  wire _al_u874_o;
  wire _al_u876_o;
  wire _al_u877_o;
  wire _al_u879_o;
  wire _al_u881_o;
  wire _al_u883_o;
  wire _al_u884_o;
  wire _al_u886_o;
  wire _al_u888_o;
  wire _al_u890_o;
  wire _al_u891_o;
  wire _al_u893_o;
  wire _al_u895_o;
  wire _al_u897_o;
  wire _al_u898_o;
  wire _al_u900_o;
  wire _al_u901_o;
  wire _al_u903_o;
  wire _al_u905_o;
  wire _al_u907_o;
  wire _al_u908_o;
  wire _al_u910_o;
  wire _al_u912_o;
  wire _al_u914_o;
  wire _al_u916_o;
  wire _al_u918_o;
  wire _al_u920_o;
  wire _al_u921_o;
  wire _al_u923_o;
  wire _al_u924_o;
  wire _al_u925_o;
  wire _al_u926_o;
  wire _al_u927_o;
  wire _al_u929_o;
  wire _al_u931_o;
  wire _al_u933_o;
  wire _al_u935_o;
  wire _al_u937_o;
  wire _al_u939_o;
  wire _al_u940_o;
  wire _al_u942_o;
  wire _al_u944_o;
  wire _al_u946_o;
  wire _al_u948_o;
  wire _al_u950_o;
  wire _al_u952_o;
  wire _al_u953_o;
  wire _al_u955_o;
  wire _al_u957_o;
  wire _al_u959_o;
  wire _al_u961_o;
  wire _al_u963_o;
  wire _al_u965_o;
  wire _al_u966_o;
  wire _al_u968_o;
  wire _al_u969_o;
  wire _al_u970_o;
  wire _al_u971_o;
  wire _al_u972_o;
  wire _al_u974_o;
  wire _al_u975_o;
  wire _al_u976_o;
  wire _al_u977_o;
  wire _al_u978_o;
  wire _al_u979_o;
  wire _al_u980_o;
  wire _al_u981_o;
  wire _al_u982_o;
  wire _al_u983_o;
  wire _al_u985_o;
  wire _al_u986_o;
  wire _al_u987_o;
  wire _al_u988_o;
  wire _al_u989_o;
  wire _al_u990_o;
  wire _al_u991_o;
  wire _al_u992_o;
  wire _al_u993_o;
  wire _al_u995_o;
  wire _al_u997_o;
  wire _al_u999_o;
  wire n1;
  wire n10;
  wire n13;
  wire n16;
  wire n19;
  wire n22;
  wire n25;
  wire n28;
  wire n31;
  wire n34;
  wire n37;
  wire n4;
  wire n40;
  wire n43;
  wire n46;
  wire n49;
  wire n52;
  wire n55;
  wire n58;
  wire n61;
  wire n64;
  wire n67;
  wire n7;
  wire n70;
  wire n73;
  wire n76;
  wire n79;
  wire n82;
  wire n85;
  wire n88;
  wire n91;
  wire n94;
  wire n98;

  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*A)"),
    .INIT(32'h20000000))
    _al_u100 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n43));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1000 (
    .a(\mux34_b31/B1_4 ),
    .b(\mux34_b31/B1_5 ),
    .c(_al_u999_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b31/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1001 (
    .a(\rfxs[14] [31]),
    .b(\rfxs[15] [31]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1001_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1002 (
    .a(\rfxs[12] [31]),
    .b(\rfxs[13] [31]),
    .c(_al_u1001_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b31/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1003 (
    .a(\rfxs[8] [31]),
    .b(\rfxs[10] [31]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1003_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1004 (
    .a(\rfxs[11] [31]),
    .b(\rfxs[9] [31]),
    .c(_al_u1003_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b31/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1005 (
    .a(\mux34_b31/B1_1 ),
    .b(\mux34_b31/B1_2 ),
    .c(_al_u806_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1005_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1006 (
    .a(\mux34_b31/B3_1 ),
    .b(_al_u1005_o),
    .c(\mux34_b31/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1006_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1007 (
    .a(n98),
    .b(_al_u1006_o),
    .c(i_rd_wdata[31]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[31]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1008 (
    .a(\rfxs[26] [30]),
    .b(\rfxs[27] [30]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1008_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1009 (
    .a(\rfxs[24] [30]),
    .b(\rfxs[25] [30]),
    .c(_al_u1008_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b30/B1_6 ));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*A)"),
    .INIT(32'h20000000))
    _al_u101 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n40));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1010 (
    .a(\rfxs[30] [30]),
    .b(\rfxs[31] [30]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1010_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1011 (
    .a(\rfxs[28] [30]),
    .b(\rfxs[29] [30]),
    .c(_al_u1010_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b30/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1012 (
    .a(\mux34_b30/B1_6 ),
    .b(\mux34_b30/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1012_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1013 (
    .a(\mux34_b30/B1_4 ),
    .b(\mux34_b30/B1_5 ),
    .c(_al_u1012_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b30/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1014 (
    .a(\rfxs[14] [30]),
    .b(\rfxs[15] [30]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1014_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1015 (
    .a(\rfxs[12] [30]),
    .b(\rfxs[13] [30]),
    .c(_al_u1014_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b30/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1016 (
    .a(\rfxs[8] [30]),
    .b(\rfxs[10] [30]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1016_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1017 (
    .a(\rfxs[11] [30]),
    .b(\rfxs[9] [30]),
    .c(_al_u1016_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b30/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1018 (
    .a(\mux34_b30/B1_1 ),
    .b(\mux34_b30/B1_2 ),
    .c(_al_u813_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1018_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1019 (
    .a(\mux34_b30/B3_1 ),
    .b(_al_u1018_o),
    .c(\mux34_b30/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1019_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*~B*A)"),
    .INIT(32'h00002000))
    _al_u102 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n37));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1020 (
    .a(n98),
    .b(_al_u1019_o),
    .c(i_rd_wdata[30]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[30]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1021 (
    .a(\rfxs[22] [3]),
    .b(\rfxs[23] [3]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1021_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1022 (
    .a(\rfxs[20] [3]),
    .b(\rfxs[21] [3]),
    .c(_al_u1021_o),
    .d(i_rs2idx[1]),
    .o(_al_u1022_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1023 (
    .a(\rfxs[18] [3]),
    .b(\rfxs[19] [3]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1023_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1024 (
    .a(\rfxs[16] [3]),
    .b(\rfxs[17] [3]),
    .c(_al_u1023_o),
    .d(i_rs2idx[1]),
    .o(_al_u1024_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1025 (
    .a(_al_u1022_o),
    .b(_al_u1024_o),
    .c(i_rs2idx[2]),
    .o(_al_u1025_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1026 (
    .a(\rfxs[1] [3]),
    .b(\rfxs[2] [3]),
    .c(\rfxs[3] [3]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1026_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1027 (
    .a(\rfxs[5] [3]),
    .b(\rfxs[6] [3]),
    .c(\rfxs[7] [3]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1027_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u1028 (
    .a(_al_u1026_o),
    .b(_al_u1027_o),
    .c(_al_u776_o),
    .d(\rfxs[4] [3]),
    .e(i_rs2idx[2]),
    .o(_al_u1028_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1029 (
    .a(_al_u1025_o),
    .b(_al_u1028_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1029_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*~B*A)"),
    .INIT(32'h00002000))
    _al_u103 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n34));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1030 (
    .a(\rfxs[8] [3]),
    .b(\rfxs[10] [3]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1030_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1031 (
    .a(\rfxs[11] [3]),
    .b(\rfxs[9] [3]),
    .c(_al_u1030_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b3/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1032 (
    .a(\rfxs[14] [3]),
    .b(\rfxs[15] [3]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1032_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1033 (
    .a(\rfxs[12] [3]),
    .b(\rfxs[13] [3]),
    .c(_al_u1032_o),
    .d(i_rs2idx[1]),
    .o(_al_u1033_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u1034 (
    .a(\mux34_b3/B1_2 ),
    .b(_al_u1033_o),
    .c(i_rs2idx[2]),
    .o(_al_u1034_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1035 (
    .a(\rfxs[26] [3]),
    .b(\rfxs[27] [3]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1035_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1036 (
    .a(\rfxs[24] [3]),
    .b(\rfxs[25] [3]),
    .c(_al_u1035_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b3/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1037 (
    .a(\rfxs[30] [3]),
    .b(\rfxs[31] [3]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1037_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1038 (
    .a(\rfxs[28] [3]),
    .b(\rfxs[29] [3]),
    .c(_al_u1037_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b3/B1_7 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u1039 (
    .a(\mux34_b3/B1_6 ),
    .b(\mux34_b3/B1_7 ),
    .c(i_rs2idx[2]),
    .o(_al_u1039_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*A)"),
    .INIT(32'h00200000))
    _al_u104 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n28));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u1040 (
    .a(_al_u1034_o),
    .b(_al_u1039_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1040_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u1041 (
    .a(n98),
    .b(_al_u1040_o),
    .c(_al_u1029_o),
    .d(i_rd_wdata[3]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[3]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1042 (
    .a(\rfxs[26] [29]),
    .b(\rfxs[27] [29]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1042_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1043 (
    .a(\rfxs[24] [29]),
    .b(\rfxs[25] [29]),
    .c(_al_u1042_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b29/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1044 (
    .a(\rfxs[30] [29]),
    .b(\rfxs[31] [29]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1044_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1045 (
    .a(\rfxs[28] [29]),
    .b(\rfxs[29] [29]),
    .c(_al_u1044_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b29/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1046 (
    .a(\rfxs[18] [29]),
    .b(\rfxs[19] [29]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1046_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1047 (
    .a(\rfxs[16] [29]),
    .b(\rfxs[17] [29]),
    .c(_al_u1046_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b29/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1048 (
    .a(\rfxs[22] [29]),
    .b(\rfxs[23] [29]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1048_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1049 (
    .a(\rfxs[20] [29]),
    .b(\rfxs[21] [29]),
    .c(_al_u1048_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b29/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    _al_u105 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n25));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fca))
    _al_u1050 (
    .a(\mux34_b29/B1_4 ),
    .b(\mux34_b29/B1_5 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1050_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u1051 (
    .a(\mux34_b29/B1_6 ),
    .b(\mux34_b29/B1_7 ),
    .c(_al_u1050_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b29/B3_1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1052 (
    .a(\mux34_b29/B3_1 ),
    .b(i_rs2idx[4]),
    .o(_al_u1052_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1053 (
    .a(\rfxs[8] [29]),
    .b(\rfxs[10] [29]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1053_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1054 (
    .a(\rfxs[11] [29]),
    .b(\rfxs[9] [29]),
    .c(_al_u1053_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b29/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1055 (
    .a(\rfxs[1] [29]),
    .b(\rfxs[2] [29]),
    .c(\rfxs[3] [29]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1055_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h005c))
    _al_u1056 (
    .a(\mux34_b29/B1_2 ),
    .b(_al_u1055_o),
    .c(i_rs2idx[3]),
    .d(i_rs2idx[2]),
    .o(_al_u1056_o));
  AL_MAP_LUT5 #(
    .EQN("(D*(~(A)*B*~(C)*~(E)+A*~(B)*C*~(E)+~(A)*B*C*~(E)+A*B*C*~(E)+A*~(B)*~(C)*E+A*B*~(C)*E+A*~(B)*C*E+A*B*C*E))"),
    .INIT(32'haa00e400))
    _al_u1057 (
    .a(_al_u773_o),
    .b(\rfxs[12] [29]),
    .c(\rfxs[13] [29]),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[1]),
    .o(_al_u1057_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*(~(A)*B*~(C)*~(E)+A*~(B)*C*~(E)+~(A)*B*C*~(E)+A*B*C*~(E)+A*~(B)*~(C)*E+A*B*~(C)*E+A*~(B)*C*E+A*B*C*E))"),
    .INIT(32'h00aa00e4))
    _al_u1058 (
    .a(_al_u772_o),
    .b(\rfxs[4] [29]),
    .c(\rfxs[5] [29]),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[1]),
    .o(_al_u1058_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~A*~(E*~C*~B)))"),
    .INIT(32'h00ab00aa))
    _al_u1059 (
    .a(_al_u1056_o),
    .b(_al_u1057_o),
    .c(_al_u1058_o),
    .d(i_rs2idx[4]),
    .e(i_rs2idx[2]),
    .o(_al_u1059_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    _al_u106 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n22));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u1060 (
    .a(n98),
    .b(_al_u1052_o),
    .c(_al_u1059_o),
    .d(i_rd_wdata[29]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[29]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1061 (
    .a(\rfxs[26] [28]),
    .b(\rfxs[27] [28]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1061_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1062 (
    .a(\rfxs[24] [28]),
    .b(\rfxs[25] [28]),
    .c(_al_u1061_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b28/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1063 (
    .a(\rfxs[30] [28]),
    .b(\rfxs[31] [28]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1063_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1064 (
    .a(\rfxs[28] [28]),
    .b(\rfxs[29] [28]),
    .c(_al_u1063_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b28/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1065 (
    .a(\mux34_b28/B1_6 ),
    .b(\mux34_b28/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1065_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1066 (
    .a(\mux34_b28/B1_4 ),
    .b(\mux34_b28/B1_5 ),
    .c(_al_u1065_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b28/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1067 (
    .a(\rfxs[14] [28]),
    .b(\rfxs[15] [28]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1067_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1068 (
    .a(\rfxs[12] [28]),
    .b(\rfxs[13] [28]),
    .c(_al_u1067_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b28/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1069 (
    .a(\rfxs[8] [28]),
    .b(\rfxs[10] [28]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1069_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*A)"),
    .INIT(32'h00200000))
    _al_u107 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n31));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1070 (
    .a(\rfxs[11] [28]),
    .b(\rfxs[9] [28]),
    .c(_al_u1069_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b28/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1071 (
    .a(\mux34_b28/B1_1 ),
    .b(\mux34_b28/B1_2 ),
    .c(_al_u820_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1071_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1072 (
    .a(\mux34_b28/B3_1 ),
    .b(_al_u1071_o),
    .c(\mux34_b28/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1072_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1073 (
    .a(n98),
    .b(_al_u1072_o),
    .c(i_rd_wdata[28]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[28]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1074 (
    .a(\rfxs[26] [27]),
    .b(\rfxs[27] [27]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1074_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1075 (
    .a(\rfxs[24] [27]),
    .b(\rfxs[25] [27]),
    .c(_al_u1074_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b27/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1076 (
    .a(\rfxs[30] [27]),
    .b(\rfxs[31] [27]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1076_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1077 (
    .a(\rfxs[28] [27]),
    .b(\rfxs[29] [27]),
    .c(_al_u1076_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b27/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1078 (
    .a(\mux34_b27/B1_6 ),
    .b(\mux34_b27/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1078_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1079 (
    .a(\mux34_b27/B1_4 ),
    .b(\mux34_b27/B1_5 ),
    .c(_al_u1078_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b27/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u108 (
    .a(i_rdidx[4]),
    .b(i_rdidx[3]),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u108_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1080 (
    .a(\rfxs[14] [27]),
    .b(\rfxs[15] [27]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1080_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1081 (
    .a(\rfxs[12] [27]),
    .b(\rfxs[13] [27]),
    .c(_al_u1080_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b27/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1082 (
    .a(\rfxs[8] [27]),
    .b(\rfxs[10] [27]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1082_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1083 (
    .a(\rfxs[11] [27]),
    .b(\rfxs[9] [27]),
    .c(_al_u1082_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b27/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1084 (
    .a(\mux34_b27/B1_1 ),
    .b(\mux34_b27/B1_2 ),
    .c(_al_u827_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1084_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1085 (
    .a(\mux34_b27/B3_1 ),
    .b(_al_u1084_o),
    .c(\mux34_b27/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1085_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1086 (
    .a(n98),
    .b(_al_u1085_o),
    .c(i_rd_wdata[27]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[27]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1087 (
    .a(\rfxs[18] [26]),
    .b(\rfxs[19] [26]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1087_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1088 (
    .a(\rfxs[16] [26]),
    .b(\rfxs[17] [26]),
    .c(_al_u1087_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b26/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1089 (
    .a(\rfxs[22] [26]),
    .b(\rfxs[23] [26]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1089_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u109 (
    .a(i_rdidx[1]),
    .b(i_rdidx[0]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u109_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1090 (
    .a(\rfxs[20] [26]),
    .b(\rfxs[21] [26]),
    .c(_al_u1089_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b26/B1_5 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u1091 (
    .a(\mux34_b26/B1_4 ),
    .b(\mux34_b26/B1_5 ),
    .c(i_rs2idx[2]),
    .o(_al_u1091_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1092 (
    .a(\rfxs[1] [26]),
    .b(\rfxs[2] [26]),
    .c(\rfxs[3] [26]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1092_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1093 (
    .a(\rfxs[5] [26]),
    .b(\rfxs[6] [26]),
    .c(\rfxs[7] [26]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1093_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u1094 (
    .a(_al_u1092_o),
    .b(_al_u1093_o),
    .c(_al_u776_o),
    .d(\rfxs[4] [26]),
    .e(i_rs2idx[2]),
    .o(_al_u1094_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1095 (
    .a(_al_u1091_o),
    .b(_al_u1094_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1095_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1096 (
    .a(\rfxs[8] [26]),
    .b(\rfxs[10] [26]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1096_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1097 (
    .a(\rfxs[11] [26]),
    .b(\rfxs[9] [26]),
    .c(_al_u1096_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b26/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1098 (
    .a(\rfxs[14] [26]),
    .b(\rfxs[15] [26]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1098_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1099 (
    .a(\rfxs[12] [26]),
    .b(\rfxs[13] [26]),
    .c(_al_u1098_o),
    .d(i_rs2idx[1]),
    .o(_al_u1099_o));
  AL_MAP_LUT5 #(
    .EQN("(D*B*A*~(E@C))"),
    .INIT(32'h80000800))
    _al_u110 (
    .a(_al_u108_o),
    .b(_al_u109_o),
    .c(i_rdidx[2]),
    .d(i_rdwen),
    .e(i_rs1idx[2]),
    .o(n94));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u1100 (
    .a(\mux34_b26/B1_2 ),
    .b(_al_u1099_o),
    .c(i_rs2idx[2]),
    .o(_al_u1100_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1101 (
    .a(\rfxs[30] [26]),
    .b(\rfxs[31] [26]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1101_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1102 (
    .a(\rfxs[28] [26]),
    .b(\rfxs[29] [26]),
    .c(_al_u1101_o),
    .d(i_rs2idx[1]),
    .o(_al_u1102_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1103 (
    .a(\rfxs[26] [26]),
    .b(\rfxs[27] [26]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1103_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1104 (
    .a(\rfxs[24] [26]),
    .b(\rfxs[25] [26]),
    .c(_al_u1103_o),
    .d(i_rs2idx[1]),
    .o(_al_u1104_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1105 (
    .a(_al_u1102_o),
    .b(_al_u1104_o),
    .c(i_rs2idx[2]),
    .o(_al_u1105_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u1106 (
    .a(_al_u1100_o),
    .b(_al_u1105_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1106_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u1107 (
    .a(n98),
    .b(_al_u1106_o),
    .c(_al_u1095_o),
    .d(i_rd_wdata[26]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[26]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1108 (
    .a(\rfxs[26] [25]),
    .b(\rfxs[27] [25]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1108_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1109 (
    .a(\rfxs[24] [25]),
    .b(\rfxs[25] [25]),
    .c(_al_u1108_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b25/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u111 (
    .a(\rfxs[6] [31]),
    .b(\rfxs[7] [31]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u111_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1110 (
    .a(\rfxs[30] [25]),
    .b(\rfxs[31] [25]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1110_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1111 (
    .a(\rfxs[28] [25]),
    .b(\rfxs[29] [25]),
    .c(_al_u1110_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b25/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1112 (
    .a(\mux34_b25/B1_6 ),
    .b(\mux34_b25/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1112_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1113 (
    .a(\mux34_b25/B1_4 ),
    .b(\mux34_b25/B1_5 ),
    .c(_al_u1112_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b25/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1114 (
    .a(\rfxs[14] [25]),
    .b(\rfxs[15] [25]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1114_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1115 (
    .a(\rfxs[12] [25]),
    .b(\rfxs[13] [25]),
    .c(_al_u1114_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b25/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1116 (
    .a(\rfxs[8] [25]),
    .b(\rfxs[10] [25]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1116_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1117 (
    .a(\rfxs[11] [25]),
    .b(\rfxs[9] [25]),
    .c(_al_u1116_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b25/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1118 (
    .a(\mux34_b25/B1_1 ),
    .b(\mux34_b25/B1_2 ),
    .c(_al_u834_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1118_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1119 (
    .a(\mux34_b25/B3_1 ),
    .b(_al_u1118_o),
    .c(\mux34_b25/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1119_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u112 (
    .a(\rfxs[14] [31]),
    .b(\rfxs[15] [31]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u112_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1120 (
    .a(n98),
    .b(_al_u1119_o),
    .c(i_rd_wdata[25]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[25]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1121 (
    .a(\rfxs[26] [24]),
    .b(\rfxs[27] [24]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1121_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1122 (
    .a(\rfxs[24] [24]),
    .b(\rfxs[25] [24]),
    .c(_al_u1121_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b24/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1123 (
    .a(\rfxs[30] [24]),
    .b(\rfxs[31] [24]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1123_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1124 (
    .a(\rfxs[28] [24]),
    .b(\rfxs[29] [24]),
    .c(_al_u1123_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b24/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1125 (
    .a(\mux34_b24/B1_6 ),
    .b(\mux34_b24/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1125_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1126 (
    .a(\mux34_b24/B1_4 ),
    .b(\mux34_b24/B1_5 ),
    .c(_al_u1125_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b24/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1127 (
    .a(\rfxs[14] [24]),
    .b(\rfxs[15] [24]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1127_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1128 (
    .a(\rfxs[12] [24]),
    .b(\rfxs[13] [24]),
    .c(_al_u1127_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b24/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1129 (
    .a(\rfxs[8] [24]),
    .b(\rfxs[10] [24]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1129_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u113 (
    .a(\rfxs[14] [27]),
    .b(\rfxs[15] [27]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u113_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1130 (
    .a(\rfxs[11] [24]),
    .b(\rfxs[9] [24]),
    .c(_al_u1129_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b24/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1131 (
    .a(\mux34_b24/B1_1 ),
    .b(\mux34_b24/B1_2 ),
    .c(_al_u841_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1131_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1132 (
    .a(\mux34_b24/B3_1 ),
    .b(_al_u1131_o),
    .c(\mux34_b24/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1132_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1133 (
    .a(n98),
    .b(_al_u1132_o),
    .c(i_rd_wdata[24]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[24]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1134 (
    .a(\rfxs[26] [23]),
    .b(\rfxs[27] [23]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1134_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1135 (
    .a(\rfxs[24] [23]),
    .b(\rfxs[25] [23]),
    .c(_al_u1134_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b23/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1136 (
    .a(\rfxs[30] [23]),
    .b(\rfxs[31] [23]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1136_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1137 (
    .a(\rfxs[28] [23]),
    .b(\rfxs[29] [23]),
    .c(_al_u1136_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b23/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1138 (
    .a(\rfxs[18] [23]),
    .b(\rfxs[19] [23]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1138_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1139 (
    .a(\rfxs[16] [23]),
    .b(\rfxs[17] [23]),
    .c(_al_u1138_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b23/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u114 (
    .a(\rfxs[14] [25]),
    .b(\rfxs[15] [25]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u114_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1140 (
    .a(\rfxs[22] [23]),
    .b(\rfxs[23] [23]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1140_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1141 (
    .a(\rfxs[20] [23]),
    .b(\rfxs[21] [23]),
    .c(_al_u1140_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b23/B1_5 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fca))
    _al_u1142 (
    .a(\mux34_b23/B1_4 ),
    .b(\mux34_b23/B1_5 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1142_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u1143 (
    .a(\mux34_b23/B1_6 ),
    .b(\mux34_b23/B1_7 ),
    .c(_al_u1142_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b23/B3_1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u1144 (
    .a(\mux34_b23/B3_1 ),
    .b(i_rs2idx[4]),
    .o(_al_u1144_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1145 (
    .a(\rfxs[8] [23]),
    .b(\rfxs[10] [23]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1145_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1146 (
    .a(\rfxs[11] [23]),
    .b(\rfxs[9] [23]),
    .c(_al_u1145_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b23/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1147 (
    .a(\rfxs[1] [23]),
    .b(\rfxs[2] [23]),
    .c(\rfxs[3] [23]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1147_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h005c))
    _al_u1148 (
    .a(\mux34_b23/B1_2 ),
    .b(_al_u1147_o),
    .c(i_rs2idx[3]),
    .d(i_rs2idx[2]),
    .o(_al_u1148_o));
  AL_MAP_LUT5 #(
    .EQN("(D*(~(A)*B*~(C)*~(E)+A*~(B)*C*~(E)+~(A)*B*C*~(E)+A*B*C*~(E)+A*~(B)*~(C)*E+A*B*~(C)*E+A*~(B)*C*E+A*B*C*E))"),
    .INIT(32'haa00e400))
    _al_u1149 (
    .a(_al_u775_o),
    .b(\rfxs[12] [23]),
    .c(\rfxs[13] [23]),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[1]),
    .o(_al_u1149_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u115 (
    .a(\rfxs[14] [18]),
    .b(\rfxs[15] [18]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u115_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*(~(A)*B*~(C)*~(E)+A*~(B)*C*~(E)+~(A)*B*C*~(E)+A*B*C*~(E)+A*~(B)*~(C)*E+A*B*~(C)*E+A*~(B)*C*E+A*B*C*E))"),
    .INIT(32'h00aa00e4))
    _al_u1150 (
    .a(_al_u774_o),
    .b(\rfxs[4] [23]),
    .c(\rfxs[5] [23]),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[1]),
    .o(_al_u1150_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~A*~(E*~C*~B)))"),
    .INIT(32'h00ab00aa))
    _al_u1151 (
    .a(_al_u1148_o),
    .b(_al_u1149_o),
    .c(_al_u1150_o),
    .d(i_rs2idx[4]),
    .e(i_rs2idx[2]),
    .o(_al_u1151_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u1152 (
    .a(n98),
    .b(_al_u1144_o),
    .c(_al_u1151_o),
    .d(i_rd_wdata[23]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[23]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1153 (
    .a(\rfxs[26] [22]),
    .b(\rfxs[27] [22]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1153_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1154 (
    .a(\rfxs[24] [22]),
    .b(\rfxs[25] [22]),
    .c(_al_u1153_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b22/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1155 (
    .a(\rfxs[30] [22]),
    .b(\rfxs[31] [22]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1155_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1156 (
    .a(\rfxs[28] [22]),
    .b(\rfxs[29] [22]),
    .c(_al_u1155_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b22/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1157 (
    .a(\mux34_b22/B1_6 ),
    .b(\mux34_b22/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1157_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1158 (
    .a(\mux34_b22/B1_4 ),
    .b(\mux34_b22/B1_5 ),
    .c(_al_u1157_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b22/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1159 (
    .a(\rfxs[14] [22]),
    .b(\rfxs[15] [22]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1159_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u116 (
    .a(i_rs1idx[1]),
    .b(i_rs1idx[0]),
    .o(_al_u116_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1160 (
    .a(\rfxs[12] [22]),
    .b(\rfxs[13] [22]),
    .c(_al_u1159_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b22/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1161 (
    .a(\rfxs[8] [22]),
    .b(\rfxs[10] [22]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1161_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1162 (
    .a(\rfxs[11] [22]),
    .b(\rfxs[9] [22]),
    .c(_al_u1161_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b22/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1163 (
    .a(\mux34_b22/B1_1 ),
    .b(\mux34_b22/B1_2 ),
    .c(_al_u848_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1163_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1164 (
    .a(\mux34_b22/B3_1 ),
    .b(_al_u1163_o),
    .c(\mux34_b22/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1164_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1165 (
    .a(n98),
    .b(_al_u1164_o),
    .c(i_rd_wdata[22]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[22]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1166 (
    .a(\rfxs[22] [21]),
    .b(\rfxs[23] [21]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1166_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1167 (
    .a(\rfxs[20] [21]),
    .b(\rfxs[21] [21]),
    .c(_al_u1166_o),
    .d(i_rs2idx[1]),
    .o(_al_u1167_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1168 (
    .a(\rfxs[18] [21]),
    .b(\rfxs[19] [21]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1168_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1169 (
    .a(\rfxs[16] [21]),
    .b(\rfxs[17] [21]),
    .c(_al_u1168_o),
    .d(i_rs2idx[1]),
    .o(_al_u1169_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u117 (
    .a(\rfxs[18] [9]),
    .b(\rfxs[19] [9]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u117_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1170 (
    .a(_al_u1167_o),
    .b(_al_u1169_o),
    .c(i_rs2idx[2]),
    .o(_al_u1170_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1171 (
    .a(\rfxs[1] [21]),
    .b(\rfxs[2] [21]),
    .c(\rfxs[3] [21]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1171_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1172 (
    .a(\rfxs[5] [21]),
    .b(\rfxs[6] [21]),
    .c(\rfxs[7] [21]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1172_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u1173 (
    .a(_al_u1171_o),
    .b(_al_u1172_o),
    .c(_al_u776_o),
    .d(\rfxs[4] [21]),
    .e(i_rs2idx[2]),
    .o(_al_u1173_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1174 (
    .a(_al_u1170_o),
    .b(_al_u1173_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1174_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1175 (
    .a(\rfxs[8] [21]),
    .b(\rfxs[10] [21]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1175_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1176 (
    .a(\rfxs[11] [21]),
    .b(\rfxs[9] [21]),
    .c(_al_u1175_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b21/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1177 (
    .a(\rfxs[14] [21]),
    .b(\rfxs[15] [21]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1177_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1178 (
    .a(\rfxs[12] [21]),
    .b(\rfxs[13] [21]),
    .c(_al_u1177_o),
    .d(i_rs2idx[1]),
    .o(_al_u1178_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u1179 (
    .a(\mux34_b21/B1_2 ),
    .b(_al_u1178_o),
    .c(i_rs2idx[2]),
    .o(_al_u1179_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u118 (
    .a(\rfxs[16] [9]),
    .b(\rfxs[17] [9]),
    .c(_al_u117_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b9/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1180 (
    .a(\rfxs[30] [21]),
    .b(\rfxs[31] [21]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1180_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1181 (
    .a(\rfxs[28] [21]),
    .b(\rfxs[29] [21]),
    .c(_al_u1180_o),
    .d(i_rs2idx[1]),
    .o(_al_u1181_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1182 (
    .a(\rfxs[26] [21]),
    .b(\rfxs[27] [21]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1182_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1183 (
    .a(\rfxs[24] [21]),
    .b(\rfxs[25] [21]),
    .c(_al_u1182_o),
    .d(i_rs2idx[1]),
    .o(_al_u1183_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1184 (
    .a(_al_u1181_o),
    .b(_al_u1183_o),
    .c(i_rs2idx[2]),
    .o(_al_u1184_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u1185 (
    .a(_al_u1179_o),
    .b(_al_u1184_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1185_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u1186 (
    .a(n98),
    .b(_al_u1185_o),
    .c(_al_u1174_o),
    .d(i_rd_wdata[21]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[21]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1187 (
    .a(\rfxs[22] [20]),
    .b(\rfxs[23] [20]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1187_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1188 (
    .a(\rfxs[20] [20]),
    .b(\rfxs[21] [20]),
    .c(_al_u1187_o),
    .d(i_rs2idx[1]),
    .o(_al_u1188_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1189 (
    .a(\rfxs[18] [20]),
    .b(\rfxs[19] [20]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1189_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u119 (
    .a(\rfxs[22] [9]),
    .b(\rfxs[23] [9]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u119_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1190 (
    .a(\rfxs[16] [20]),
    .b(\rfxs[17] [20]),
    .c(_al_u1189_o),
    .d(i_rs2idx[1]),
    .o(_al_u1190_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1191 (
    .a(_al_u1188_o),
    .b(_al_u1190_o),
    .c(i_rs2idx[2]),
    .o(_al_u1191_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1192 (
    .a(\rfxs[1] [20]),
    .b(\rfxs[2] [20]),
    .c(\rfxs[3] [20]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1192_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1193 (
    .a(\rfxs[5] [20]),
    .b(\rfxs[6] [20]),
    .c(\rfxs[7] [20]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1193_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u1194 (
    .a(_al_u1192_o),
    .b(_al_u1193_o),
    .c(_al_u776_o),
    .d(\rfxs[4] [20]),
    .e(i_rs2idx[2]),
    .o(_al_u1194_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1195 (
    .a(_al_u1191_o),
    .b(_al_u1194_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1195_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1196 (
    .a(\rfxs[8] [20]),
    .b(\rfxs[10] [20]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1196_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1197 (
    .a(\rfxs[11] [20]),
    .b(\rfxs[9] [20]),
    .c(_al_u1196_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b20/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1198 (
    .a(\rfxs[14] [20]),
    .b(\rfxs[15] [20]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1198_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1199 (
    .a(\rfxs[12] [20]),
    .b(\rfxs[13] [20]),
    .c(_al_u1198_o),
    .d(i_rs2idx[1]),
    .o(_al_u1199_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u120 (
    .a(\rfxs[20] [9]),
    .b(\rfxs[21] [9]),
    .c(_al_u119_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b9/B1_5 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u1200 (
    .a(\mux34_b20/B1_2 ),
    .b(_al_u1199_o),
    .c(i_rs2idx[2]),
    .o(_al_u1200_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1201 (
    .a(\rfxs[30] [20]),
    .b(\rfxs[31] [20]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1201_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1202 (
    .a(\rfxs[28] [20]),
    .b(\rfxs[29] [20]),
    .c(_al_u1201_o),
    .d(i_rs2idx[1]),
    .o(_al_u1202_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1203 (
    .a(\rfxs[26] [20]),
    .b(\rfxs[27] [20]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1203_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1204 (
    .a(\rfxs[24] [20]),
    .b(\rfxs[25] [20]),
    .c(_al_u1203_o),
    .d(i_rs2idx[1]),
    .o(_al_u1204_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1205 (
    .a(_al_u1202_o),
    .b(_al_u1204_o),
    .c(i_rs2idx[2]),
    .o(_al_u1205_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u1206 (
    .a(_al_u1200_o),
    .b(_al_u1205_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1206_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u1207 (
    .a(n98),
    .b(_al_u1206_o),
    .c(_al_u1195_o),
    .d(i_rd_wdata[20]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[20]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1208 (
    .a(\rfxs[22] [2]),
    .b(\rfxs[23] [2]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1208_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1209 (
    .a(\rfxs[20] [2]),
    .b(\rfxs[21] [2]),
    .c(_al_u1208_o),
    .d(i_rs2idx[1]),
    .o(_al_u1209_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u121 (
    .a(\rfxs[26] [9]),
    .b(\rfxs[27] [9]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u121_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1210 (
    .a(\rfxs[18] [2]),
    .b(\rfxs[19] [2]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1210_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1211 (
    .a(\rfxs[16] [2]),
    .b(\rfxs[17] [2]),
    .c(_al_u1210_o),
    .d(i_rs2idx[1]),
    .o(_al_u1211_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1212 (
    .a(_al_u1209_o),
    .b(_al_u1211_o),
    .c(i_rs2idx[2]),
    .o(_al_u1212_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1213 (
    .a(\rfxs[1] [2]),
    .b(\rfxs[2] [2]),
    .c(\rfxs[3] [2]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1213_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1214 (
    .a(\rfxs[5] [2]),
    .b(\rfxs[6] [2]),
    .c(\rfxs[7] [2]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1214_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u1215 (
    .a(_al_u1213_o),
    .b(_al_u1214_o),
    .c(_al_u776_o),
    .d(\rfxs[4] [2]),
    .e(i_rs2idx[2]),
    .o(_al_u1215_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1216 (
    .a(_al_u1212_o),
    .b(_al_u1215_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1216_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1217 (
    .a(\rfxs[8] [2]),
    .b(\rfxs[10] [2]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1217_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1218 (
    .a(\rfxs[11] [2]),
    .b(\rfxs[9] [2]),
    .c(_al_u1217_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b2/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1219 (
    .a(\rfxs[14] [2]),
    .b(\rfxs[15] [2]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1219_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u122 (
    .a(\rfxs[24] [9]),
    .b(\rfxs[25] [9]),
    .c(_al_u121_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b9/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1220 (
    .a(\rfxs[12] [2]),
    .b(\rfxs[13] [2]),
    .c(_al_u1219_o),
    .d(i_rs2idx[1]),
    .o(_al_u1220_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u1221 (
    .a(\mux34_b2/B1_2 ),
    .b(_al_u1220_o),
    .c(i_rs2idx[2]),
    .o(_al_u1221_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1222 (
    .a(\rfxs[30] [2]),
    .b(\rfxs[31] [2]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1222_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1223 (
    .a(\rfxs[28] [2]),
    .b(\rfxs[29] [2]),
    .c(_al_u1222_o),
    .d(i_rs2idx[1]),
    .o(_al_u1223_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1224 (
    .a(\rfxs[26] [2]),
    .b(\rfxs[27] [2]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1224_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1225 (
    .a(\rfxs[24] [2]),
    .b(\rfxs[25] [2]),
    .c(_al_u1224_o),
    .d(i_rs2idx[1]),
    .o(_al_u1225_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1226 (
    .a(_al_u1223_o),
    .b(_al_u1225_o),
    .c(i_rs2idx[2]),
    .o(_al_u1226_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u1227 (
    .a(_al_u1221_o),
    .b(_al_u1226_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1227_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u1228 (
    .a(n98),
    .b(_al_u1227_o),
    .c(_al_u1216_o),
    .d(i_rd_wdata[2]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[2]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1229 (
    .a(\rfxs[22] [19]),
    .b(\rfxs[23] [19]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1229_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u123 (
    .a(\rfxs[30] [9]),
    .b(\rfxs[31] [9]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u123_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1230 (
    .a(\rfxs[20] [19]),
    .b(\rfxs[21] [19]),
    .c(_al_u1229_o),
    .d(i_rs2idx[1]),
    .o(_al_u1230_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1231 (
    .a(\rfxs[18] [19]),
    .b(\rfxs[19] [19]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1231_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1232 (
    .a(\rfxs[16] [19]),
    .b(\rfxs[17] [19]),
    .c(_al_u1231_o),
    .d(i_rs2idx[1]),
    .o(_al_u1232_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1233 (
    .a(_al_u1230_o),
    .b(_al_u1232_o),
    .c(i_rs2idx[2]),
    .o(_al_u1233_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1234 (
    .a(\rfxs[1] [19]),
    .b(\rfxs[2] [19]),
    .c(\rfxs[3] [19]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1234_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1235 (
    .a(\rfxs[5] [19]),
    .b(\rfxs[6] [19]),
    .c(\rfxs[7] [19]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1235_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u1236 (
    .a(_al_u1234_o),
    .b(_al_u1235_o),
    .c(_al_u776_o),
    .d(\rfxs[4] [19]),
    .e(i_rs2idx[2]),
    .o(_al_u1236_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1237 (
    .a(_al_u1233_o),
    .b(_al_u1236_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1237_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1238 (
    .a(\rfxs[8] [19]),
    .b(\rfxs[10] [19]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1238_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1239 (
    .a(\rfxs[11] [19]),
    .b(\rfxs[9] [19]),
    .c(_al_u1238_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b19/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u124 (
    .a(\rfxs[28] [9]),
    .b(\rfxs[29] [9]),
    .c(_al_u123_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b9/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1240 (
    .a(\rfxs[14] [19]),
    .b(\rfxs[15] [19]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1240_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1241 (
    .a(\rfxs[12] [19]),
    .b(\rfxs[13] [19]),
    .c(_al_u1240_o),
    .d(i_rs2idx[1]),
    .o(_al_u1241_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u1242 (
    .a(\mux34_b19/B1_2 ),
    .b(_al_u1241_o),
    .c(i_rs2idx[2]),
    .o(_al_u1242_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1243 (
    .a(\rfxs[26] [19]),
    .b(\rfxs[27] [19]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1243_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1244 (
    .a(\rfxs[24] [19]),
    .b(\rfxs[25] [19]),
    .c(_al_u1243_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b19/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1245 (
    .a(\rfxs[30] [19]),
    .b(\rfxs[31] [19]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1245_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1246 (
    .a(\rfxs[28] [19]),
    .b(\rfxs[29] [19]),
    .c(_al_u1245_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b19/B1_7 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u1247 (
    .a(\mux34_b19/B1_6 ),
    .b(\mux34_b19/B1_7 ),
    .c(i_rs2idx[2]),
    .o(_al_u1247_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u1248 (
    .a(_al_u1242_o),
    .b(_al_u1247_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1248_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u1249 (
    .a(n98),
    .b(_al_u1248_o),
    .c(_al_u1237_o),
    .d(i_rd_wdata[19]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[19]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u125 (
    .a(i_rs1idx[1]),
    .b(i_rs1idx[0]),
    .o(_al_u125_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1250 (
    .a(\rfxs[26] [18]),
    .b(\rfxs[27] [18]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1250_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1251 (
    .a(\rfxs[24] [18]),
    .b(\rfxs[25] [18]),
    .c(_al_u1250_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b18/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1252 (
    .a(\rfxs[30] [18]),
    .b(\rfxs[31] [18]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1252_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1253 (
    .a(\rfxs[28] [18]),
    .b(\rfxs[29] [18]),
    .c(_al_u1252_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b18/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1254 (
    .a(\mux34_b18/B1_6 ),
    .b(\mux34_b18/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1254_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1255 (
    .a(\mux34_b18/B1_4 ),
    .b(\mux34_b18/B1_5 ),
    .c(_al_u1254_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b18/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1256 (
    .a(\rfxs[14] [18]),
    .b(\rfxs[15] [18]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1256_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1257 (
    .a(\rfxs[12] [18]),
    .b(\rfxs[13] [18]),
    .c(_al_u1256_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b18/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1258 (
    .a(\rfxs[8] [18]),
    .b(\rfxs[10] [18]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1258_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1259 (
    .a(\rfxs[11] [18]),
    .b(\rfxs[9] [18]),
    .c(_al_u1258_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b18/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u126 (
    .a(\rfxs[1] [9]),
    .b(\rfxs[2] [9]),
    .c(\rfxs[3] [9]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u126_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1260 (
    .a(\mux34_b18/B1_1 ),
    .b(\mux34_b18/B1_2 ),
    .c(_al_u855_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1260_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1261 (
    .a(\mux34_b18/B3_1 ),
    .b(_al_u1260_o),
    .c(\mux34_b18/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1261_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1262 (
    .a(n98),
    .b(_al_u1261_o),
    .c(i_rd_wdata[18]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[18]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1263 (
    .a(\rfxs[26] [17]),
    .b(\rfxs[27] [17]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1263_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1264 (
    .a(\rfxs[24] [17]),
    .b(\rfxs[25] [17]),
    .c(_al_u1263_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b17/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1265 (
    .a(\rfxs[30] [17]),
    .b(\rfxs[31] [17]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1265_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1266 (
    .a(\rfxs[28] [17]),
    .b(\rfxs[29] [17]),
    .c(_al_u1265_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b17/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1267 (
    .a(\mux34_b17/B1_6 ),
    .b(\mux34_b17/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1267_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1268 (
    .a(\mux34_b17/B1_4 ),
    .b(\mux34_b17/B1_5 ),
    .c(_al_u1267_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b17/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1269 (
    .a(\rfxs[14] [17]),
    .b(\rfxs[15] [17]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1269_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u127 (
    .a(\rfxs[6] [9]),
    .b(\rfxs[7] [9]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u127_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1270 (
    .a(\rfxs[12] [17]),
    .b(\rfxs[13] [17]),
    .c(_al_u1269_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b17/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1271 (
    .a(\rfxs[8] [17]),
    .b(\rfxs[10] [17]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1271_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1272 (
    .a(\rfxs[11] [17]),
    .b(\rfxs[9] [17]),
    .c(_al_u1271_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b17/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1273 (
    .a(\mux34_b17/B1_1 ),
    .b(\mux34_b17/B1_2 ),
    .c(_al_u862_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1273_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1274 (
    .a(\mux34_b17/B3_1 ),
    .b(_al_u1273_o),
    .c(\mux34_b17/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1274_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1275 (
    .a(n98),
    .b(_al_u1274_o),
    .c(i_rd_wdata[17]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[17]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1276 (
    .a(\rfxs[22] [16]),
    .b(\rfxs[23] [16]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1276_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1277 (
    .a(\rfxs[20] [16]),
    .b(\rfxs[21] [16]),
    .c(_al_u1276_o),
    .d(i_rs2idx[1]),
    .o(_al_u1277_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1278 (
    .a(\rfxs[18] [16]),
    .b(\rfxs[19] [16]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1278_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1279 (
    .a(\rfxs[16] [16]),
    .b(\rfxs[17] [16]),
    .c(_al_u1278_o),
    .d(i_rs2idx[1]),
    .o(_al_u1279_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u128 (
    .a(\rfxs[4] [9]),
    .b(\rfxs[5] [9]),
    .c(_al_u127_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b9/B1_1 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1280 (
    .a(_al_u1277_o),
    .b(_al_u1279_o),
    .c(i_rs2idx[2]),
    .o(_al_u1280_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1281 (
    .a(\rfxs[1] [16]),
    .b(\rfxs[2] [16]),
    .c(\rfxs[3] [16]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1281_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1282 (
    .a(\rfxs[5] [16]),
    .b(\rfxs[6] [16]),
    .c(\rfxs[7] [16]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1282_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u1283 (
    .a(_al_u1281_o),
    .b(_al_u1282_o),
    .c(_al_u776_o),
    .d(\rfxs[4] [16]),
    .e(i_rs2idx[2]),
    .o(_al_u1283_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1284 (
    .a(_al_u1280_o),
    .b(_al_u1283_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1284_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1285 (
    .a(\rfxs[8] [16]),
    .b(\rfxs[10] [16]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1285_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1286 (
    .a(\rfxs[11] [16]),
    .b(\rfxs[9] [16]),
    .c(_al_u1285_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b16/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1287 (
    .a(\rfxs[14] [16]),
    .b(\rfxs[15] [16]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1287_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1288 (
    .a(\rfxs[12] [16]),
    .b(\rfxs[13] [16]),
    .c(_al_u1287_o),
    .d(i_rs2idx[1]),
    .o(_al_u1288_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u1289 (
    .a(\mux34_b16/B1_2 ),
    .b(_al_u1288_o),
    .c(i_rs2idx[2]),
    .o(_al_u1289_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u129 (
    .a(\rfxs[18] [8]),
    .b(\rfxs[19] [8]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u129_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1290 (
    .a(\rfxs[30] [16]),
    .b(\rfxs[31] [16]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1290_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1291 (
    .a(\rfxs[28] [16]),
    .b(\rfxs[29] [16]),
    .c(_al_u1290_o),
    .d(i_rs2idx[1]),
    .o(_al_u1291_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1292 (
    .a(\rfxs[26] [16]),
    .b(\rfxs[27] [16]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1292_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1293 (
    .a(\rfxs[24] [16]),
    .b(\rfxs[25] [16]),
    .c(_al_u1292_o),
    .d(i_rs2idx[1]),
    .o(_al_u1293_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1294 (
    .a(_al_u1291_o),
    .b(_al_u1293_o),
    .c(i_rs2idx[2]),
    .o(_al_u1294_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u1295 (
    .a(_al_u1289_o),
    .b(_al_u1294_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1295_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u1296 (
    .a(n98),
    .b(_al_u1295_o),
    .c(_al_u1284_o),
    .d(i_rd_wdata[16]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[16]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1297 (
    .a(\rfxs[26] [15]),
    .b(\rfxs[27] [15]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1297_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1298 (
    .a(\rfxs[24] [15]),
    .b(\rfxs[25] [15]),
    .c(_al_u1297_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b15/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1299 (
    .a(\rfxs[30] [15]),
    .b(\rfxs[31] [15]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1299_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u130 (
    .a(\rfxs[16] [8]),
    .b(\rfxs[17] [8]),
    .c(_al_u129_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b8/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1300 (
    .a(\rfxs[28] [15]),
    .b(\rfxs[29] [15]),
    .c(_al_u1299_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b15/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1301 (
    .a(\mux34_b15/B1_6 ),
    .b(\mux34_b15/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1301_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1302 (
    .a(\mux34_b15/B1_4 ),
    .b(\mux34_b15/B1_5 ),
    .c(_al_u1301_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b15/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1303 (
    .a(\rfxs[14] [15]),
    .b(\rfxs[15] [15]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1303_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1304 (
    .a(\rfxs[12] [15]),
    .b(\rfxs[13] [15]),
    .c(_al_u1303_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b15/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1305 (
    .a(\rfxs[8] [15]),
    .b(\rfxs[10] [15]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1305_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1306 (
    .a(\rfxs[11] [15]),
    .b(\rfxs[9] [15]),
    .c(_al_u1305_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b15/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1307 (
    .a(\mux34_b15/B1_1 ),
    .b(\mux34_b15/B1_2 ),
    .c(_al_u869_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1307_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1308 (
    .a(\mux34_b15/B3_1 ),
    .b(_al_u1307_o),
    .c(\mux34_b15/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1308_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1309 (
    .a(n98),
    .b(_al_u1308_o),
    .c(i_rd_wdata[15]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[15]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u131 (
    .a(\rfxs[22] [8]),
    .b(\rfxs[23] [8]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u131_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1310 (
    .a(\rfxs[26] [14]),
    .b(\rfxs[27] [14]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1310_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1311 (
    .a(\rfxs[24] [14]),
    .b(\rfxs[25] [14]),
    .c(_al_u1310_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b14/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1312 (
    .a(\rfxs[30] [14]),
    .b(\rfxs[31] [14]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1312_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1313 (
    .a(\rfxs[28] [14]),
    .b(\rfxs[29] [14]),
    .c(_al_u1312_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b14/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1314 (
    .a(\mux34_b14/B1_6 ),
    .b(\mux34_b14/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1314_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1315 (
    .a(\mux34_b14/B1_4 ),
    .b(\mux34_b14/B1_5 ),
    .c(_al_u1314_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b14/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1316 (
    .a(\rfxs[14] [14]),
    .b(\rfxs[15] [14]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1316_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1317 (
    .a(\rfxs[12] [14]),
    .b(\rfxs[13] [14]),
    .c(_al_u1316_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b14/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1318 (
    .a(\rfxs[8] [14]),
    .b(\rfxs[10] [14]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1318_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1319 (
    .a(\rfxs[11] [14]),
    .b(\rfxs[9] [14]),
    .c(_al_u1318_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b14/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u132 (
    .a(\rfxs[20] [8]),
    .b(\rfxs[21] [8]),
    .c(_al_u131_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b8/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1320 (
    .a(\mux34_b14/B1_1 ),
    .b(\mux34_b14/B1_2 ),
    .c(_al_u876_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1320_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1321 (
    .a(\mux34_b14/B3_1 ),
    .b(_al_u1320_o),
    .c(\mux34_b14/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1321_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1322 (
    .a(n98),
    .b(_al_u1321_o),
    .c(i_rd_wdata[14]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[14]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1323 (
    .a(\rfxs[26] [13]),
    .b(\rfxs[27] [13]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1323_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1324 (
    .a(\rfxs[24] [13]),
    .b(\rfxs[25] [13]),
    .c(_al_u1323_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b13/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1325 (
    .a(\rfxs[30] [13]),
    .b(\rfxs[31] [13]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1325_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1326 (
    .a(\rfxs[28] [13]),
    .b(\rfxs[29] [13]),
    .c(_al_u1325_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b13/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1327 (
    .a(\mux34_b13/B1_6 ),
    .b(\mux34_b13/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1327_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1328 (
    .a(\mux34_b13/B1_4 ),
    .b(\mux34_b13/B1_5 ),
    .c(_al_u1327_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b13/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1329 (
    .a(\rfxs[14] [13]),
    .b(\rfxs[15] [13]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1329_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u133 (
    .a(\rfxs[1] [8]),
    .b(\rfxs[2] [8]),
    .c(\rfxs[3] [8]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u133_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1330 (
    .a(\rfxs[12] [13]),
    .b(\rfxs[13] [13]),
    .c(_al_u1329_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b13/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1331 (
    .a(\rfxs[8] [13]),
    .b(\rfxs[10] [13]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1331_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1332 (
    .a(\rfxs[11] [13]),
    .b(\rfxs[9] [13]),
    .c(_al_u1331_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b13/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1333 (
    .a(\mux34_b13/B1_1 ),
    .b(\mux34_b13/B1_2 ),
    .c(_al_u883_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1333_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1334 (
    .a(\mux34_b13/B3_1 ),
    .b(_al_u1333_o),
    .c(\mux34_b13/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1334_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1335 (
    .a(n98),
    .b(_al_u1334_o),
    .c(i_rd_wdata[13]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[13]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1336 (
    .a(\rfxs[26] [12]),
    .b(\rfxs[27] [12]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1336_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1337 (
    .a(\rfxs[24] [12]),
    .b(\rfxs[25] [12]),
    .c(_al_u1336_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b12/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1338 (
    .a(\rfxs[30] [12]),
    .b(\rfxs[31] [12]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1338_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1339 (
    .a(\rfxs[28] [12]),
    .b(\rfxs[29] [12]),
    .c(_al_u1338_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b12/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u134 (
    .a(\rfxs[6] [8]),
    .b(\rfxs[7] [8]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u134_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1340 (
    .a(\mux34_b12/B1_6 ),
    .b(\mux34_b12/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1340_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1341 (
    .a(\mux34_b12/B1_4 ),
    .b(\mux34_b12/B1_5 ),
    .c(_al_u1340_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b12/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1342 (
    .a(\rfxs[14] [12]),
    .b(\rfxs[15] [12]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1342_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1343 (
    .a(\rfxs[12] [12]),
    .b(\rfxs[13] [12]),
    .c(_al_u1342_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b12/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1344 (
    .a(\rfxs[8] [12]),
    .b(\rfxs[10] [12]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1344_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1345 (
    .a(\rfxs[11] [12]),
    .b(\rfxs[9] [12]),
    .c(_al_u1344_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b12/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u1346 (
    .a(\mux34_b12/B1_1 ),
    .b(\mux34_b12/B1_2 ),
    .c(_al_u890_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1346_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u1347 (
    .a(\mux34_b12/B3_1 ),
    .b(_al_u1346_o),
    .c(\mux34_b12/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u1347_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1348 (
    .a(n98),
    .b(_al_u1347_o),
    .c(i_rd_wdata[12]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[12]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1349 (
    .a(\rfxs[18] [11]),
    .b(\rfxs[19] [11]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1349_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u135 (
    .a(\rfxs[4] [8]),
    .b(\rfxs[5] [8]),
    .c(_al_u134_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b8/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1350 (
    .a(\rfxs[16] [11]),
    .b(\rfxs[17] [11]),
    .c(_al_u1349_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b11/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1351 (
    .a(\rfxs[22] [11]),
    .b(\rfxs[23] [11]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1351_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1352 (
    .a(\rfxs[20] [11]),
    .b(\rfxs[21] [11]),
    .c(_al_u1351_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b11/B1_5 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u1353 (
    .a(\mux34_b11/B1_4 ),
    .b(\mux34_b11/B1_5 ),
    .c(i_rs2idx[2]),
    .o(_al_u1353_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1354 (
    .a(\rfxs[1] [11]),
    .b(\rfxs[2] [11]),
    .c(\rfxs[3] [11]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1354_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1355 (
    .a(\rfxs[5] [11]),
    .b(\rfxs[6] [11]),
    .c(\rfxs[7] [11]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1355_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u1356 (
    .a(_al_u1354_o),
    .b(_al_u1355_o),
    .c(_al_u776_o),
    .d(\rfxs[4] [11]),
    .e(i_rs2idx[2]),
    .o(_al_u1356_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1357 (
    .a(_al_u1353_o),
    .b(_al_u1356_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1357_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1358 (
    .a(\rfxs[8] [11]),
    .b(\rfxs[10] [11]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1358_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1359 (
    .a(\rfxs[11] [11]),
    .b(\rfxs[9] [11]),
    .c(_al_u1358_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b11/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u136 (
    .a(\rfxs[18] [4]),
    .b(\rfxs[19] [4]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u136_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1360 (
    .a(\rfxs[14] [11]),
    .b(\rfxs[15] [11]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1360_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1361 (
    .a(\rfxs[12] [11]),
    .b(\rfxs[13] [11]),
    .c(_al_u1360_o),
    .d(i_rs2idx[1]),
    .o(_al_u1361_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u1362 (
    .a(\mux34_b11/B1_2 ),
    .b(_al_u1361_o),
    .c(i_rs2idx[2]),
    .o(_al_u1362_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1363 (
    .a(\rfxs[30] [11]),
    .b(\rfxs[31] [11]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1363_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1364 (
    .a(\rfxs[28] [11]),
    .b(\rfxs[29] [11]),
    .c(_al_u1363_o),
    .d(i_rs2idx[1]),
    .o(_al_u1364_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1365 (
    .a(\rfxs[26] [11]),
    .b(\rfxs[27] [11]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1365_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1366 (
    .a(\rfxs[24] [11]),
    .b(\rfxs[25] [11]),
    .c(_al_u1365_o),
    .d(i_rs2idx[1]),
    .o(_al_u1366_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1367 (
    .a(_al_u1364_o),
    .b(_al_u1366_o),
    .c(i_rs2idx[2]),
    .o(_al_u1367_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u1368 (
    .a(_al_u1362_o),
    .b(_al_u1367_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1368_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u1369 (
    .a(n98),
    .b(_al_u1368_o),
    .c(_al_u1357_o),
    .d(i_rd_wdata[11]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[11]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u137 (
    .a(\rfxs[16] [4]),
    .b(\rfxs[17] [4]),
    .c(_al_u136_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b4/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1370 (
    .a(\rfxs[18] [10]),
    .b(\rfxs[19] [10]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1370_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1371 (
    .a(\rfxs[16] [10]),
    .b(\rfxs[17] [10]),
    .c(_al_u1370_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b10/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1372 (
    .a(\rfxs[22] [10]),
    .b(\rfxs[23] [10]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1372_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1373 (
    .a(\rfxs[20] [10]),
    .b(\rfxs[21] [10]),
    .c(_al_u1372_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b10/B1_5 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u1374 (
    .a(\mux34_b10/B1_4 ),
    .b(\mux34_b10/B1_5 ),
    .c(i_rs2idx[2]),
    .o(_al_u1374_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1375 (
    .a(\rfxs[1] [10]),
    .b(\rfxs[2] [10]),
    .c(\rfxs[3] [10]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1375_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1376 (
    .a(\rfxs[5] [10]),
    .b(\rfxs[6] [10]),
    .c(\rfxs[7] [10]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1376_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u1377 (
    .a(_al_u1375_o),
    .b(_al_u1376_o),
    .c(_al_u776_o),
    .d(\rfxs[4] [10]),
    .e(i_rs2idx[2]),
    .o(_al_u1377_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1378 (
    .a(_al_u1374_o),
    .b(_al_u1377_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1378_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1379 (
    .a(\rfxs[8] [10]),
    .b(\rfxs[10] [10]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1379_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u138 (
    .a(\rfxs[22] [4]),
    .b(\rfxs[23] [4]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u138_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1380 (
    .a(\rfxs[11] [10]),
    .b(\rfxs[9] [10]),
    .c(_al_u1379_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b10/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1381 (
    .a(\rfxs[14] [10]),
    .b(\rfxs[15] [10]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1381_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1382 (
    .a(\rfxs[12] [10]),
    .b(\rfxs[13] [10]),
    .c(_al_u1381_o),
    .d(i_rs2idx[1]),
    .o(_al_u1382_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u1383 (
    .a(\mux34_b10/B1_2 ),
    .b(_al_u1382_o),
    .c(i_rs2idx[2]),
    .o(_al_u1383_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1384 (
    .a(\rfxs[30] [10]),
    .b(\rfxs[31] [10]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1384_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1385 (
    .a(\rfxs[28] [10]),
    .b(\rfxs[29] [10]),
    .c(_al_u1384_o),
    .d(i_rs2idx[1]),
    .o(_al_u1385_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1386 (
    .a(\rfxs[26] [10]),
    .b(\rfxs[27] [10]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1386_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1387 (
    .a(\rfxs[24] [10]),
    .b(\rfxs[25] [10]),
    .c(_al_u1386_o),
    .d(i_rs2idx[1]),
    .o(_al_u1387_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1388 (
    .a(_al_u1385_o),
    .b(_al_u1387_o),
    .c(i_rs2idx[2]),
    .o(_al_u1388_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u1389 (
    .a(_al_u1383_o),
    .b(_al_u1388_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1389_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u139 (
    .a(\rfxs[20] [4]),
    .b(\rfxs[21] [4]),
    .c(_al_u138_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b4/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u1390 (
    .a(n98),
    .b(_al_u1389_o),
    .c(_al_u1378_o),
    .d(i_rd_wdata[10]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[10]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1391 (
    .a(\rfxs[22] [1]),
    .b(\rfxs[23] [1]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1391_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1392 (
    .a(\rfxs[20] [1]),
    .b(\rfxs[21] [1]),
    .c(_al_u1391_o),
    .d(i_rs2idx[1]),
    .o(_al_u1392_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1393 (
    .a(\rfxs[17] [1]),
    .b(\rfxs[18] [1]),
    .c(\rfxs[19] [1]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1393_o));
  AL_MAP_LUT5 #(
    .EQN("((B*~(D*C))*~(A)*~(E)+(B*~(D*C))*A*~(E)+~((B*~(D*C)))*A*E+(B*~(D*C))*A*E)"),
    .INIT(32'haaaa0ccc))
    _al_u1394 (
    .a(_al_u1392_o),
    .b(_al_u1393_o),
    .c(_al_u776_o),
    .d(\rfxs[16] [1]),
    .e(i_rs2idx[2]),
    .o(_al_u1394_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1395 (
    .a(\rfxs[1] [1]),
    .b(\rfxs[2] [1]),
    .c(\rfxs[3] [1]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1395_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u1396 (
    .a(\rfxs[5] [1]),
    .b(\rfxs[6] [1]),
    .c(\rfxs[7] [1]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1396_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u1397 (
    .a(_al_u1395_o),
    .b(_al_u1396_o),
    .c(_al_u776_o),
    .d(\rfxs[4] [1]),
    .e(i_rs2idx[2]),
    .o(_al_u1397_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u1398 (
    .a(_al_u1394_o),
    .b(_al_u1397_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1398_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u1399 (
    .a(\rfxs[8] [1]),
    .b(\rfxs[10] [1]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u1399_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u140 (
    .a(\rfxs[1] [4]),
    .b(\rfxs[2] [4]),
    .c(\rfxs[3] [4]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u140_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1400 (
    .a(\rfxs[11] [1]),
    .b(\rfxs[9] [1]),
    .c(_al_u1399_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b1/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1401 (
    .a(\rfxs[14] [1]),
    .b(\rfxs[15] [1]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1401_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1402 (
    .a(\rfxs[12] [1]),
    .b(\rfxs[13] [1]),
    .c(_al_u1401_o),
    .d(i_rs2idx[1]),
    .o(_al_u1402_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u1403 (
    .a(\mux34_b1/B1_2 ),
    .b(_al_u1402_o),
    .c(i_rs2idx[2]),
    .o(_al_u1403_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1404 (
    .a(\rfxs[30] [1]),
    .b(\rfxs[31] [1]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1404_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1405 (
    .a(\rfxs[28] [1]),
    .b(\rfxs[29] [1]),
    .c(_al_u1404_o),
    .d(i_rs2idx[1]),
    .o(_al_u1405_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1406 (
    .a(\rfxs[26] [1]),
    .b(\rfxs[27] [1]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1406_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u1407 (
    .a(\rfxs[24] [1]),
    .b(\rfxs[25] [1]),
    .c(_al_u1406_o),
    .d(i_rs2idx[1]),
    .o(_al_u1407_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u1408 (
    .a(_al_u1405_o),
    .b(_al_u1407_o),
    .c(i_rs2idx[2]),
    .o(_al_u1408_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u1409 (
    .a(_al_u1403_o),
    .b(_al_u1408_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u1409_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u141 (
    .a(\rfxs[6] [4]),
    .b(\rfxs[7] [4]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u141_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u1410 (
    .a(n98),
    .b(_al_u1409_o),
    .c(_al_u1398_o),
    .d(i_rd_wdata[1]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1411 (
    .a(\rfxs[26] [0]),
    .b(\rfxs[27] [0]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1411_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1412 (
    .a(\rfxs[24] [0]),
    .b(\rfxs[25] [0]),
    .c(_al_u1411_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b0/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1413 (
    .a(\rfxs[30] [0]),
    .b(\rfxs[31] [0]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1413_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1414 (
    .a(\rfxs[28] [0]),
    .b(\rfxs[29] [0]),
    .c(_al_u1413_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b0/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u1415 (
    .a(\mux34_b0/B1_6 ),
    .b(\mux34_b0/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u1415_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u1416 (
    .a(\mux34_b0/B1_4 ),
    .b(\mux34_b0/B1_5 ),
    .c(_al_u1415_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b0/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u1417 (
    .a(\rfxs[14] [0]),
    .b(\rfxs[15] [0]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u1417_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u1418 (
    .a(\rfxs[12] [0]),
    .b(\rfxs[13] [0]),
    .c(_al_u1417_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b0/B1_3 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hccaaff0f))
    _al_u1419 (
    .a(\mux34_b0/B1_1 ),
    .b(\mux34_b0/B1_3 ),
    .c(_al_u897_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u1419_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u142 (
    .a(\rfxs[4] [4]),
    .b(\rfxs[5] [4]),
    .c(_al_u141_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b4/B1_1 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55ff0f33))
    _al_u1420 (
    .a(\rfxs[11] [0]),
    .b(\rfxs[8] [0]),
    .c(\rfxs[10] [0]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u1420_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u1421 (
    .a(\rfxs[9] [0]),
    .b(i_rs2idx[1]),
    .c(i_rs2idx[0]),
    .o(_al_u1421_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u1422 (
    .a(_al_u1420_o),
    .b(_al_u1421_o),
    .c(i_rs2idx[3]),
    .d(i_rs2idx[2]),
    .o(_al_u1422_o));
  AL_MAP_LUT4 #(
    .EQN("~((~C*B)*~(A)*~(D)+(~C*B)*A*~(D)+~((~C*B))*A*D+(~C*B)*A*D)"),
    .INIT(16'h55f3))
    _al_u1423 (
    .a(\mux34_b0/B3_1 ),
    .b(_al_u1419_o),
    .c(_al_u1422_o),
    .d(i_rs2idx[4]),
    .o(_al_u1423_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u1424 (
    .a(n98),
    .b(_al_u1423_o),
    .c(i_rd_wdata[0]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[0]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u143 (
    .a(\rfxs[18] [30]),
    .b(\rfxs[19] [30]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u143_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u144 (
    .a(\rfxs[16] [30]),
    .b(\rfxs[17] [30]),
    .c(_al_u143_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b30/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u145 (
    .a(\rfxs[22] [30]),
    .b(\rfxs[23] [30]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u145_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u146 (
    .a(\rfxs[20] [30]),
    .b(\rfxs[21] [30]),
    .c(_al_u145_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b30/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u147 (
    .a(\rfxs[1] [30]),
    .b(\rfxs[2] [30]),
    .c(\rfxs[3] [30]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u147_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u148 (
    .a(\rfxs[6] [30]),
    .b(\rfxs[7] [30]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u148_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u149 (
    .a(\rfxs[4] [30]),
    .b(\rfxs[5] [30]),
    .c(_al_u148_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b30/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u150 (
    .a(\rfxs[18] [29]),
    .b(\rfxs[19] [29]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u150_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u151 (
    .a(\rfxs[16] [29]),
    .b(\rfxs[17] [29]),
    .c(_al_u150_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b29/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u152 (
    .a(\rfxs[22] [29]),
    .b(\rfxs[23] [29]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u152_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u153 (
    .a(\rfxs[20] [29]),
    .b(\rfxs[21] [29]),
    .c(_al_u152_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b29/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u154 (
    .a(\rfxs[1] [29]),
    .b(\rfxs[2] [29]),
    .c(\rfxs[3] [29]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u154_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u155 (
    .a(\rfxs[6] [29]),
    .b(\rfxs[7] [29]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u155_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u156 (
    .a(\rfxs[4] [29]),
    .b(\rfxs[5] [29]),
    .c(_al_u155_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b29/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u157 (
    .a(\rfxs[18] [28]),
    .b(\rfxs[19] [28]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u157_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u158 (
    .a(\rfxs[16] [28]),
    .b(\rfxs[17] [28]),
    .c(_al_u157_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b28/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u159 (
    .a(\rfxs[22] [28]),
    .b(\rfxs[23] [28]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u159_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u160 (
    .a(\rfxs[20] [28]),
    .b(\rfxs[21] [28]),
    .c(_al_u159_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b28/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u161 (
    .a(\rfxs[1] [28]),
    .b(\rfxs[2] [28]),
    .c(\rfxs[3] [28]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u161_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u162 (
    .a(\rfxs[6] [28]),
    .b(\rfxs[7] [28]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u162_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u163 (
    .a(\rfxs[4] [28]),
    .b(\rfxs[5] [28]),
    .c(_al_u162_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b28/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u164 (
    .a(\rfxs[18] [26]),
    .b(\rfxs[19] [26]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u164_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u165 (
    .a(\rfxs[16] [26]),
    .b(\rfxs[17] [26]),
    .c(_al_u164_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b26/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u166 (
    .a(\rfxs[22] [26]),
    .b(\rfxs[23] [26]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u166_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u167 (
    .a(\rfxs[20] [26]),
    .b(\rfxs[21] [26]),
    .c(_al_u166_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b26/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u168 (
    .a(\rfxs[1] [26]),
    .b(\rfxs[2] [26]),
    .c(\rfxs[3] [26]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u168_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u169 (
    .a(\rfxs[6] [26]),
    .b(\rfxs[7] [26]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u169_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u170 (
    .a(\rfxs[4] [26]),
    .b(\rfxs[5] [26]),
    .c(_al_u169_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b26/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u171 (
    .a(\rfxs[18] [24]),
    .b(\rfxs[19] [24]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u171_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u172 (
    .a(\rfxs[16] [24]),
    .b(\rfxs[17] [24]),
    .c(_al_u171_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b24/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u173 (
    .a(\rfxs[22] [24]),
    .b(\rfxs[23] [24]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u173_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u174 (
    .a(\rfxs[20] [24]),
    .b(\rfxs[21] [24]),
    .c(_al_u173_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b24/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u175 (
    .a(\rfxs[1] [24]),
    .b(\rfxs[2] [24]),
    .c(\rfxs[3] [24]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u175_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u176 (
    .a(\rfxs[6] [24]),
    .b(\rfxs[7] [24]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u176_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u177 (
    .a(\rfxs[4] [24]),
    .b(\rfxs[5] [24]),
    .c(_al_u176_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b24/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u178 (
    .a(\rfxs[18] [23]),
    .b(\rfxs[19] [23]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u178_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u179 (
    .a(\rfxs[16] [23]),
    .b(\rfxs[17] [23]),
    .c(_al_u178_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b23/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u180 (
    .a(\rfxs[22] [23]),
    .b(\rfxs[23] [23]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u180_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u181 (
    .a(\rfxs[20] [23]),
    .b(\rfxs[21] [23]),
    .c(_al_u180_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b23/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u182 (
    .a(\rfxs[1] [23]),
    .b(\rfxs[2] [23]),
    .c(\rfxs[3] [23]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u182_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u183 (
    .a(\rfxs[6] [23]),
    .b(\rfxs[7] [23]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u183_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u184 (
    .a(\rfxs[4] [23]),
    .b(\rfxs[5] [23]),
    .c(_al_u183_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b23/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u185 (
    .a(\rfxs[18] [16]),
    .b(\rfxs[19] [16]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u185_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u186 (
    .a(\rfxs[16] [16]),
    .b(\rfxs[17] [16]),
    .c(_al_u185_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b16/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u187 (
    .a(\rfxs[22] [16]),
    .b(\rfxs[23] [16]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u187_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u188 (
    .a(\rfxs[20] [16]),
    .b(\rfxs[21] [16]),
    .c(_al_u187_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b16/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u189 (
    .a(\rfxs[1] [16]),
    .b(\rfxs[2] [16]),
    .c(\rfxs[3] [16]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u189_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u190 (
    .a(\rfxs[6] [16]),
    .b(\rfxs[7] [16]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u190_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u191 (
    .a(\rfxs[4] [16]),
    .b(\rfxs[5] [16]),
    .c(_al_u190_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b16/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u192 (
    .a(\rfxs[18] [15]),
    .b(\rfxs[19] [15]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u192_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u193 (
    .a(\rfxs[16] [15]),
    .b(\rfxs[17] [15]),
    .c(_al_u192_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b15/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u194 (
    .a(\rfxs[22] [15]),
    .b(\rfxs[23] [15]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u194_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u195 (
    .a(\rfxs[20] [15]),
    .b(\rfxs[21] [15]),
    .c(_al_u194_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b15/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u196 (
    .a(\rfxs[1] [15]),
    .b(\rfxs[2] [15]),
    .c(\rfxs[3] [15]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u196_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u197 (
    .a(\rfxs[6] [15]),
    .b(\rfxs[7] [15]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u197_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u198 (
    .a(\rfxs[4] [15]),
    .b(\rfxs[5] [15]),
    .c(_al_u197_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b15/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u199 (
    .a(\rfxs[18] [14]),
    .b(\rfxs[19] [14]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u199_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u200 (
    .a(\rfxs[16] [14]),
    .b(\rfxs[17] [14]),
    .c(_al_u199_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b14/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u201 (
    .a(\rfxs[22] [14]),
    .b(\rfxs[23] [14]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u201_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u202 (
    .a(\rfxs[20] [14]),
    .b(\rfxs[21] [14]),
    .c(_al_u201_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b14/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u203 (
    .a(\rfxs[1] [14]),
    .b(\rfxs[2] [14]),
    .c(\rfxs[3] [14]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u203_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u204 (
    .a(\rfxs[6] [14]),
    .b(\rfxs[7] [14]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u204_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u205 (
    .a(\rfxs[4] [14]),
    .b(\rfxs[5] [14]),
    .c(_al_u204_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b14/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u206 (
    .a(\rfxs[18] [13]),
    .b(\rfxs[19] [13]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u206_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u207 (
    .a(\rfxs[16] [13]),
    .b(\rfxs[17] [13]),
    .c(_al_u206_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b13/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u208 (
    .a(\rfxs[22] [13]),
    .b(\rfxs[23] [13]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u208_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u209 (
    .a(\rfxs[20] [13]),
    .b(\rfxs[21] [13]),
    .c(_al_u208_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b13/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u210 (
    .a(\rfxs[1] [13]),
    .b(\rfxs[2] [13]),
    .c(\rfxs[3] [13]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u210_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u211 (
    .a(\rfxs[6] [13]),
    .b(\rfxs[7] [13]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u211_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u212 (
    .a(\rfxs[4] [13]),
    .b(\rfxs[5] [13]),
    .c(_al_u211_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b13/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u213 (
    .a(\rfxs[18] [12]),
    .b(\rfxs[19] [12]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u213_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u214 (
    .a(\rfxs[16] [12]),
    .b(\rfxs[17] [12]),
    .c(_al_u213_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b12/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u215 (
    .a(\rfxs[22] [12]),
    .b(\rfxs[23] [12]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u215_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u216 (
    .a(\rfxs[20] [12]),
    .b(\rfxs[21] [12]),
    .c(_al_u215_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b12/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u217 (
    .a(\rfxs[1] [12]),
    .b(\rfxs[2] [12]),
    .c(\rfxs[3] [12]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u217_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u218 (
    .a(\rfxs[6] [12]),
    .b(\rfxs[7] [12]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u218_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u219 (
    .a(\rfxs[4] [12]),
    .b(\rfxs[5] [12]),
    .c(_al_u218_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b12/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u220 (
    .a(\rfxs[18] [0]),
    .b(\rfxs[19] [0]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u220_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u221 (
    .a(\rfxs[16] [0]),
    .b(\rfxs[17] [0]),
    .c(_al_u220_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b0/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u222 (
    .a(\rfxs[22] [0]),
    .b(\rfxs[23] [0]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u222_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u223 (
    .a(\rfxs[20] [0]),
    .b(\rfxs[21] [0]),
    .c(_al_u222_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b0/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u224 (
    .a(\rfxs[1] [0]),
    .b(\rfxs[2] [0]),
    .c(\rfxs[3] [0]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u224_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u225 (
    .a(\rfxs[6] [0]),
    .b(\rfxs[7] [0]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u225_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u226 (
    .a(\rfxs[4] [0]),
    .b(\rfxs[5] [0]),
    .c(_al_u225_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b0/B1_1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u227 (
    .a(i_rs1idx[3]),
    .b(i_rs1idx[2]),
    .o(_al_u227_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u228 (
    .a(\mux31_b9/B1_6 ),
    .b(\mux31_b9/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u228_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u229 (
    .a(\mux31_b9/B1_4 ),
    .b(\mux31_b9/B1_5 ),
    .c(_al_u228_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b9/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u230 (
    .a(\rfxs[14] [9]),
    .b(\rfxs[15] [9]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u230_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u231 (
    .a(\rfxs[12] [9]),
    .b(\rfxs[13] [9]),
    .c(_al_u230_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b9/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u232 (
    .a(\rfxs[8] [9]),
    .b(\rfxs[10] [9]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u232_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u233 (
    .a(\rfxs[11] [9]),
    .b(\rfxs[9] [9]),
    .c(_al_u232_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b9/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u234 (
    .a(\mux31_b9/B1_1 ),
    .b(\mux31_b9/B1_2 ),
    .c(_al_u126_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u234_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u235 (
    .a(\mux31_b9/B3_1 ),
    .b(_al_u234_o),
    .c(\mux31_b9/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u235_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u236 (
    .a(n94),
    .b(_al_u235_o),
    .c(i_rd_wdata[9]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[9]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u237 (
    .a(\rfxs[26] [8]),
    .b(\rfxs[27] [8]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u237_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u238 (
    .a(\rfxs[24] [8]),
    .b(\rfxs[25] [8]),
    .c(_al_u237_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b8/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u239 (
    .a(\rfxs[30] [8]),
    .b(\rfxs[31] [8]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u239_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u240 (
    .a(\rfxs[28] [8]),
    .b(\rfxs[29] [8]),
    .c(_al_u239_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b8/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u241 (
    .a(\mux31_b8/B1_6 ),
    .b(\mux31_b8/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u241_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u242 (
    .a(\mux31_b8/B1_4 ),
    .b(\mux31_b8/B1_5 ),
    .c(_al_u241_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b8/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u243 (
    .a(\rfxs[14] [8]),
    .b(\rfxs[15] [8]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u243_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u244 (
    .a(\rfxs[12] [8]),
    .b(\rfxs[13] [8]),
    .c(_al_u243_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b8/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u245 (
    .a(\rfxs[8] [8]),
    .b(\rfxs[10] [8]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u245_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u246 (
    .a(\rfxs[11] [8]),
    .b(\rfxs[9] [8]),
    .c(_al_u245_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b8/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u247 (
    .a(\mux31_b8/B1_1 ),
    .b(\mux31_b8/B1_2 ),
    .c(_al_u133_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u247_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u248 (
    .a(\mux31_b8/B3_1 ),
    .b(_al_u247_o),
    .c(\mux31_b8/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u248_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u249 (
    .a(n94),
    .b(_al_u248_o),
    .c(i_rd_wdata[8]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[8]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u250 (
    .a(\rfxs[22] [7]),
    .b(\rfxs[23] [7]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u250_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u251 (
    .a(\rfxs[20] [7]),
    .b(\rfxs[21] [7]),
    .c(_al_u250_o),
    .d(i_rs1idx[1]),
    .o(_al_u251_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u252 (
    .a(\rfxs[18] [7]),
    .b(\rfxs[19] [7]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u252_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u253 (
    .a(\rfxs[16] [7]),
    .b(\rfxs[17] [7]),
    .c(_al_u252_o),
    .d(i_rs1idx[1]),
    .o(_al_u253_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u254 (
    .a(_al_u251_o),
    .b(_al_u253_o),
    .c(i_rs1idx[2]),
    .o(_al_u254_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u255 (
    .a(\rfxs[1] [7]),
    .b(\rfxs[2] [7]),
    .c(\rfxs[3] [7]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u255_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u256 (
    .a(\rfxs[5] [7]),
    .b(\rfxs[6] [7]),
    .c(\rfxs[7] [7]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u256_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u257 (
    .a(_al_u255_o),
    .b(_al_u256_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [7]),
    .e(i_rs1idx[2]),
    .o(_al_u257_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u258 (
    .a(_al_u254_o),
    .b(_al_u257_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u258_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u259 (
    .a(\rfxs[8] [7]),
    .b(\rfxs[10] [7]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u259_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u260 (
    .a(\rfxs[11] [7]),
    .b(\rfxs[9] [7]),
    .c(_al_u259_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b7/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u261 (
    .a(\rfxs[14] [7]),
    .b(\rfxs[15] [7]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u261_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u262 (
    .a(\rfxs[12] [7]),
    .b(\rfxs[13] [7]),
    .c(_al_u261_o),
    .d(i_rs1idx[1]),
    .o(_al_u262_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u263 (
    .a(\mux31_b7/B1_2 ),
    .b(_al_u262_o),
    .c(i_rs1idx[2]),
    .o(_al_u263_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u264 (
    .a(\rfxs[26] [7]),
    .b(\rfxs[27] [7]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u264_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u265 (
    .a(\rfxs[24] [7]),
    .b(\rfxs[25] [7]),
    .c(_al_u264_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b7/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u266 (
    .a(\rfxs[30] [7]),
    .b(\rfxs[31] [7]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u266_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u267 (
    .a(\rfxs[28] [7]),
    .b(\rfxs[29] [7]),
    .c(_al_u266_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b7/B1_7 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u268 (
    .a(\mux31_b7/B1_6 ),
    .b(\mux31_b7/B1_7 ),
    .c(i_rs1idx[2]),
    .o(_al_u268_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u269 (
    .a(_al_u263_o),
    .b(_al_u268_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u269_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u270 (
    .a(n94),
    .b(_al_u269_o),
    .c(_al_u258_o),
    .d(i_rd_wdata[7]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[7]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u271 (
    .a(\rfxs[22] [6]),
    .b(\rfxs[23] [6]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u271_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u272 (
    .a(\rfxs[20] [6]),
    .b(\rfxs[21] [6]),
    .c(_al_u271_o),
    .d(i_rs1idx[1]),
    .o(_al_u272_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u273 (
    .a(\rfxs[18] [6]),
    .b(\rfxs[19] [6]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u273_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u274 (
    .a(\rfxs[16] [6]),
    .b(\rfxs[17] [6]),
    .c(_al_u273_o),
    .d(i_rs1idx[1]),
    .o(_al_u274_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u275 (
    .a(_al_u272_o),
    .b(_al_u274_o),
    .c(i_rs1idx[2]),
    .o(_al_u275_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u276 (
    .a(\rfxs[1] [6]),
    .b(\rfxs[2] [6]),
    .c(\rfxs[3] [6]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u276_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u277 (
    .a(\rfxs[5] [6]),
    .b(\rfxs[6] [6]),
    .c(\rfxs[7] [6]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u277_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u278 (
    .a(_al_u276_o),
    .b(_al_u277_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [6]),
    .e(i_rs1idx[2]),
    .o(_al_u278_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u279 (
    .a(_al_u275_o),
    .b(_al_u278_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u279_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u280 (
    .a(\rfxs[8] [6]),
    .b(\rfxs[10] [6]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u280_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u281 (
    .a(\rfxs[11] [6]),
    .b(\rfxs[9] [6]),
    .c(_al_u280_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b6/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u282 (
    .a(\rfxs[14] [6]),
    .b(\rfxs[15] [6]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u282_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u283 (
    .a(\rfxs[12] [6]),
    .b(\rfxs[13] [6]),
    .c(_al_u282_o),
    .d(i_rs1idx[1]),
    .o(_al_u283_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u284 (
    .a(\mux31_b6/B1_2 ),
    .b(_al_u283_o),
    .c(i_rs1idx[2]),
    .o(_al_u284_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u285 (
    .a(\rfxs[30] [6]),
    .b(\rfxs[31] [6]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u285_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u286 (
    .a(\rfxs[28] [6]),
    .b(\rfxs[29] [6]),
    .c(_al_u285_o),
    .d(i_rs1idx[1]),
    .o(_al_u286_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u287 (
    .a(\rfxs[26] [6]),
    .b(\rfxs[27] [6]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u287_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u288 (
    .a(\rfxs[24] [6]),
    .b(\rfxs[25] [6]),
    .c(_al_u287_o),
    .d(i_rs1idx[1]),
    .o(_al_u288_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u289 (
    .a(_al_u286_o),
    .b(_al_u288_o),
    .c(i_rs1idx[2]),
    .o(_al_u289_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u290 (
    .a(_al_u284_o),
    .b(_al_u289_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u290_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u291 (
    .a(n94),
    .b(_al_u290_o),
    .c(_al_u279_o),
    .d(i_rd_wdata[6]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[6]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u292 (
    .a(\rfxs[22] [5]),
    .b(\rfxs[23] [5]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u292_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u293 (
    .a(\rfxs[20] [5]),
    .b(\rfxs[21] [5]),
    .c(_al_u292_o),
    .d(i_rs1idx[1]),
    .o(_al_u293_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u294 (
    .a(\rfxs[18] [5]),
    .b(\rfxs[19] [5]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u294_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u295 (
    .a(\rfxs[16] [5]),
    .b(\rfxs[17] [5]),
    .c(_al_u294_o),
    .d(i_rs1idx[1]),
    .o(_al_u295_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u296 (
    .a(_al_u293_o),
    .b(_al_u295_o),
    .c(i_rs1idx[2]),
    .o(_al_u296_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u297 (
    .a(\rfxs[1] [5]),
    .b(\rfxs[2] [5]),
    .c(\rfxs[3] [5]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u297_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u298 (
    .a(\rfxs[5] [5]),
    .b(\rfxs[6] [5]),
    .c(\rfxs[7] [5]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u298_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u299 (
    .a(_al_u297_o),
    .b(_al_u298_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [5]),
    .e(i_rs1idx[2]),
    .o(_al_u299_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u300 (
    .a(_al_u296_o),
    .b(_al_u299_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u300_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u301 (
    .a(\rfxs[8] [5]),
    .b(\rfxs[10] [5]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u301_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u302 (
    .a(\rfxs[11] [5]),
    .b(\rfxs[9] [5]),
    .c(_al_u301_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b5/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u303 (
    .a(\rfxs[14] [5]),
    .b(\rfxs[15] [5]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u303_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u304 (
    .a(\rfxs[12] [5]),
    .b(\rfxs[13] [5]),
    .c(_al_u303_o),
    .d(i_rs1idx[1]),
    .o(_al_u304_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u305 (
    .a(\mux31_b5/B1_2 ),
    .b(_al_u304_o),
    .c(i_rs1idx[2]),
    .o(_al_u305_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u306 (
    .a(\rfxs[30] [5]),
    .b(\rfxs[31] [5]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u306_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u307 (
    .a(\rfxs[28] [5]),
    .b(\rfxs[29] [5]),
    .c(_al_u306_o),
    .d(i_rs1idx[1]),
    .o(_al_u307_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u308 (
    .a(\rfxs[26] [5]),
    .b(\rfxs[27] [5]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u308_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u309 (
    .a(\rfxs[24] [5]),
    .b(\rfxs[25] [5]),
    .c(_al_u308_o),
    .d(i_rs1idx[1]),
    .o(_al_u309_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u310 (
    .a(_al_u307_o),
    .b(_al_u309_o),
    .c(i_rs1idx[2]),
    .o(_al_u310_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u311 (
    .a(_al_u305_o),
    .b(_al_u310_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u311_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u312 (
    .a(n94),
    .b(_al_u311_o),
    .c(_al_u300_o),
    .d(i_rd_wdata[5]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[5]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u313 (
    .a(\rfxs[26] [4]),
    .b(\rfxs[27] [4]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u313_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u314 (
    .a(\rfxs[24] [4]),
    .b(\rfxs[25] [4]),
    .c(_al_u313_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b4/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u315 (
    .a(\rfxs[30] [4]),
    .b(\rfxs[31] [4]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u315_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u316 (
    .a(\rfxs[28] [4]),
    .b(\rfxs[29] [4]),
    .c(_al_u315_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b4/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u317 (
    .a(\mux31_b4/B1_6 ),
    .b(\mux31_b4/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u317_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u318 (
    .a(\mux31_b4/B1_4 ),
    .b(\mux31_b4/B1_5 ),
    .c(_al_u317_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b4/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u319 (
    .a(\rfxs[14] [4]),
    .b(\rfxs[15] [4]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u319_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u320 (
    .a(\rfxs[12] [4]),
    .b(\rfxs[13] [4]),
    .c(_al_u319_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b4/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u321 (
    .a(\rfxs[8] [4]),
    .b(\rfxs[10] [4]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u321_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u322 (
    .a(\rfxs[11] [4]),
    .b(\rfxs[9] [4]),
    .c(_al_u321_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b4/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u323 (
    .a(\mux31_b4/B1_1 ),
    .b(\mux31_b4/B1_2 ),
    .c(_al_u140_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u323_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u324 (
    .a(\mux31_b4/B3_1 ),
    .b(_al_u323_o),
    .c(\mux31_b4/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u324_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u325 (
    .a(n94),
    .b(_al_u324_o),
    .c(i_rd_wdata[4]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[4]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u326 (
    .a(\rfxs[26] [31]),
    .b(\rfxs[27] [31]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u326_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u327 (
    .a(\rfxs[24] [31]),
    .b(\rfxs[25] [31]),
    .c(_al_u326_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b31/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u328 (
    .a(\rfxs[30] [31]),
    .b(\rfxs[31] [31]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u328_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u329 (
    .a(\rfxs[28] [31]),
    .b(\rfxs[29] [31]),
    .c(_al_u328_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b31/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u330 (
    .a(\rfxs[18] [31]),
    .b(\rfxs[19] [31]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u330_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u331 (
    .a(\rfxs[16] [31]),
    .b(\rfxs[17] [31]),
    .c(_al_u330_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b31/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u332 (
    .a(\rfxs[22] [31]),
    .b(\rfxs[23] [31]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u332_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u333 (
    .a(\rfxs[20] [31]),
    .b(\rfxs[21] [31]),
    .c(_al_u332_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b31/B1_5 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fca))
    _al_u334 (
    .a(\mux31_b31/B1_4 ),
    .b(\mux31_b31/B1_5 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u334_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u335 (
    .a(\mux31_b31/B1_6 ),
    .b(\mux31_b31/B1_7 ),
    .c(_al_u334_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b31/B3_1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u336 (
    .a(\mux31_b31/B3_1 ),
    .b(i_rs1idx[4]),
    .o(_al_u336_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u337 (
    .a(\rfxs[8] [31]),
    .b(\rfxs[10] [31]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u337_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u338 (
    .a(\rfxs[11] [31]),
    .b(\rfxs[9] [31]),
    .c(_al_u337_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b31/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u339 (
    .a(\rfxs[1] [31]),
    .b(\rfxs[2] [31]),
    .c(\rfxs[3] [31]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u339_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h005c))
    _al_u340 (
    .a(\mux31_b31/B1_2 ),
    .b(_al_u339_o),
    .c(i_rs1idx[3]),
    .d(i_rs1idx[2]),
    .o(_al_u340_o));
  AL_MAP_LUT5 #(
    .EQN("(D*(~(A)*B*~(C)*~(E)+A*~(B)*C*~(E)+~(A)*B*C*~(E)+A*B*C*~(E)+A*~(B)*~(C)*E+A*B*~(C)*E+A*~(B)*C*E+A*B*C*E))"),
    .INIT(32'haa00e400))
    _al_u341 (
    .a(_al_u112_o),
    .b(\rfxs[12] [31]),
    .c(\rfxs[13] [31]),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[1]),
    .o(_al_u341_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*(~(A)*B*~(C)*~(E)+A*~(B)*C*~(E)+~(A)*B*C*~(E)+A*B*C*~(E)+A*~(B)*~(C)*E+A*B*~(C)*E+A*~(B)*C*E+A*B*C*E))"),
    .INIT(32'h00aa00e4))
    _al_u342 (
    .a(_al_u111_o),
    .b(\rfxs[4] [31]),
    .c(\rfxs[5] [31]),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[1]),
    .o(_al_u342_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~A*~(E*~C*~B)))"),
    .INIT(32'h00ab00aa))
    _al_u343 (
    .a(_al_u340_o),
    .b(_al_u341_o),
    .c(_al_u342_o),
    .d(i_rs1idx[4]),
    .e(i_rs1idx[2]),
    .o(_al_u343_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u344 (
    .a(n94),
    .b(_al_u336_o),
    .c(_al_u343_o),
    .d(i_rd_wdata[31]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[31]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u345 (
    .a(\rfxs[26] [30]),
    .b(\rfxs[27] [30]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u345_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u346 (
    .a(\rfxs[24] [30]),
    .b(\rfxs[25] [30]),
    .c(_al_u345_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b30/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u347 (
    .a(\rfxs[30] [30]),
    .b(\rfxs[31] [30]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u347_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u348 (
    .a(\rfxs[28] [30]),
    .b(\rfxs[29] [30]),
    .c(_al_u347_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b30/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u349 (
    .a(\mux31_b30/B1_6 ),
    .b(\mux31_b30/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u349_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u350 (
    .a(\mux31_b30/B1_4 ),
    .b(\mux31_b30/B1_5 ),
    .c(_al_u349_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b30/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u351 (
    .a(\rfxs[14] [30]),
    .b(\rfxs[15] [30]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u351_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u352 (
    .a(\rfxs[12] [30]),
    .b(\rfxs[13] [30]),
    .c(_al_u351_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b30/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u353 (
    .a(\rfxs[8] [30]),
    .b(\rfxs[10] [30]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u353_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u354 (
    .a(\rfxs[11] [30]),
    .b(\rfxs[9] [30]),
    .c(_al_u353_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b30/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u355 (
    .a(\mux31_b30/B1_1 ),
    .b(\mux31_b30/B1_2 ),
    .c(_al_u147_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u355_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u356 (
    .a(\mux31_b30/B3_1 ),
    .b(_al_u355_o),
    .c(\mux31_b30/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u356_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u357 (
    .a(n94),
    .b(_al_u356_o),
    .c(i_rd_wdata[30]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[30]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u358 (
    .a(\rfxs[22] [3]),
    .b(\rfxs[23] [3]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u358_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u359 (
    .a(\rfxs[20] [3]),
    .b(\rfxs[21] [3]),
    .c(_al_u358_o),
    .d(i_rs1idx[1]),
    .o(_al_u359_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u360 (
    .a(\rfxs[18] [3]),
    .b(\rfxs[19] [3]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u360_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u361 (
    .a(\rfxs[16] [3]),
    .b(\rfxs[17] [3]),
    .c(_al_u360_o),
    .d(i_rs1idx[1]),
    .o(_al_u361_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u362 (
    .a(_al_u359_o),
    .b(_al_u361_o),
    .c(i_rs1idx[2]),
    .o(_al_u362_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u363 (
    .a(\rfxs[1] [3]),
    .b(\rfxs[2] [3]),
    .c(\rfxs[3] [3]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u363_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u364 (
    .a(\rfxs[5] [3]),
    .b(\rfxs[6] [3]),
    .c(\rfxs[7] [3]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u364_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u365 (
    .a(_al_u363_o),
    .b(_al_u364_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [3]),
    .e(i_rs1idx[2]),
    .o(_al_u365_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u366 (
    .a(_al_u362_o),
    .b(_al_u365_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u366_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u367 (
    .a(\rfxs[8] [3]),
    .b(\rfxs[10] [3]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u367_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u368 (
    .a(\rfxs[11] [3]),
    .b(\rfxs[9] [3]),
    .c(_al_u367_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b3/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u369 (
    .a(\rfxs[14] [3]),
    .b(\rfxs[15] [3]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u369_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u370 (
    .a(\rfxs[12] [3]),
    .b(\rfxs[13] [3]),
    .c(_al_u369_o),
    .d(i_rs1idx[1]),
    .o(_al_u370_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u371 (
    .a(\mux31_b3/B1_2 ),
    .b(_al_u370_o),
    .c(i_rs1idx[2]),
    .o(_al_u371_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u372 (
    .a(\rfxs[30] [3]),
    .b(\rfxs[31] [3]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u372_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u373 (
    .a(\rfxs[28] [3]),
    .b(\rfxs[29] [3]),
    .c(_al_u372_o),
    .d(i_rs1idx[1]),
    .o(_al_u373_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u374 (
    .a(\rfxs[26] [3]),
    .b(\rfxs[27] [3]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u374_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u375 (
    .a(\rfxs[24] [3]),
    .b(\rfxs[25] [3]),
    .c(_al_u374_o),
    .d(i_rs1idx[1]),
    .o(_al_u375_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u376 (
    .a(_al_u373_o),
    .b(_al_u375_o),
    .c(i_rs1idx[2]),
    .o(_al_u376_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u377 (
    .a(_al_u371_o),
    .b(_al_u376_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u377_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u378 (
    .a(n94),
    .b(_al_u377_o),
    .c(_al_u366_o),
    .d(i_rd_wdata[3]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[3]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u379 (
    .a(\rfxs[26] [29]),
    .b(\rfxs[27] [29]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u379_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u380 (
    .a(\rfxs[24] [29]),
    .b(\rfxs[25] [29]),
    .c(_al_u379_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b29/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u381 (
    .a(\rfxs[30] [29]),
    .b(\rfxs[31] [29]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u381_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u382 (
    .a(\rfxs[28] [29]),
    .b(\rfxs[29] [29]),
    .c(_al_u381_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b29/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u383 (
    .a(\mux31_b29/B1_6 ),
    .b(\mux31_b29/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u383_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u384 (
    .a(\mux31_b29/B1_4 ),
    .b(\mux31_b29/B1_5 ),
    .c(_al_u383_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b29/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u385 (
    .a(\rfxs[14] [29]),
    .b(\rfxs[15] [29]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u385_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u386 (
    .a(\rfxs[12] [29]),
    .b(\rfxs[13] [29]),
    .c(_al_u385_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b29/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u387 (
    .a(\rfxs[8] [29]),
    .b(\rfxs[10] [29]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u387_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u388 (
    .a(\rfxs[11] [29]),
    .b(\rfxs[9] [29]),
    .c(_al_u387_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b29/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u389 (
    .a(\mux31_b29/B1_1 ),
    .b(\mux31_b29/B1_2 ),
    .c(_al_u154_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u389_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u390 (
    .a(\mux31_b29/B3_1 ),
    .b(_al_u389_o),
    .c(\mux31_b29/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u390_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u391 (
    .a(n94),
    .b(_al_u390_o),
    .c(i_rd_wdata[29]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[29]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u392 (
    .a(\rfxs[26] [28]),
    .b(\rfxs[27] [28]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u392_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u393 (
    .a(\rfxs[24] [28]),
    .b(\rfxs[25] [28]),
    .c(_al_u392_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b28/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u394 (
    .a(\rfxs[30] [28]),
    .b(\rfxs[31] [28]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u394_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u395 (
    .a(\rfxs[28] [28]),
    .b(\rfxs[29] [28]),
    .c(_al_u394_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b28/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u396 (
    .a(\mux31_b28/B1_6 ),
    .b(\mux31_b28/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u396_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u397 (
    .a(\mux31_b28/B1_4 ),
    .b(\mux31_b28/B1_5 ),
    .c(_al_u396_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b28/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u398 (
    .a(\rfxs[14] [28]),
    .b(\rfxs[15] [28]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u398_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u399 (
    .a(\rfxs[12] [28]),
    .b(\rfxs[13] [28]),
    .c(_al_u398_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b28/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u400 (
    .a(\rfxs[8] [28]),
    .b(\rfxs[10] [28]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u400_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u401 (
    .a(\rfxs[11] [28]),
    .b(\rfxs[9] [28]),
    .c(_al_u400_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b28/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u402 (
    .a(\mux31_b28/B1_1 ),
    .b(\mux31_b28/B1_2 ),
    .c(_al_u161_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u402_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u403 (
    .a(\mux31_b28/B3_1 ),
    .b(_al_u402_o),
    .c(\mux31_b28/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u403_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u404 (
    .a(n94),
    .b(_al_u403_o),
    .c(i_rd_wdata[28]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[28]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u405 (
    .a(\rfxs[22] [27]),
    .b(\rfxs[23] [27]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u405_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u406 (
    .a(\rfxs[20] [27]),
    .b(\rfxs[21] [27]),
    .c(_al_u405_o),
    .d(i_rs1idx[1]),
    .o(_al_u406_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u407 (
    .a(\rfxs[18] [27]),
    .b(\rfxs[19] [27]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u407_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u408 (
    .a(\rfxs[16] [27]),
    .b(\rfxs[17] [27]),
    .c(_al_u407_o),
    .d(i_rs1idx[1]),
    .o(_al_u408_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u409 (
    .a(\rfxs[1] [27]),
    .b(\rfxs[2] [27]),
    .c(\rfxs[3] [27]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u409_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u410 (
    .a(\rfxs[6] [27]),
    .b(\rfxs[7] [27]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u410_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u411 (
    .a(\rfxs[4] [27]),
    .b(\rfxs[5] [27]),
    .c(_al_u410_o),
    .d(i_rs1idx[1]),
    .o(_al_u411_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f53))
    _al_u412 (
    .a(_al_u411_o),
    .b(_al_u409_o),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[4]),
    .o(_al_u412_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u413 (
    .a(_al_u406_o),
    .b(_al_u408_o),
    .c(_al_u412_o),
    .d(i_rs1idx[4]),
    .o(_al_u413_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55ff0f33))
    _al_u414 (
    .a(\rfxs[11] [27]),
    .b(\rfxs[8] [27]),
    .c(\rfxs[10] [27]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u414_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(C*B))"),
    .INIT(16'h002a))
    _al_u415 (
    .a(_al_u414_o),
    .b(_al_u125_o),
    .c(\rfxs[9] [27]),
    .d(i_rs1idx[2]),
    .o(_al_u415_o));
  AL_MAP_LUT5 #(
    .EQN("(D*(~(A)*~(B)*~(C)*~(E)+A*~(B)*~(C)*~(E)+A*B*~(C)*~(E)+~(A)*~(B)*C*~(E)+~(A)*~(B)*~(C)*E+~(A)*B*~(C)*E+~(A)*~(B)*C*E+~(A)*B*C*E))"),
    .INIT(32'h55001b00))
    _al_u416 (
    .a(_al_u113_o),
    .b(\rfxs[12] [27]),
    .c(\rfxs[13] [27]),
    .d(i_rs1idx[2]),
    .e(i_rs1idx[1]),
    .o(_al_u416_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u417 (
    .a(\rfxs[29] [27]),
    .b(\rfxs[30] [27]),
    .c(\rfxs[31] [27]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u417_o));
  AL_MAP_LUT4 #(
    .EQN("(D*A*~(C*B))"),
    .INIT(16'h2a00))
    _al_u418 (
    .a(_al_u417_o),
    .b(_al_u116_o),
    .c(\rfxs[28] [27]),
    .d(i_rs1idx[2]),
    .o(_al_u418_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u419 (
    .a(\rfxs[25] [27]),
    .b(\rfxs[26] [27]),
    .c(\rfxs[27] [27]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u419_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(C*B))"),
    .INIT(16'h002a))
    _al_u420 (
    .a(_al_u419_o),
    .b(_al_u116_o),
    .c(\rfxs[24] [27]),
    .d(i_rs1idx[2]),
    .o(_al_u420_o));
  AL_MAP_LUT5 #(
    .EQN("~((~D*~A)*~((~C*~B))*~(E)+(~D*~A)*(~C*~B)*~(E)+~((~D*~A))*(~C*~B)*E+(~D*~A)*(~C*~B)*E)"),
    .INIT(32'hfcfcffaa))
    _al_u421 (
    .a(_al_u415_o),
    .b(_al_u418_o),
    .c(_al_u420_o),
    .d(_al_u416_o),
    .e(i_rs1idx[4]),
    .o(_al_u421_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u422 (
    .a(_al_u413_o),
    .b(_al_u421_o),
    .c(i_rs1idx[3]),
    .o(_al_u422_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u423 (
    .a(n94),
    .b(_al_u422_o),
    .c(i_rd_wdata[27]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[27]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u424 (
    .a(\rfxs[26] [26]),
    .b(\rfxs[27] [26]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u424_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u425 (
    .a(\rfxs[24] [26]),
    .b(\rfxs[25] [26]),
    .c(_al_u424_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b26/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u426 (
    .a(\rfxs[30] [26]),
    .b(\rfxs[31] [26]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u426_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u427 (
    .a(\rfxs[28] [26]),
    .b(\rfxs[29] [26]),
    .c(_al_u426_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b26/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u428 (
    .a(\mux31_b26/B1_6 ),
    .b(\mux31_b26/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u428_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u429 (
    .a(\mux31_b26/B1_4 ),
    .b(\mux31_b26/B1_5 ),
    .c(_al_u428_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b26/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u430 (
    .a(\rfxs[14] [26]),
    .b(\rfxs[15] [26]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u430_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u431 (
    .a(\rfxs[12] [26]),
    .b(\rfxs[13] [26]),
    .c(_al_u430_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b26/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u432 (
    .a(\rfxs[8] [26]),
    .b(\rfxs[10] [26]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u432_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u433 (
    .a(\rfxs[11] [26]),
    .b(\rfxs[9] [26]),
    .c(_al_u432_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b26/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u434 (
    .a(\mux31_b26/B1_1 ),
    .b(\mux31_b26/B1_2 ),
    .c(_al_u168_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u434_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u435 (
    .a(\mux31_b26/B3_1 ),
    .b(_al_u434_o),
    .c(\mux31_b26/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u435_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u436 (
    .a(n94),
    .b(_al_u435_o),
    .c(i_rd_wdata[26]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[26]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u437 (
    .a(\rfxs[22] [25]),
    .b(\rfxs[23] [25]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u437_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u438 (
    .a(\rfxs[20] [25]),
    .b(\rfxs[21] [25]),
    .c(_al_u437_o),
    .d(i_rs1idx[1]),
    .o(_al_u438_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u439 (
    .a(\rfxs[18] [25]),
    .b(\rfxs[19] [25]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u439_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u440 (
    .a(\rfxs[16] [25]),
    .b(\rfxs[17] [25]),
    .c(_al_u439_o),
    .d(i_rs1idx[1]),
    .o(_al_u440_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u441 (
    .a(\rfxs[1] [25]),
    .b(\rfxs[2] [25]),
    .c(\rfxs[3] [25]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u441_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u442 (
    .a(\rfxs[6] [25]),
    .b(\rfxs[7] [25]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u442_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u443 (
    .a(\rfxs[4] [25]),
    .b(\rfxs[5] [25]),
    .c(_al_u442_o),
    .d(i_rs1idx[1]),
    .o(_al_u443_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f53))
    _al_u444 (
    .a(_al_u443_o),
    .b(_al_u441_o),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[4]),
    .o(_al_u444_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u445 (
    .a(_al_u438_o),
    .b(_al_u440_o),
    .c(_al_u444_o),
    .d(i_rs1idx[4]),
    .o(_al_u445_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55ff0f33))
    _al_u446 (
    .a(\rfxs[11] [25]),
    .b(\rfxs[8] [25]),
    .c(\rfxs[10] [25]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u446_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(C*B))"),
    .INIT(16'h002a))
    _al_u447 (
    .a(_al_u446_o),
    .b(_al_u125_o),
    .c(\rfxs[9] [25]),
    .d(i_rs1idx[2]),
    .o(_al_u447_o));
  AL_MAP_LUT5 #(
    .EQN("(D*(~(A)*~(B)*~(C)*~(E)+A*~(B)*~(C)*~(E)+A*B*~(C)*~(E)+~(A)*~(B)*C*~(E)+~(A)*~(B)*~(C)*E+~(A)*B*~(C)*E+~(A)*~(B)*C*E+~(A)*B*C*E))"),
    .INIT(32'h55001b00))
    _al_u448 (
    .a(_al_u114_o),
    .b(\rfxs[12] [25]),
    .c(\rfxs[13] [25]),
    .d(i_rs1idx[2]),
    .e(i_rs1idx[1]),
    .o(_al_u448_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u449 (
    .a(\rfxs[29] [25]),
    .b(\rfxs[30] [25]),
    .c(\rfxs[31] [25]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u449_o));
  AL_MAP_LUT4 #(
    .EQN("(D*A*~(C*B))"),
    .INIT(16'h2a00))
    _al_u450 (
    .a(_al_u449_o),
    .b(_al_u116_o),
    .c(\rfxs[28] [25]),
    .d(i_rs1idx[2]),
    .o(_al_u450_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u451 (
    .a(\rfxs[25] [25]),
    .b(\rfxs[26] [25]),
    .c(\rfxs[27] [25]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u451_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(C*B))"),
    .INIT(16'h002a))
    _al_u452 (
    .a(_al_u451_o),
    .b(_al_u116_o),
    .c(\rfxs[24] [25]),
    .d(i_rs1idx[2]),
    .o(_al_u452_o));
  AL_MAP_LUT5 #(
    .EQN("~((~D*~A)*~((~C*~B))*~(E)+(~D*~A)*(~C*~B)*~(E)+~((~D*~A))*(~C*~B)*E+(~D*~A)*(~C*~B)*E)"),
    .INIT(32'hfcfcffaa))
    _al_u453 (
    .a(_al_u447_o),
    .b(_al_u450_o),
    .c(_al_u452_o),
    .d(_al_u448_o),
    .e(i_rs1idx[4]),
    .o(_al_u453_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u454 (
    .a(_al_u445_o),
    .b(_al_u453_o),
    .c(i_rs1idx[3]),
    .o(_al_u454_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u455 (
    .a(n94),
    .b(_al_u454_o),
    .c(i_rd_wdata[25]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[25]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u456 (
    .a(\rfxs[26] [24]),
    .b(\rfxs[27] [24]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u456_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u457 (
    .a(\rfxs[24] [24]),
    .b(\rfxs[25] [24]),
    .c(_al_u456_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b24/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u458 (
    .a(\rfxs[30] [24]),
    .b(\rfxs[31] [24]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u458_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u459 (
    .a(\rfxs[28] [24]),
    .b(\rfxs[29] [24]),
    .c(_al_u458_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b24/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u460 (
    .a(\mux31_b24/B1_6 ),
    .b(\mux31_b24/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u460_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u461 (
    .a(\mux31_b24/B1_4 ),
    .b(\mux31_b24/B1_5 ),
    .c(_al_u460_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b24/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u462 (
    .a(\rfxs[14] [24]),
    .b(\rfxs[15] [24]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u462_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u463 (
    .a(\rfxs[12] [24]),
    .b(\rfxs[13] [24]),
    .c(_al_u462_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b24/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u464 (
    .a(\rfxs[8] [24]),
    .b(\rfxs[10] [24]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u464_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u465 (
    .a(\rfxs[11] [24]),
    .b(\rfxs[9] [24]),
    .c(_al_u464_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b24/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u466 (
    .a(\mux31_b24/B1_1 ),
    .b(\mux31_b24/B1_2 ),
    .c(_al_u175_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u466_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u467 (
    .a(\mux31_b24/B3_1 ),
    .b(_al_u466_o),
    .c(\mux31_b24/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u467_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u468 (
    .a(n94),
    .b(_al_u467_o),
    .c(i_rd_wdata[24]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[24]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u469 (
    .a(\rfxs[26] [23]),
    .b(\rfxs[27] [23]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u469_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u470 (
    .a(\rfxs[24] [23]),
    .b(\rfxs[25] [23]),
    .c(_al_u469_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b23/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u471 (
    .a(\rfxs[30] [23]),
    .b(\rfxs[31] [23]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u471_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u472 (
    .a(\rfxs[28] [23]),
    .b(\rfxs[29] [23]),
    .c(_al_u471_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b23/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u473 (
    .a(\mux31_b23/B1_6 ),
    .b(\mux31_b23/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u473_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u474 (
    .a(\mux31_b23/B1_4 ),
    .b(\mux31_b23/B1_5 ),
    .c(_al_u473_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b23/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u475 (
    .a(\rfxs[14] [23]),
    .b(\rfxs[15] [23]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u475_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u476 (
    .a(\rfxs[12] [23]),
    .b(\rfxs[13] [23]),
    .c(_al_u475_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b23/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u477 (
    .a(\rfxs[8] [23]),
    .b(\rfxs[10] [23]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u477_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u478 (
    .a(\rfxs[11] [23]),
    .b(\rfxs[9] [23]),
    .c(_al_u477_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b23/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u479 (
    .a(\mux31_b23/B1_1 ),
    .b(\mux31_b23/B1_2 ),
    .c(_al_u182_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u479_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u480 (
    .a(\mux31_b23/B3_1 ),
    .b(_al_u479_o),
    .c(\mux31_b23/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u480_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u481 (
    .a(n94),
    .b(_al_u480_o),
    .c(i_rd_wdata[23]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[23]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u482 (
    .a(\rfxs[22] [22]),
    .b(\rfxs[23] [22]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u482_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u483 (
    .a(\rfxs[20] [22]),
    .b(\rfxs[21] [22]),
    .c(_al_u482_o),
    .d(i_rs1idx[1]),
    .o(_al_u483_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u484 (
    .a(\rfxs[18] [22]),
    .b(\rfxs[19] [22]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u484_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u485 (
    .a(\rfxs[16] [22]),
    .b(\rfxs[17] [22]),
    .c(_al_u484_o),
    .d(i_rs1idx[1]),
    .o(_al_u485_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u486 (
    .a(_al_u483_o),
    .b(_al_u485_o),
    .c(i_rs1idx[2]),
    .o(_al_u486_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u487 (
    .a(\rfxs[1] [22]),
    .b(\rfxs[2] [22]),
    .c(\rfxs[3] [22]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u487_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u488 (
    .a(\rfxs[5] [22]),
    .b(\rfxs[6] [22]),
    .c(\rfxs[7] [22]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u488_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u489 (
    .a(_al_u487_o),
    .b(_al_u488_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [22]),
    .e(i_rs1idx[2]),
    .o(_al_u489_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u490 (
    .a(_al_u486_o),
    .b(_al_u489_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u490_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u491 (
    .a(\rfxs[8] [22]),
    .b(\rfxs[10] [22]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u491_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u492 (
    .a(\rfxs[11] [22]),
    .b(\rfxs[9] [22]),
    .c(_al_u491_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b22/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u493 (
    .a(\rfxs[14] [22]),
    .b(\rfxs[15] [22]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u493_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u494 (
    .a(\rfxs[12] [22]),
    .b(\rfxs[13] [22]),
    .c(_al_u493_o),
    .d(i_rs1idx[1]),
    .o(_al_u494_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u495 (
    .a(\mux31_b22/B1_2 ),
    .b(_al_u494_o),
    .c(i_rs1idx[2]),
    .o(_al_u495_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u496 (
    .a(\rfxs[30] [22]),
    .b(\rfxs[31] [22]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u496_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u497 (
    .a(\rfxs[28] [22]),
    .b(\rfxs[29] [22]),
    .c(_al_u496_o),
    .d(i_rs1idx[1]),
    .o(_al_u497_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u498 (
    .a(\rfxs[26] [22]),
    .b(\rfxs[27] [22]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u498_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u499 (
    .a(\rfxs[24] [22]),
    .b(\rfxs[25] [22]),
    .c(_al_u498_o),
    .d(i_rs1idx[1]),
    .o(_al_u499_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u500 (
    .a(_al_u497_o),
    .b(_al_u499_o),
    .c(i_rs1idx[2]),
    .o(_al_u500_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u501 (
    .a(_al_u495_o),
    .b(_al_u500_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u501_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u502 (
    .a(n94),
    .b(_al_u501_o),
    .c(_al_u490_o),
    .d(i_rd_wdata[22]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[22]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u503 (
    .a(\rfxs[22] [21]),
    .b(\rfxs[23] [21]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u503_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u504 (
    .a(\rfxs[20] [21]),
    .b(\rfxs[21] [21]),
    .c(_al_u503_o),
    .d(i_rs1idx[1]),
    .o(_al_u504_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u505 (
    .a(\rfxs[18] [21]),
    .b(\rfxs[19] [21]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u505_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u506 (
    .a(\rfxs[16] [21]),
    .b(\rfxs[17] [21]),
    .c(_al_u505_o),
    .d(i_rs1idx[1]),
    .o(_al_u506_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u507 (
    .a(_al_u504_o),
    .b(_al_u506_o),
    .c(i_rs1idx[2]),
    .o(_al_u507_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u508 (
    .a(\rfxs[1] [21]),
    .b(\rfxs[2] [21]),
    .c(\rfxs[3] [21]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u508_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u509 (
    .a(\rfxs[5] [21]),
    .b(\rfxs[6] [21]),
    .c(\rfxs[7] [21]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u509_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u510 (
    .a(_al_u508_o),
    .b(_al_u509_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [21]),
    .e(i_rs1idx[2]),
    .o(_al_u510_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u511 (
    .a(_al_u507_o),
    .b(_al_u510_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u511_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u512 (
    .a(\rfxs[8] [21]),
    .b(\rfxs[10] [21]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u512_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u513 (
    .a(\rfxs[11] [21]),
    .b(\rfxs[9] [21]),
    .c(_al_u512_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b21/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u514 (
    .a(\rfxs[14] [21]),
    .b(\rfxs[15] [21]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u514_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u515 (
    .a(\rfxs[12] [21]),
    .b(\rfxs[13] [21]),
    .c(_al_u514_o),
    .d(i_rs1idx[1]),
    .o(_al_u515_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u516 (
    .a(\mux31_b21/B1_2 ),
    .b(_al_u515_o),
    .c(i_rs1idx[2]),
    .o(_al_u516_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u517 (
    .a(\rfxs[30] [21]),
    .b(\rfxs[31] [21]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u517_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u518 (
    .a(\rfxs[28] [21]),
    .b(\rfxs[29] [21]),
    .c(_al_u517_o),
    .d(i_rs1idx[1]),
    .o(_al_u518_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u519 (
    .a(\rfxs[26] [21]),
    .b(\rfxs[27] [21]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u519_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u520 (
    .a(\rfxs[24] [21]),
    .b(\rfxs[25] [21]),
    .c(_al_u519_o),
    .d(i_rs1idx[1]),
    .o(_al_u520_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u521 (
    .a(_al_u518_o),
    .b(_al_u520_o),
    .c(i_rs1idx[2]),
    .o(_al_u521_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u522 (
    .a(_al_u516_o),
    .b(_al_u521_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u522_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u523 (
    .a(n94),
    .b(_al_u522_o),
    .c(_al_u511_o),
    .d(i_rd_wdata[21]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[21]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u524 (
    .a(\rfxs[22] [20]),
    .b(\rfxs[23] [20]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u524_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u525 (
    .a(\rfxs[20] [20]),
    .b(\rfxs[21] [20]),
    .c(_al_u524_o),
    .d(i_rs1idx[1]),
    .o(_al_u525_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u526 (
    .a(\rfxs[18] [20]),
    .b(\rfxs[19] [20]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u526_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u527 (
    .a(\rfxs[16] [20]),
    .b(\rfxs[17] [20]),
    .c(_al_u526_o),
    .d(i_rs1idx[1]),
    .o(_al_u527_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u528 (
    .a(_al_u525_o),
    .b(_al_u527_o),
    .c(i_rs1idx[2]),
    .o(_al_u528_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u529 (
    .a(\rfxs[1] [20]),
    .b(\rfxs[2] [20]),
    .c(\rfxs[3] [20]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u529_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u530 (
    .a(\rfxs[5] [20]),
    .b(\rfxs[6] [20]),
    .c(\rfxs[7] [20]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u530_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u531 (
    .a(_al_u529_o),
    .b(_al_u530_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [20]),
    .e(i_rs1idx[2]),
    .o(_al_u531_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u532 (
    .a(_al_u528_o),
    .b(_al_u531_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u532_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u533 (
    .a(\rfxs[8] [20]),
    .b(\rfxs[10] [20]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u533_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u534 (
    .a(\rfxs[11] [20]),
    .b(\rfxs[9] [20]),
    .c(_al_u533_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b20/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u535 (
    .a(\rfxs[14] [20]),
    .b(\rfxs[15] [20]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u535_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u536 (
    .a(\rfxs[12] [20]),
    .b(\rfxs[13] [20]),
    .c(_al_u535_o),
    .d(i_rs1idx[1]),
    .o(_al_u536_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u537 (
    .a(\mux31_b20/B1_2 ),
    .b(_al_u536_o),
    .c(i_rs1idx[2]),
    .o(_al_u537_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u538 (
    .a(\rfxs[30] [20]),
    .b(\rfxs[31] [20]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u538_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u539 (
    .a(\rfxs[28] [20]),
    .b(\rfxs[29] [20]),
    .c(_al_u538_o),
    .d(i_rs1idx[1]),
    .o(_al_u539_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u540 (
    .a(\rfxs[26] [20]),
    .b(\rfxs[27] [20]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u540_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u541 (
    .a(\rfxs[24] [20]),
    .b(\rfxs[25] [20]),
    .c(_al_u540_o),
    .d(i_rs1idx[1]),
    .o(_al_u541_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u542 (
    .a(_al_u539_o),
    .b(_al_u541_o),
    .c(i_rs1idx[2]),
    .o(_al_u542_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u543 (
    .a(_al_u537_o),
    .b(_al_u542_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u543_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u544 (
    .a(n94),
    .b(_al_u543_o),
    .c(_al_u532_o),
    .d(i_rd_wdata[20]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[20]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u545 (
    .a(\rfxs[22] [2]),
    .b(\rfxs[23] [2]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u545_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u546 (
    .a(\rfxs[20] [2]),
    .b(\rfxs[21] [2]),
    .c(_al_u545_o),
    .d(i_rs1idx[1]),
    .o(_al_u546_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u547 (
    .a(\rfxs[18] [2]),
    .b(\rfxs[19] [2]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u547_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u548 (
    .a(\rfxs[16] [2]),
    .b(\rfxs[17] [2]),
    .c(_al_u547_o),
    .d(i_rs1idx[1]),
    .o(_al_u548_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u549 (
    .a(_al_u546_o),
    .b(_al_u548_o),
    .c(i_rs1idx[2]),
    .o(_al_u549_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u550 (
    .a(\rfxs[1] [2]),
    .b(\rfxs[2] [2]),
    .c(\rfxs[3] [2]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u550_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u551 (
    .a(\rfxs[5] [2]),
    .b(\rfxs[6] [2]),
    .c(\rfxs[7] [2]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u551_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u552 (
    .a(_al_u550_o),
    .b(_al_u551_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [2]),
    .e(i_rs1idx[2]),
    .o(_al_u552_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u553 (
    .a(_al_u549_o),
    .b(_al_u552_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u553_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u554 (
    .a(\rfxs[8] [2]),
    .b(\rfxs[10] [2]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u554_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u555 (
    .a(\rfxs[11] [2]),
    .b(\rfxs[9] [2]),
    .c(_al_u554_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b2/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u556 (
    .a(\rfxs[14] [2]),
    .b(\rfxs[15] [2]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u556_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u557 (
    .a(\rfxs[12] [2]),
    .b(\rfxs[13] [2]),
    .c(_al_u556_o),
    .d(i_rs1idx[1]),
    .o(_al_u557_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u558 (
    .a(\mux31_b2/B1_2 ),
    .b(_al_u557_o),
    .c(i_rs1idx[2]),
    .o(_al_u558_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u559 (
    .a(\rfxs[26] [2]),
    .b(\rfxs[27] [2]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u559_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u560 (
    .a(\rfxs[24] [2]),
    .b(\rfxs[25] [2]),
    .c(_al_u559_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b2/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u561 (
    .a(\rfxs[30] [2]),
    .b(\rfxs[31] [2]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u561_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u562 (
    .a(\rfxs[28] [2]),
    .b(\rfxs[29] [2]),
    .c(_al_u561_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b2/B1_7 ));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u563 (
    .a(\mux31_b2/B1_6 ),
    .b(\mux31_b2/B1_7 ),
    .c(i_rs1idx[2]),
    .o(_al_u563_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u564 (
    .a(_al_u558_o),
    .b(_al_u563_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u564_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u565 (
    .a(n94),
    .b(_al_u564_o),
    .c(_al_u553_o),
    .d(i_rd_wdata[2]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[2]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u566 (
    .a(\rfxs[22] [19]),
    .b(\rfxs[23] [19]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u566_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u567 (
    .a(\rfxs[20] [19]),
    .b(\rfxs[21] [19]),
    .c(_al_u566_o),
    .d(i_rs1idx[1]),
    .o(_al_u567_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u568 (
    .a(\rfxs[18] [19]),
    .b(\rfxs[19] [19]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u568_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u569 (
    .a(\rfxs[16] [19]),
    .b(\rfxs[17] [19]),
    .c(_al_u568_o),
    .d(i_rs1idx[1]),
    .o(_al_u569_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u570 (
    .a(_al_u567_o),
    .b(_al_u569_o),
    .c(i_rs1idx[2]),
    .o(_al_u570_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u571 (
    .a(\rfxs[1] [19]),
    .b(\rfxs[2] [19]),
    .c(\rfxs[3] [19]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u571_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u572 (
    .a(\rfxs[5] [19]),
    .b(\rfxs[6] [19]),
    .c(\rfxs[7] [19]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u572_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u573 (
    .a(_al_u571_o),
    .b(_al_u572_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [19]),
    .e(i_rs1idx[2]),
    .o(_al_u573_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u574 (
    .a(_al_u570_o),
    .b(_al_u573_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u574_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u575 (
    .a(\rfxs[8] [19]),
    .b(\rfxs[10] [19]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u575_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u576 (
    .a(\rfxs[11] [19]),
    .b(\rfxs[9] [19]),
    .c(_al_u575_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b19/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u577 (
    .a(\rfxs[14] [19]),
    .b(\rfxs[15] [19]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u577_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u578 (
    .a(\rfxs[12] [19]),
    .b(\rfxs[13] [19]),
    .c(_al_u577_o),
    .d(i_rs1idx[1]),
    .o(_al_u578_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u579 (
    .a(\mux31_b19/B1_2 ),
    .b(_al_u578_o),
    .c(i_rs1idx[2]),
    .o(_al_u579_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u580 (
    .a(\rfxs[30] [19]),
    .b(\rfxs[31] [19]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u580_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u581 (
    .a(\rfxs[28] [19]),
    .b(\rfxs[29] [19]),
    .c(_al_u580_o),
    .d(i_rs1idx[1]),
    .o(_al_u581_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u582 (
    .a(\rfxs[26] [19]),
    .b(\rfxs[27] [19]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u582_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u583 (
    .a(\rfxs[24] [19]),
    .b(\rfxs[25] [19]),
    .c(_al_u582_o),
    .d(i_rs1idx[1]),
    .o(_al_u583_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u584 (
    .a(_al_u581_o),
    .b(_al_u583_o),
    .c(i_rs1idx[2]),
    .o(_al_u584_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u585 (
    .a(_al_u579_o),
    .b(_al_u584_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u585_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u586 (
    .a(n94),
    .b(_al_u585_o),
    .c(_al_u574_o),
    .d(i_rd_wdata[19]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[19]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u587 (
    .a(\rfxs[22] [18]),
    .b(\rfxs[23] [18]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u587_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u588 (
    .a(\rfxs[20] [18]),
    .b(\rfxs[21] [18]),
    .c(_al_u587_o),
    .d(i_rs1idx[1]),
    .o(_al_u588_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u589 (
    .a(\rfxs[18] [18]),
    .b(\rfxs[19] [18]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u589_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u590 (
    .a(\rfxs[16] [18]),
    .b(\rfxs[17] [18]),
    .c(_al_u589_o),
    .d(i_rs1idx[1]),
    .o(_al_u590_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u591 (
    .a(\rfxs[1] [18]),
    .b(\rfxs[2] [18]),
    .c(\rfxs[3] [18]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u591_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u592 (
    .a(\rfxs[6] [18]),
    .b(\rfxs[7] [18]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u592_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u593 (
    .a(\rfxs[4] [18]),
    .b(\rfxs[5] [18]),
    .c(_al_u592_o),
    .d(i_rs1idx[1]),
    .o(_al_u593_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f53))
    _al_u594 (
    .a(_al_u593_o),
    .b(_al_u591_o),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[4]),
    .o(_al_u594_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u595 (
    .a(_al_u588_o),
    .b(_al_u590_o),
    .c(_al_u594_o),
    .d(i_rs1idx[4]),
    .o(_al_u595_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h55ff0f33))
    _al_u596 (
    .a(\rfxs[11] [18]),
    .b(\rfxs[8] [18]),
    .c(\rfxs[10] [18]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u596_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(C*B))"),
    .INIT(16'h002a))
    _al_u597 (
    .a(_al_u596_o),
    .b(_al_u125_o),
    .c(\rfxs[9] [18]),
    .d(i_rs1idx[2]),
    .o(_al_u597_o));
  AL_MAP_LUT5 #(
    .EQN("(D*(~(A)*~(B)*~(C)*~(E)+A*~(B)*~(C)*~(E)+A*B*~(C)*~(E)+~(A)*~(B)*C*~(E)+~(A)*~(B)*~(C)*E+~(A)*B*~(C)*E+~(A)*~(B)*C*E+~(A)*B*C*E))"),
    .INIT(32'h55001b00))
    _al_u598 (
    .a(_al_u115_o),
    .b(\rfxs[12] [18]),
    .c(\rfxs[13] [18]),
    .d(i_rs1idx[2]),
    .e(i_rs1idx[1]),
    .o(_al_u598_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u599 (
    .a(\rfxs[29] [18]),
    .b(\rfxs[30] [18]),
    .c(\rfxs[31] [18]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u599_o));
  AL_MAP_LUT4 #(
    .EQN("(D*A*~(C*B))"),
    .INIT(16'h2a00))
    _al_u600 (
    .a(_al_u599_o),
    .b(_al_u116_o),
    .c(\rfxs[28] [18]),
    .d(i_rs1idx[2]),
    .o(_al_u600_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u601 (
    .a(\rfxs[25] [18]),
    .b(\rfxs[26] [18]),
    .c(\rfxs[27] [18]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u601_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(C*B))"),
    .INIT(16'h002a))
    _al_u602 (
    .a(_al_u601_o),
    .b(_al_u116_o),
    .c(\rfxs[24] [18]),
    .d(i_rs1idx[2]),
    .o(_al_u602_o));
  AL_MAP_LUT5 #(
    .EQN("~((~D*~A)*~((~C*~B))*~(E)+(~D*~A)*(~C*~B)*~(E)+~((~D*~A))*(~C*~B)*E+(~D*~A)*(~C*~B)*E)"),
    .INIT(32'hfcfcffaa))
    _al_u603 (
    .a(_al_u597_o),
    .b(_al_u600_o),
    .c(_al_u602_o),
    .d(_al_u598_o),
    .e(i_rs1idx[4]),
    .o(_al_u603_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'hca))
    _al_u604 (
    .a(_al_u595_o),
    .b(_al_u603_o),
    .c(i_rs1idx[3]),
    .o(_al_u604_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u605 (
    .a(n94),
    .b(_al_u604_o),
    .c(i_rd_wdata[18]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[18]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u606 (
    .a(\rfxs[22] [17]),
    .b(\rfxs[23] [17]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u606_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u607 (
    .a(\rfxs[20] [17]),
    .b(\rfxs[21] [17]),
    .c(_al_u606_o),
    .d(i_rs1idx[1]),
    .o(_al_u607_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u608 (
    .a(\rfxs[18] [17]),
    .b(\rfxs[19] [17]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u608_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u609 (
    .a(\rfxs[16] [17]),
    .b(\rfxs[17] [17]),
    .c(_al_u608_o),
    .d(i_rs1idx[1]),
    .o(_al_u609_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u610 (
    .a(_al_u607_o),
    .b(_al_u609_o),
    .c(i_rs1idx[2]),
    .o(_al_u610_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u611 (
    .a(\rfxs[1] [17]),
    .b(\rfxs[2] [17]),
    .c(\rfxs[3] [17]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u611_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u612 (
    .a(\rfxs[5] [17]),
    .b(\rfxs[6] [17]),
    .c(\rfxs[7] [17]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u612_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u613 (
    .a(_al_u611_o),
    .b(_al_u612_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [17]),
    .e(i_rs1idx[2]),
    .o(_al_u613_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u614 (
    .a(_al_u610_o),
    .b(_al_u613_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u614_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u615 (
    .a(\rfxs[8] [17]),
    .b(\rfxs[10] [17]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u615_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u616 (
    .a(\rfxs[11] [17]),
    .b(\rfxs[9] [17]),
    .c(_al_u615_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b17/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u617 (
    .a(\rfxs[14] [17]),
    .b(\rfxs[15] [17]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u617_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u618 (
    .a(\rfxs[12] [17]),
    .b(\rfxs[13] [17]),
    .c(_al_u617_o),
    .d(i_rs1idx[1]),
    .o(_al_u618_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u619 (
    .a(\mux31_b17/B1_2 ),
    .b(_al_u618_o),
    .c(i_rs1idx[2]),
    .o(_al_u619_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u620 (
    .a(\rfxs[30] [17]),
    .b(\rfxs[31] [17]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u620_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u621 (
    .a(\rfxs[28] [17]),
    .b(\rfxs[29] [17]),
    .c(_al_u620_o),
    .d(i_rs1idx[1]),
    .o(_al_u621_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u622 (
    .a(\rfxs[26] [17]),
    .b(\rfxs[27] [17]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u622_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u623 (
    .a(\rfxs[24] [17]),
    .b(\rfxs[25] [17]),
    .c(_al_u622_o),
    .d(i_rs1idx[1]),
    .o(_al_u623_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u624 (
    .a(_al_u621_o),
    .b(_al_u623_o),
    .c(i_rs1idx[2]),
    .o(_al_u624_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u625 (
    .a(_al_u619_o),
    .b(_al_u624_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u625_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u626 (
    .a(n94),
    .b(_al_u625_o),
    .c(_al_u614_o),
    .d(i_rd_wdata[17]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[17]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u627 (
    .a(\rfxs[26] [16]),
    .b(\rfxs[27] [16]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u627_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u628 (
    .a(\rfxs[24] [16]),
    .b(\rfxs[25] [16]),
    .c(_al_u627_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b16/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u629 (
    .a(\rfxs[30] [16]),
    .b(\rfxs[31] [16]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u629_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u630 (
    .a(\rfxs[28] [16]),
    .b(\rfxs[29] [16]),
    .c(_al_u629_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b16/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u631 (
    .a(\mux31_b16/B1_6 ),
    .b(\mux31_b16/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u631_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u632 (
    .a(\mux31_b16/B1_4 ),
    .b(\mux31_b16/B1_5 ),
    .c(_al_u631_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b16/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u633 (
    .a(\rfxs[14] [16]),
    .b(\rfxs[15] [16]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u633_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u634 (
    .a(\rfxs[12] [16]),
    .b(\rfxs[13] [16]),
    .c(_al_u633_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b16/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u635 (
    .a(\rfxs[8] [16]),
    .b(\rfxs[10] [16]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u635_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u636 (
    .a(\rfxs[11] [16]),
    .b(\rfxs[9] [16]),
    .c(_al_u635_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b16/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u637 (
    .a(\mux31_b16/B1_1 ),
    .b(\mux31_b16/B1_2 ),
    .c(_al_u189_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u637_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u638 (
    .a(\mux31_b16/B3_1 ),
    .b(_al_u637_o),
    .c(\mux31_b16/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u638_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u639 (
    .a(n94),
    .b(_al_u638_o),
    .c(i_rd_wdata[16]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[16]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u640 (
    .a(\rfxs[26] [15]),
    .b(\rfxs[27] [15]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u640_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u641 (
    .a(\rfxs[24] [15]),
    .b(\rfxs[25] [15]),
    .c(_al_u640_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b15/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u642 (
    .a(\rfxs[30] [15]),
    .b(\rfxs[31] [15]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u642_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u643 (
    .a(\rfxs[28] [15]),
    .b(\rfxs[29] [15]),
    .c(_al_u642_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b15/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u644 (
    .a(\mux31_b15/B1_6 ),
    .b(\mux31_b15/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u644_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u645 (
    .a(\mux31_b15/B1_4 ),
    .b(\mux31_b15/B1_5 ),
    .c(_al_u644_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b15/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u646 (
    .a(\rfxs[14] [15]),
    .b(\rfxs[15] [15]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u646_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u647 (
    .a(\rfxs[12] [15]),
    .b(\rfxs[13] [15]),
    .c(_al_u646_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b15/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u648 (
    .a(\rfxs[8] [15]),
    .b(\rfxs[10] [15]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u648_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u649 (
    .a(\rfxs[11] [15]),
    .b(\rfxs[9] [15]),
    .c(_al_u648_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b15/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u650 (
    .a(\mux31_b15/B1_1 ),
    .b(\mux31_b15/B1_2 ),
    .c(_al_u196_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u650_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u651 (
    .a(\mux31_b15/B3_1 ),
    .b(_al_u650_o),
    .c(\mux31_b15/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u651_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u652 (
    .a(n94),
    .b(_al_u651_o),
    .c(i_rd_wdata[15]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[15]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u653 (
    .a(\rfxs[26] [14]),
    .b(\rfxs[27] [14]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u653_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u654 (
    .a(\rfxs[24] [14]),
    .b(\rfxs[25] [14]),
    .c(_al_u653_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b14/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u655 (
    .a(\rfxs[30] [14]),
    .b(\rfxs[31] [14]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u655_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u656 (
    .a(\rfxs[28] [14]),
    .b(\rfxs[29] [14]),
    .c(_al_u655_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b14/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u657 (
    .a(\mux31_b14/B1_6 ),
    .b(\mux31_b14/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u657_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u658 (
    .a(\mux31_b14/B1_4 ),
    .b(\mux31_b14/B1_5 ),
    .c(_al_u657_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b14/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u659 (
    .a(\rfxs[14] [14]),
    .b(\rfxs[15] [14]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u659_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u660 (
    .a(\rfxs[12] [14]),
    .b(\rfxs[13] [14]),
    .c(_al_u659_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b14/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u661 (
    .a(\rfxs[8] [14]),
    .b(\rfxs[10] [14]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u661_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u662 (
    .a(\rfxs[11] [14]),
    .b(\rfxs[9] [14]),
    .c(_al_u661_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b14/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u663 (
    .a(\mux31_b14/B1_1 ),
    .b(\mux31_b14/B1_2 ),
    .c(_al_u203_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u663_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u664 (
    .a(\mux31_b14/B3_1 ),
    .b(_al_u663_o),
    .c(\mux31_b14/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u664_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u665 (
    .a(n94),
    .b(_al_u664_o),
    .c(i_rd_wdata[14]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[14]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u666 (
    .a(\rfxs[26] [13]),
    .b(\rfxs[27] [13]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u666_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u667 (
    .a(\rfxs[24] [13]),
    .b(\rfxs[25] [13]),
    .c(_al_u666_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b13/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u668 (
    .a(\rfxs[30] [13]),
    .b(\rfxs[31] [13]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u668_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u669 (
    .a(\rfxs[28] [13]),
    .b(\rfxs[29] [13]),
    .c(_al_u668_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b13/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u670 (
    .a(\mux31_b13/B1_6 ),
    .b(\mux31_b13/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u670_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u671 (
    .a(\mux31_b13/B1_4 ),
    .b(\mux31_b13/B1_5 ),
    .c(_al_u670_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b13/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u672 (
    .a(\rfxs[14] [13]),
    .b(\rfxs[15] [13]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u672_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u673 (
    .a(\rfxs[12] [13]),
    .b(\rfxs[13] [13]),
    .c(_al_u672_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b13/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u674 (
    .a(\rfxs[8] [13]),
    .b(\rfxs[10] [13]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u674_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u675 (
    .a(\rfxs[11] [13]),
    .b(\rfxs[9] [13]),
    .c(_al_u674_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b13/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u676 (
    .a(\mux31_b13/B1_1 ),
    .b(\mux31_b13/B1_2 ),
    .c(_al_u210_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u676_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u677 (
    .a(\mux31_b13/B3_1 ),
    .b(_al_u676_o),
    .c(\mux31_b13/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u677_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u678 (
    .a(n94),
    .b(_al_u677_o),
    .c(i_rd_wdata[13]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[13]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u679 (
    .a(\rfxs[26] [12]),
    .b(\rfxs[27] [12]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u679_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u680 (
    .a(\rfxs[24] [12]),
    .b(\rfxs[25] [12]),
    .c(_al_u679_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b12/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u681 (
    .a(\rfxs[30] [12]),
    .b(\rfxs[31] [12]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u681_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u682 (
    .a(\rfxs[28] [12]),
    .b(\rfxs[29] [12]),
    .c(_al_u681_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b12/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u683 (
    .a(\mux31_b12/B1_6 ),
    .b(\mux31_b12/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u683_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u684 (
    .a(\mux31_b12/B1_4 ),
    .b(\mux31_b12/B1_5 ),
    .c(_al_u683_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b12/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u685 (
    .a(\rfxs[14] [12]),
    .b(\rfxs[15] [12]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u685_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u686 (
    .a(\rfxs[12] [12]),
    .b(\rfxs[13] [12]),
    .c(_al_u685_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b12/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u687 (
    .a(\rfxs[8] [12]),
    .b(\rfxs[10] [12]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u687_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u688 (
    .a(\rfxs[11] [12]),
    .b(\rfxs[9] [12]),
    .c(_al_u687_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b12/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u689 (
    .a(\mux31_b12/B1_1 ),
    .b(\mux31_b12/B1_2 ),
    .c(_al_u217_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u689_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u690 (
    .a(\mux31_b12/B3_1 ),
    .b(_al_u689_o),
    .c(\mux31_b12/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u690_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u691 (
    .a(n94),
    .b(_al_u690_o),
    .c(i_rd_wdata[12]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[12]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u692 (
    .a(\rfxs[22] [11]),
    .b(\rfxs[23] [11]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u692_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u693 (
    .a(\rfxs[20] [11]),
    .b(\rfxs[21] [11]),
    .c(_al_u692_o),
    .d(i_rs1idx[1]),
    .o(_al_u693_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u694 (
    .a(\rfxs[17] [11]),
    .b(\rfxs[18] [11]),
    .c(\rfxs[19] [11]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u694_o));
  AL_MAP_LUT5 #(
    .EQN("((B*~(D*C))*~(A)*~(E)+(B*~(D*C))*A*~(E)+~((B*~(D*C)))*A*E+(B*~(D*C))*A*E)"),
    .INIT(32'haaaa0ccc))
    _al_u695 (
    .a(_al_u693_o),
    .b(_al_u694_o),
    .c(_al_u116_o),
    .d(\rfxs[16] [11]),
    .e(i_rs1idx[2]),
    .o(_al_u695_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u696 (
    .a(\rfxs[1] [11]),
    .b(\rfxs[2] [11]),
    .c(\rfxs[3] [11]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u696_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u697 (
    .a(\rfxs[5] [11]),
    .b(\rfxs[6] [11]),
    .c(\rfxs[7] [11]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u697_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u698 (
    .a(_al_u696_o),
    .b(_al_u697_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [11]),
    .e(i_rs1idx[2]),
    .o(_al_u698_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u699 (
    .a(_al_u695_o),
    .b(_al_u698_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u699_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u700 (
    .a(\rfxs[8] [11]),
    .b(\rfxs[10] [11]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u700_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u701 (
    .a(\rfxs[11] [11]),
    .b(\rfxs[9] [11]),
    .c(_al_u700_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b11/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u702 (
    .a(\rfxs[14] [11]),
    .b(\rfxs[15] [11]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u702_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u703 (
    .a(\rfxs[12] [11]),
    .b(\rfxs[13] [11]),
    .c(_al_u702_o),
    .d(i_rs1idx[1]),
    .o(_al_u703_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u704 (
    .a(\mux31_b11/B1_2 ),
    .b(_al_u703_o),
    .c(i_rs1idx[2]),
    .o(_al_u704_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u705 (
    .a(\rfxs[30] [11]),
    .b(\rfxs[31] [11]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u705_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u706 (
    .a(\rfxs[28] [11]),
    .b(\rfxs[29] [11]),
    .c(_al_u705_o),
    .d(i_rs1idx[1]),
    .o(_al_u706_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u707 (
    .a(\rfxs[26] [11]),
    .b(\rfxs[27] [11]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u707_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u708 (
    .a(\rfxs[24] [11]),
    .b(\rfxs[25] [11]),
    .c(_al_u707_o),
    .d(i_rs1idx[1]),
    .o(_al_u708_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u709 (
    .a(_al_u706_o),
    .b(_al_u708_o),
    .c(i_rs1idx[2]),
    .o(_al_u709_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u710 (
    .a(_al_u704_o),
    .b(_al_u709_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u710_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u711 (
    .a(n94),
    .b(_al_u710_o),
    .c(_al_u699_o),
    .d(i_rd_wdata[11]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[11]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u712 (
    .a(\rfxs[22] [10]),
    .b(\rfxs[23] [10]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u712_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u713 (
    .a(\rfxs[20] [10]),
    .b(\rfxs[21] [10]),
    .c(_al_u712_o),
    .d(i_rs1idx[1]),
    .o(_al_u713_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u714 (
    .a(\rfxs[17] [10]),
    .b(\rfxs[18] [10]),
    .c(\rfxs[19] [10]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u714_o));
  AL_MAP_LUT5 #(
    .EQN("((B*~(D*C))*~(A)*~(E)+(B*~(D*C))*A*~(E)+~((B*~(D*C)))*A*E+(B*~(D*C))*A*E)"),
    .INIT(32'haaaa0ccc))
    _al_u715 (
    .a(_al_u713_o),
    .b(_al_u714_o),
    .c(_al_u116_o),
    .d(\rfxs[16] [10]),
    .e(i_rs1idx[2]),
    .o(_al_u715_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u716 (
    .a(\rfxs[1] [10]),
    .b(\rfxs[2] [10]),
    .c(\rfxs[3] [10]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u716_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u717 (
    .a(\rfxs[5] [10]),
    .b(\rfxs[6] [10]),
    .c(\rfxs[7] [10]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u717_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u718 (
    .a(_al_u716_o),
    .b(_al_u717_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [10]),
    .e(i_rs1idx[2]),
    .o(_al_u718_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u719 (
    .a(_al_u715_o),
    .b(_al_u718_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u719_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u720 (
    .a(\rfxs[8] [10]),
    .b(\rfxs[10] [10]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u720_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u721 (
    .a(\rfxs[11] [10]),
    .b(\rfxs[9] [10]),
    .c(_al_u720_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b10/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u722 (
    .a(\rfxs[14] [10]),
    .b(\rfxs[15] [10]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u722_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u723 (
    .a(\rfxs[12] [10]),
    .b(\rfxs[13] [10]),
    .c(_al_u722_o),
    .d(i_rs1idx[1]),
    .o(_al_u723_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u724 (
    .a(\mux31_b10/B1_2 ),
    .b(_al_u723_o),
    .c(i_rs1idx[2]),
    .o(_al_u724_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u725 (
    .a(\rfxs[30] [10]),
    .b(\rfxs[31] [10]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u725_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u726 (
    .a(\rfxs[28] [10]),
    .b(\rfxs[29] [10]),
    .c(_al_u725_o),
    .d(i_rs1idx[1]),
    .o(_al_u726_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u727 (
    .a(\rfxs[26] [10]),
    .b(\rfxs[27] [10]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u727_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u728 (
    .a(\rfxs[24] [10]),
    .b(\rfxs[25] [10]),
    .c(_al_u727_o),
    .d(i_rs1idx[1]),
    .o(_al_u728_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u729 (
    .a(_al_u726_o),
    .b(_al_u728_o),
    .c(i_rs1idx[2]),
    .o(_al_u729_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u730 (
    .a(_al_u724_o),
    .b(_al_u729_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u730_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u731 (
    .a(n94),
    .b(_al_u730_o),
    .c(_al_u719_o),
    .d(i_rd_wdata[10]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[10]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u732 (
    .a(\rfxs[22] [1]),
    .b(\rfxs[23] [1]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u732_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u733 (
    .a(\rfxs[20] [1]),
    .b(\rfxs[21] [1]),
    .c(_al_u732_o),
    .d(i_rs1idx[1]),
    .o(_al_u733_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u734 (
    .a(\rfxs[17] [1]),
    .b(\rfxs[18] [1]),
    .c(\rfxs[19] [1]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u734_o));
  AL_MAP_LUT5 #(
    .EQN("((B*~(D*C))*~(A)*~(E)+(B*~(D*C))*A*~(E)+~((B*~(D*C)))*A*E+(B*~(D*C))*A*E)"),
    .INIT(32'haaaa0ccc))
    _al_u735 (
    .a(_al_u733_o),
    .b(_al_u734_o),
    .c(_al_u116_o),
    .d(\rfxs[16] [1]),
    .e(i_rs1idx[2]),
    .o(_al_u735_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u736 (
    .a(\rfxs[1] [1]),
    .b(\rfxs[2] [1]),
    .c(\rfxs[3] [1]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u736_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u737 (
    .a(\rfxs[5] [1]),
    .b(\rfxs[6] [1]),
    .c(\rfxs[7] [1]),
    .d(i_rs1idx[1]),
    .e(i_rs1idx[0]),
    .o(_al_u737_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u738 (
    .a(_al_u736_o),
    .b(_al_u737_o),
    .c(_al_u116_o),
    .d(\rfxs[4] [1]),
    .e(i_rs1idx[2]),
    .o(_al_u738_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u739 (
    .a(_al_u735_o),
    .b(_al_u738_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u739_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u740 (
    .a(\rfxs[8] [1]),
    .b(\rfxs[10] [1]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u740_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u741 (
    .a(\rfxs[11] [1]),
    .b(\rfxs[9] [1]),
    .c(_al_u740_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b1/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u742 (
    .a(\rfxs[14] [1]),
    .b(\rfxs[15] [1]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u742_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u743 (
    .a(\rfxs[12] [1]),
    .b(\rfxs[13] [1]),
    .c(_al_u742_o),
    .d(i_rs1idx[1]),
    .o(_al_u743_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u744 (
    .a(\mux31_b1/B1_2 ),
    .b(_al_u743_o),
    .c(i_rs1idx[2]),
    .o(_al_u744_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u745 (
    .a(\rfxs[30] [1]),
    .b(\rfxs[31] [1]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u745_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u746 (
    .a(\rfxs[28] [1]),
    .b(\rfxs[29] [1]),
    .c(_al_u745_o),
    .d(i_rs1idx[1]),
    .o(_al_u746_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u747 (
    .a(\rfxs[26] [1]),
    .b(\rfxs[27] [1]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u747_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u748 (
    .a(\rfxs[24] [1]),
    .b(\rfxs[25] [1]),
    .c(_al_u747_o),
    .d(i_rs1idx[1]),
    .o(_al_u748_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u749 (
    .a(_al_u746_o),
    .b(_al_u748_o),
    .c(i_rs1idx[2]),
    .o(_al_u749_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u75 (
    .a(i_rdidx[0]),
    .b(i_rdwen),
    .o(_al_u75_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u750 (
    .a(_al_u744_o),
    .b(_al_u749_o),
    .c(i_rs1idx[4]),
    .d(i_rs1idx[3]),
    .o(_al_u750_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u751 (
    .a(n94),
    .b(_al_u750_o),
    .c(_al_u739_o),
    .d(i_rd_wdata[1]),
    .e(i_rs1ren),
    .o(o_rs1_rdata[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u752 (
    .a(\rfxs[26] [0]),
    .b(\rfxs[27] [0]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u752_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u753 (
    .a(\rfxs[24] [0]),
    .b(\rfxs[25] [0]),
    .c(_al_u752_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b0/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u754 (
    .a(\rfxs[30] [0]),
    .b(\rfxs[31] [0]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u754_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u755 (
    .a(\rfxs[28] [0]),
    .b(\rfxs[29] [0]),
    .c(_al_u754_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b0/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u756 (
    .a(\mux31_b0/B1_6 ),
    .b(\mux31_b0/B1_7 ),
    .c(i_rs1idx[2]),
    .d(i_rs1idx[3]),
    .o(_al_u756_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u757 (
    .a(\mux31_b0/B1_4 ),
    .b(\mux31_b0/B1_5 ),
    .c(_al_u756_o),
    .d(i_rs1idx[3]),
    .o(\mux31_b0/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u758 (
    .a(\rfxs[14] [0]),
    .b(\rfxs[15] [0]),
    .c(i_rs1idx[0]),
    .d(i_rs1idx[1]),
    .o(_al_u758_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u759 (
    .a(\rfxs[12] [0]),
    .b(\rfxs[13] [0]),
    .c(_al_u758_o),
    .d(i_rs1idx[1]),
    .o(\mux31_b0/B1_3 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*~B*A)"),
    .INIT(32'h00000200))
    _al_u76 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n10));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u760 (
    .a(\rfxs[8] [0]),
    .b(\rfxs[10] [0]),
    .c(i_rs1idx[1]),
    .d(i_rs1idx[0]),
    .o(_al_u760_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u761 (
    .a(\rfxs[11] [0]),
    .b(\rfxs[9] [0]),
    .c(_al_u760_o),
    .d(i_rs1idx[0]),
    .o(\mux31_b0/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u762 (
    .a(\mux31_b0/B1_1 ),
    .b(\mux31_b0/B1_2 ),
    .c(_al_u224_o),
    .d(i_rs1idx[3]),
    .e(i_rs1idx[2]),
    .o(_al_u762_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u763 (
    .a(\mux31_b0/B3_1 ),
    .b(_al_u762_o),
    .c(\mux31_b0/B1_3 ),
    .d(_al_u227_o),
    .e(i_rs1idx[4]),
    .o(_al_u763_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u764 (
    .a(n94),
    .b(_al_u763_o),
    .c(i_rd_wdata[0]),
    .d(i_rs1ren),
    .o(o_rs1_rdata[0]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u765 (
    .a(i_rdidx[4]),
    .b(i_rdidx[3]),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u765_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u766 (
    .a(i_rdidx[1]),
    .b(i_rdidx[0]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u766_o));
  AL_MAP_LUT5 #(
    .EQN("(D*B*A*~(E@C))"),
    .INIT(32'h80000800))
    _al_u767 (
    .a(_al_u765_o),
    .b(_al_u766_o),
    .c(i_rdidx[2]),
    .d(i_rdwen),
    .e(i_rs2idx[2]),
    .o(n98));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u768 (
    .a(\rfxs[6] [8]),
    .b(\rfxs[7] [8]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u768_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u769 (
    .a(\rfxs[14] [8]),
    .b(\rfxs[15] [8]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u769_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*A)"),
    .INIT(32'h02000000))
    _al_u77 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n16));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u770 (
    .a(\rfxs[6] [5]),
    .b(\rfxs[7] [5]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u770_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u771 (
    .a(\rfxs[14] [5]),
    .b(\rfxs[15] [5]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u771_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u772 (
    .a(\rfxs[6] [29]),
    .b(\rfxs[7] [29]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u772_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u773 (
    .a(\rfxs[14] [29]),
    .b(\rfxs[15] [29]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u773_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u774 (
    .a(\rfxs[6] [23]),
    .b(\rfxs[7] [23]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u774_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hcfa0))
    _al_u775 (
    .a(\rfxs[14] [23]),
    .b(\rfxs[15] [23]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u775_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u776 (
    .a(i_rs2idx[1]),
    .b(i_rs2idx[0]),
    .o(_al_u776_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u777 (
    .a(\rfxs[18] [9]),
    .b(\rfxs[19] [9]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u777_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u778 (
    .a(\rfxs[16] [9]),
    .b(\rfxs[17] [9]),
    .c(_al_u777_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b9/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u779 (
    .a(\rfxs[22] [9]),
    .b(\rfxs[23] [9]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u779_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    _al_u78 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n4));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u780 (
    .a(\rfxs[20] [9]),
    .b(\rfxs[21] [9]),
    .c(_al_u779_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b9/B1_5 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u781 (
    .a(\rfxs[26] [9]),
    .b(\rfxs[27] [9]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u781_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u782 (
    .a(\rfxs[24] [9]),
    .b(\rfxs[25] [9]),
    .c(_al_u781_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b9/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u783 (
    .a(\rfxs[30] [9]),
    .b(\rfxs[31] [9]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u783_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u784 (
    .a(\rfxs[28] [9]),
    .b(\rfxs[29] [9]),
    .c(_al_u783_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b9/B1_7 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u785 (
    .a(\rfxs[1] [9]),
    .b(\rfxs[2] [9]),
    .c(\rfxs[3] [9]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u785_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u786 (
    .a(\rfxs[6] [9]),
    .b(\rfxs[7] [9]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u786_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u787 (
    .a(\rfxs[4] [9]),
    .b(\rfxs[5] [9]),
    .c(_al_u786_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b9/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u788 (
    .a(\rfxs[18] [7]),
    .b(\rfxs[19] [7]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u788_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u789 (
    .a(\rfxs[16] [7]),
    .b(\rfxs[17] [7]),
    .c(_al_u788_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b7/B1_4 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u79 (
    .a(i_rdidx[0]),
    .b(i_rdwen),
    .o(_al_u79_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u790 (
    .a(\rfxs[22] [7]),
    .b(\rfxs[23] [7]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u790_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u791 (
    .a(\rfxs[20] [7]),
    .b(\rfxs[21] [7]),
    .c(_al_u790_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b7/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u792 (
    .a(\rfxs[1] [7]),
    .b(\rfxs[2] [7]),
    .c(\rfxs[3] [7]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u792_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u793 (
    .a(\rfxs[6] [7]),
    .b(\rfxs[7] [7]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u793_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u794 (
    .a(\rfxs[4] [7]),
    .b(\rfxs[5] [7]),
    .c(_al_u793_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b7/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u795 (
    .a(\rfxs[18] [6]),
    .b(\rfxs[19] [6]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u795_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u796 (
    .a(\rfxs[16] [6]),
    .b(\rfxs[17] [6]),
    .c(_al_u795_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b6/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u797 (
    .a(\rfxs[22] [6]),
    .b(\rfxs[23] [6]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u797_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u798 (
    .a(\rfxs[20] [6]),
    .b(\rfxs[21] [6]),
    .c(_al_u797_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b6/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u799 (
    .a(\rfxs[1] [6]),
    .b(\rfxs[2] [6]),
    .c(\rfxs[3] [6]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u799_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*~B*A)"),
    .INIT(32'h02000000))
    _al_u80 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n19));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u800 (
    .a(\rfxs[6] [6]),
    .b(\rfxs[7] [6]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u800_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u801 (
    .a(\rfxs[4] [6]),
    .b(\rfxs[5] [6]),
    .c(_al_u800_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b6/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u802 (
    .a(\rfxs[18] [31]),
    .b(\rfxs[19] [31]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u802_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u803 (
    .a(\rfxs[16] [31]),
    .b(\rfxs[17] [31]),
    .c(_al_u802_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b31/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u804 (
    .a(\rfxs[22] [31]),
    .b(\rfxs[23] [31]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u804_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u805 (
    .a(\rfxs[20] [31]),
    .b(\rfxs[21] [31]),
    .c(_al_u804_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b31/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u806 (
    .a(\rfxs[1] [31]),
    .b(\rfxs[2] [31]),
    .c(\rfxs[3] [31]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u806_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u807 (
    .a(\rfxs[6] [31]),
    .b(\rfxs[7] [31]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u807_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u808 (
    .a(\rfxs[4] [31]),
    .b(\rfxs[5] [31]),
    .c(_al_u807_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b31/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u809 (
    .a(\rfxs[18] [30]),
    .b(\rfxs[19] [30]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u809_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    _al_u81 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n7));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u810 (
    .a(\rfxs[16] [30]),
    .b(\rfxs[17] [30]),
    .c(_al_u809_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b30/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u811 (
    .a(\rfxs[22] [30]),
    .b(\rfxs[23] [30]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u811_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u812 (
    .a(\rfxs[20] [30]),
    .b(\rfxs[21] [30]),
    .c(_al_u811_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b30/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u813 (
    .a(\rfxs[1] [30]),
    .b(\rfxs[2] [30]),
    .c(\rfxs[3] [30]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u813_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u814 (
    .a(\rfxs[6] [30]),
    .b(\rfxs[7] [30]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u814_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u815 (
    .a(\rfxs[4] [30]),
    .b(\rfxs[5] [30]),
    .c(_al_u814_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b30/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u816 (
    .a(\rfxs[18] [28]),
    .b(\rfxs[19] [28]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u816_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u817 (
    .a(\rfxs[16] [28]),
    .b(\rfxs[17] [28]),
    .c(_al_u816_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b28/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u818 (
    .a(\rfxs[22] [28]),
    .b(\rfxs[23] [28]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u818_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u819 (
    .a(\rfxs[20] [28]),
    .b(\rfxs[21] [28]),
    .c(_al_u818_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b28/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*~B*A)"),
    .INIT(32'h00000200))
    _al_u82 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n13));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u820 (
    .a(\rfxs[1] [28]),
    .b(\rfxs[2] [28]),
    .c(\rfxs[3] [28]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u820_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u821 (
    .a(\rfxs[6] [28]),
    .b(\rfxs[7] [28]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u821_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u822 (
    .a(\rfxs[4] [28]),
    .b(\rfxs[5] [28]),
    .c(_al_u821_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b28/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u823 (
    .a(\rfxs[18] [27]),
    .b(\rfxs[19] [27]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u823_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u824 (
    .a(\rfxs[16] [27]),
    .b(\rfxs[17] [27]),
    .c(_al_u823_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b27/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u825 (
    .a(\rfxs[22] [27]),
    .b(\rfxs[23] [27]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u825_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u826 (
    .a(\rfxs[20] [27]),
    .b(\rfxs[21] [27]),
    .c(_al_u825_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b27/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u827 (
    .a(\rfxs[1] [27]),
    .b(\rfxs[2] [27]),
    .c(\rfxs[3] [27]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u827_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u828 (
    .a(\rfxs[6] [27]),
    .b(\rfxs[7] [27]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u828_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u829 (
    .a(\rfxs[4] [27]),
    .b(\rfxs[5] [27]),
    .c(_al_u828_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b27/B1_1 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u83 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n1));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u830 (
    .a(\rfxs[18] [25]),
    .b(\rfxs[19] [25]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u830_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u831 (
    .a(\rfxs[16] [25]),
    .b(\rfxs[17] [25]),
    .c(_al_u830_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b25/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u832 (
    .a(\rfxs[22] [25]),
    .b(\rfxs[23] [25]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u832_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u833 (
    .a(\rfxs[20] [25]),
    .b(\rfxs[21] [25]),
    .c(_al_u832_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b25/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u834 (
    .a(\rfxs[1] [25]),
    .b(\rfxs[2] [25]),
    .c(\rfxs[3] [25]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u834_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u835 (
    .a(\rfxs[6] [25]),
    .b(\rfxs[7] [25]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u835_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u836 (
    .a(\rfxs[4] [25]),
    .b(\rfxs[5] [25]),
    .c(_al_u835_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b25/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u837 (
    .a(\rfxs[18] [24]),
    .b(\rfxs[19] [24]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u837_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u838 (
    .a(\rfxs[16] [24]),
    .b(\rfxs[17] [24]),
    .c(_al_u837_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b24/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u839 (
    .a(\rfxs[22] [24]),
    .b(\rfxs[23] [24]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u839_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*B*A)"),
    .INIT(32'h08000000))
    _al_u84 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n67));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u840 (
    .a(\rfxs[20] [24]),
    .b(\rfxs[21] [24]),
    .c(_al_u839_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b24/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u841 (
    .a(\rfxs[1] [24]),
    .b(\rfxs[2] [24]),
    .c(\rfxs[3] [24]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u841_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u842 (
    .a(\rfxs[6] [24]),
    .b(\rfxs[7] [24]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u842_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u843 (
    .a(\rfxs[4] [24]),
    .b(\rfxs[5] [24]),
    .c(_al_u842_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b24/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u844 (
    .a(\rfxs[18] [22]),
    .b(\rfxs[19] [22]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u844_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u845 (
    .a(\rfxs[16] [22]),
    .b(\rfxs[17] [22]),
    .c(_al_u844_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b22/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u846 (
    .a(\rfxs[22] [22]),
    .b(\rfxs[23] [22]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u846_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u847 (
    .a(\rfxs[20] [22]),
    .b(\rfxs[21] [22]),
    .c(_al_u846_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b22/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u848 (
    .a(\rfxs[1] [22]),
    .b(\rfxs[2] [22]),
    .c(\rfxs[3] [22]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u848_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u849 (
    .a(\rfxs[6] [22]),
    .b(\rfxs[7] [22]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u849_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*B*A)"),
    .INIT(32'h08000000))
    _al_u85 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n64));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u850 (
    .a(\rfxs[4] [22]),
    .b(\rfxs[5] [22]),
    .c(_al_u849_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b22/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u851 (
    .a(\rfxs[18] [18]),
    .b(\rfxs[19] [18]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u851_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u852 (
    .a(\rfxs[16] [18]),
    .b(\rfxs[17] [18]),
    .c(_al_u851_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b18/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u853 (
    .a(\rfxs[22] [18]),
    .b(\rfxs[23] [18]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u853_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u854 (
    .a(\rfxs[20] [18]),
    .b(\rfxs[21] [18]),
    .c(_al_u853_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b18/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u855 (
    .a(\rfxs[1] [18]),
    .b(\rfxs[2] [18]),
    .c(\rfxs[3] [18]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u855_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u856 (
    .a(\rfxs[6] [18]),
    .b(\rfxs[7] [18]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u856_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u857 (
    .a(\rfxs[4] [18]),
    .b(\rfxs[5] [18]),
    .c(_al_u856_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b18/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u858 (
    .a(\rfxs[18] [17]),
    .b(\rfxs[19] [17]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u858_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u859 (
    .a(\rfxs[16] [17]),
    .b(\rfxs[17] [17]),
    .c(_al_u858_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b17/B1_4 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    _al_u86 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n61));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u860 (
    .a(\rfxs[22] [17]),
    .b(\rfxs[23] [17]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u860_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u861 (
    .a(\rfxs[20] [17]),
    .b(\rfxs[21] [17]),
    .c(_al_u860_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b17/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u862 (
    .a(\rfxs[1] [17]),
    .b(\rfxs[2] [17]),
    .c(\rfxs[3] [17]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u862_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u863 (
    .a(\rfxs[6] [17]),
    .b(\rfxs[7] [17]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u863_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u864 (
    .a(\rfxs[4] [17]),
    .b(\rfxs[5] [17]),
    .c(_al_u863_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b17/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u865 (
    .a(\rfxs[18] [15]),
    .b(\rfxs[19] [15]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u865_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u866 (
    .a(\rfxs[16] [15]),
    .b(\rfxs[17] [15]),
    .c(_al_u865_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b15/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u867 (
    .a(\rfxs[22] [15]),
    .b(\rfxs[23] [15]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u867_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u868 (
    .a(\rfxs[20] [15]),
    .b(\rfxs[21] [15]),
    .c(_al_u867_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b15/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u869 (
    .a(\rfxs[1] [15]),
    .b(\rfxs[2] [15]),
    .c(\rfxs[3] [15]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u869_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    _al_u87 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n58));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u870 (
    .a(\rfxs[6] [15]),
    .b(\rfxs[7] [15]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u870_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u871 (
    .a(\rfxs[4] [15]),
    .b(\rfxs[5] [15]),
    .c(_al_u870_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b15/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u872 (
    .a(\rfxs[18] [14]),
    .b(\rfxs[19] [14]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u872_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u873 (
    .a(\rfxs[16] [14]),
    .b(\rfxs[17] [14]),
    .c(_al_u872_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b14/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u874 (
    .a(\rfxs[22] [14]),
    .b(\rfxs[23] [14]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u874_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u875 (
    .a(\rfxs[20] [14]),
    .b(\rfxs[21] [14]),
    .c(_al_u874_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b14/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u876 (
    .a(\rfxs[1] [14]),
    .b(\rfxs[2] [14]),
    .c(\rfxs[3] [14]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u876_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u877 (
    .a(\rfxs[6] [14]),
    .b(\rfxs[7] [14]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u877_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u878 (
    .a(\rfxs[4] [14]),
    .b(\rfxs[5] [14]),
    .c(_al_u877_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b14/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u879 (
    .a(\rfxs[18] [13]),
    .b(\rfxs[19] [13]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u879_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'h00080000))
    _al_u88 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n55));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u880 (
    .a(\rfxs[16] [13]),
    .b(\rfxs[17] [13]),
    .c(_al_u879_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b13/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u881 (
    .a(\rfxs[22] [13]),
    .b(\rfxs[23] [13]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u881_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u882 (
    .a(\rfxs[20] [13]),
    .b(\rfxs[21] [13]),
    .c(_al_u881_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b13/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u883 (
    .a(\rfxs[1] [13]),
    .b(\rfxs[2] [13]),
    .c(\rfxs[3] [13]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u883_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u884 (
    .a(\rfxs[6] [13]),
    .b(\rfxs[7] [13]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u884_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u885 (
    .a(\rfxs[4] [13]),
    .b(\rfxs[5] [13]),
    .c(_al_u884_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b13/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u886 (
    .a(\rfxs[18] [12]),
    .b(\rfxs[19] [12]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u886_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u887 (
    .a(\rfxs[16] [12]),
    .b(\rfxs[17] [12]),
    .c(_al_u886_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b12/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u888 (
    .a(\rfxs[22] [12]),
    .b(\rfxs[23] [12]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u888_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u889 (
    .a(\rfxs[20] [12]),
    .b(\rfxs[21] [12]),
    .c(_al_u888_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b12/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'h00080000))
    _al_u89 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n52));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u890 (
    .a(\rfxs[1] [12]),
    .b(\rfxs[2] [12]),
    .c(\rfxs[3] [12]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u890_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u891 (
    .a(\rfxs[6] [12]),
    .b(\rfxs[7] [12]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u891_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u892 (
    .a(\rfxs[4] [12]),
    .b(\rfxs[5] [12]),
    .c(_al_u891_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b12/B1_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u893 (
    .a(\rfxs[18] [0]),
    .b(\rfxs[19] [0]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u893_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u894 (
    .a(\rfxs[16] [0]),
    .b(\rfxs[17] [0]),
    .c(_al_u893_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b0/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u895 (
    .a(\rfxs[22] [0]),
    .b(\rfxs[23] [0]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u895_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u896 (
    .a(\rfxs[20] [0]),
    .b(\rfxs[21] [0]),
    .c(_al_u895_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b0/B1_5 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u897 (
    .a(\rfxs[1] [0]),
    .b(\rfxs[2] [0]),
    .c(\rfxs[3] [0]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u897_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u898 (
    .a(\rfxs[6] [0]),
    .b(\rfxs[7] [0]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u898_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u899 (
    .a(\rfxs[4] [0]),
    .b(\rfxs[5] [0]),
    .c(_al_u898_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b0/B1_1 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    _al_u90 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n49));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u900 (
    .a(i_rs2idx[3]),
    .b(i_rs2idx[2]),
    .o(_al_u900_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u901 (
    .a(\mux34_b9/B1_6 ),
    .b(\mux34_b9/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u901_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u902 (
    .a(\mux34_b9/B1_4 ),
    .b(\mux34_b9/B1_5 ),
    .c(_al_u901_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b9/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u903 (
    .a(\rfxs[14] [9]),
    .b(\rfxs[15] [9]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u903_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u904 (
    .a(\rfxs[12] [9]),
    .b(\rfxs[13] [9]),
    .c(_al_u903_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b9/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u905 (
    .a(\rfxs[8] [9]),
    .b(\rfxs[10] [9]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u905_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u906 (
    .a(\rfxs[11] [9]),
    .b(\rfxs[9] [9]),
    .c(_al_u905_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b9/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u907 (
    .a(\mux34_b9/B1_1 ),
    .b(\mux34_b9/B1_2 ),
    .c(_al_u785_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u907_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u908 (
    .a(\mux34_b9/B3_1 ),
    .b(_al_u907_o),
    .c(\mux34_b9/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u908_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u909 (
    .a(n98),
    .b(_al_u908_o),
    .c(i_rd_wdata[9]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[9]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    _al_u91 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n46));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u910 (
    .a(\rfxs[26] [8]),
    .b(\rfxs[27] [8]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u910_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u911 (
    .a(\rfxs[24] [8]),
    .b(\rfxs[25] [8]),
    .c(_al_u910_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b8/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u912 (
    .a(\rfxs[30] [8]),
    .b(\rfxs[31] [8]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u912_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u913 (
    .a(\rfxs[28] [8]),
    .b(\rfxs[29] [8]),
    .c(_al_u912_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b8/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u914 (
    .a(\rfxs[18] [8]),
    .b(\rfxs[19] [8]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u914_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u915 (
    .a(\rfxs[16] [8]),
    .b(\rfxs[17] [8]),
    .c(_al_u914_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b8/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u916 (
    .a(\rfxs[22] [8]),
    .b(\rfxs[23] [8]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u916_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u917 (
    .a(\rfxs[20] [8]),
    .b(\rfxs[21] [8]),
    .c(_al_u916_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b8/B1_5 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fca))
    _al_u918 (
    .a(\mux34_b8/B1_4 ),
    .b(\mux34_b8/B1_5 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u918_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u919 (
    .a(\mux34_b8/B1_6 ),
    .b(\mux34_b8/B1_7 ),
    .c(_al_u918_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b8/B3_1 ));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u92 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n91));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u920 (
    .a(\mux34_b8/B3_1 ),
    .b(i_rs2idx[4]),
    .o(_al_u920_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u921 (
    .a(\rfxs[8] [8]),
    .b(\rfxs[10] [8]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u921_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u922 (
    .a(\rfxs[11] [8]),
    .b(\rfxs[9] [8]),
    .c(_al_u921_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b8/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u923 (
    .a(\rfxs[1] [8]),
    .b(\rfxs[2] [8]),
    .c(\rfxs[3] [8]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u923_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h005c))
    _al_u924 (
    .a(\mux34_b8/B1_2 ),
    .b(_al_u923_o),
    .c(i_rs2idx[3]),
    .d(i_rs2idx[2]),
    .o(_al_u924_o));
  AL_MAP_LUT5 #(
    .EQN("(D*(~(A)*B*~(C)*~(E)+A*~(B)*C*~(E)+~(A)*B*C*~(E)+A*B*C*~(E)+A*~(B)*~(C)*E+A*B*~(C)*E+A*~(B)*C*E+A*B*C*E))"),
    .INIT(32'haa00e400))
    _al_u925 (
    .a(_al_u769_o),
    .b(\rfxs[12] [8]),
    .c(\rfxs[13] [8]),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[1]),
    .o(_al_u925_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*(~(A)*B*~(C)*~(E)+A*~(B)*C*~(E)+~(A)*B*C*~(E)+A*B*C*~(E)+A*~(B)*~(C)*E+A*B*~(C)*E+A*~(B)*C*E+A*B*C*E))"),
    .INIT(32'h00aa00e4))
    _al_u926 (
    .a(_al_u768_o),
    .b(\rfxs[4] [8]),
    .c(\rfxs[5] [8]),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[1]),
    .o(_al_u926_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~A*~(E*~C*~B)))"),
    .INIT(32'h00ab00aa))
    _al_u927 (
    .a(_al_u924_o),
    .b(_al_u925_o),
    .c(_al_u926_o),
    .d(i_rs2idx[4]),
    .e(i_rs2idx[2]),
    .o(_al_u927_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u928 (
    .a(n98),
    .b(_al_u920_o),
    .c(_al_u927_o),
    .d(i_rd_wdata[8]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[8]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u929 (
    .a(\rfxs[26] [7]),
    .b(\rfxs[27] [7]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u929_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u93 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n88));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u930 (
    .a(\rfxs[24] [7]),
    .b(\rfxs[25] [7]),
    .c(_al_u929_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b7/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u931 (
    .a(\rfxs[30] [7]),
    .b(\rfxs[31] [7]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u931_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u932 (
    .a(\rfxs[28] [7]),
    .b(\rfxs[29] [7]),
    .c(_al_u931_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b7/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u933 (
    .a(\mux34_b7/B1_6 ),
    .b(\mux34_b7/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u933_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u934 (
    .a(\mux34_b7/B1_4 ),
    .b(\mux34_b7/B1_5 ),
    .c(_al_u933_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b7/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u935 (
    .a(\rfxs[14] [7]),
    .b(\rfxs[15] [7]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u935_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u936 (
    .a(\rfxs[12] [7]),
    .b(\rfxs[13] [7]),
    .c(_al_u935_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b7/B1_3 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u937 (
    .a(\rfxs[8] [7]),
    .b(\rfxs[10] [7]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u937_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u938 (
    .a(\rfxs[11] [7]),
    .b(\rfxs[9] [7]),
    .c(_al_u937_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b7/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u939 (
    .a(\mux34_b7/B1_1 ),
    .b(\mux34_b7/B1_2 ),
    .c(_al_u792_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u939_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    _al_u94 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n85));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u940 (
    .a(\mux34_b7/B3_1 ),
    .b(_al_u939_o),
    .c(\mux34_b7/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u940_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u941 (
    .a(n98),
    .b(_al_u940_o),
    .c(i_rd_wdata[7]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[7]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u942 (
    .a(\rfxs[26] [6]),
    .b(\rfxs[27] [6]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u942_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u943 (
    .a(\rfxs[24] [6]),
    .b(\rfxs[25] [6]),
    .c(_al_u942_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b6/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u944 (
    .a(\rfxs[30] [6]),
    .b(\rfxs[31] [6]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u944_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u945 (
    .a(\rfxs[28] [6]),
    .b(\rfxs[29] [6]),
    .c(_al_u944_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b6/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u946 (
    .a(\mux34_b6/B1_6 ),
    .b(\mux34_b6/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u946_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u947 (
    .a(\mux34_b6/B1_4 ),
    .b(\mux34_b6/B1_5 ),
    .c(_al_u946_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b6/B3_1 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u948 (
    .a(\rfxs[14] [6]),
    .b(\rfxs[15] [6]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u948_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u949 (
    .a(\rfxs[12] [6]),
    .b(\rfxs[13] [6]),
    .c(_al_u948_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b6/B1_3 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*C*B*A)"),
    .INIT(32'h00008000))
    _al_u95 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n82));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u950 (
    .a(\rfxs[8] [6]),
    .b(\rfxs[10] [6]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u950_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u951 (
    .a(\rfxs[11] [6]),
    .b(\rfxs[9] [6]),
    .c(_al_u950_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b6/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hff5533f0))
    _al_u952 (
    .a(\mux34_b6/B1_1 ),
    .b(\mux34_b6/B1_2 ),
    .c(_al_u799_o),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[2]),
    .o(_al_u952_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(B*~(D*C))*~(A)*~(E)+~(B*~(D*C))*A*~(E)+~(~(B*~(D*C)))*A*E+~(B*~(D*C))*A*E)"),
    .INIT(32'h55550ccc))
    _al_u953 (
    .a(\mux34_b6/B3_1 ),
    .b(_al_u952_o),
    .c(\mux34_b6/B1_3 ),
    .d(_al_u900_o),
    .e(i_rs2idx[4]),
    .o(_al_u953_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A))"),
    .INIT(16'hb100))
    _al_u954 (
    .a(n98),
    .b(_al_u953_o),
    .c(i_rd_wdata[6]),
    .d(i_rs2ren),
    .o(o_rs2_rdata[6]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u955 (
    .a(\rfxs[26] [5]),
    .b(\rfxs[27] [5]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u955_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u956 (
    .a(\rfxs[24] [5]),
    .b(\rfxs[25] [5]),
    .c(_al_u955_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b5/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u957 (
    .a(\rfxs[30] [5]),
    .b(\rfxs[31] [5]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u957_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u958 (
    .a(\rfxs[28] [5]),
    .b(\rfxs[29] [5]),
    .c(_al_u957_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b5/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u959 (
    .a(\rfxs[18] [5]),
    .b(\rfxs[19] [5]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u959_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*A)"),
    .INIT(32'h00800000))
    _al_u96 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n79));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u960 (
    .a(\rfxs[16] [5]),
    .b(\rfxs[17] [5]),
    .c(_al_u959_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b5/B1_4 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u961 (
    .a(\rfxs[22] [5]),
    .b(\rfxs[23] [5]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u961_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u962 (
    .a(\rfxs[20] [5]),
    .b(\rfxs[21] [5]),
    .c(_al_u961_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b5/B1_5 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fca))
    _al_u963 (
    .a(\mux34_b5/B1_4 ),
    .b(\mux34_b5/B1_5 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u963_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u964 (
    .a(\mux34_b5/B1_6 ),
    .b(\mux34_b5/B1_7 ),
    .c(_al_u963_o),
    .d(i_rs2idx[3]),
    .o(\mux34_b5/B3_1 ));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u965 (
    .a(\mux34_b5/B3_1 ),
    .b(i_rs2idx[4]),
    .o(_al_u965_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u966 (
    .a(\rfxs[8] [5]),
    .b(\rfxs[10] [5]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u966_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u967 (
    .a(\rfxs[11] [5]),
    .b(\rfxs[9] [5]),
    .c(_al_u966_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b5/B1_2 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u968 (
    .a(\rfxs[1] [5]),
    .b(\rfxs[2] [5]),
    .c(\rfxs[3] [5]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u968_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h005c))
    _al_u969 (
    .a(\mux34_b5/B1_2 ),
    .b(_al_u968_o),
    .c(i_rs2idx[3]),
    .d(i_rs2idx[2]),
    .o(_al_u969_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*A)"),
    .INIT(32'h00800000))
    _al_u97 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n76));
  AL_MAP_LUT5 #(
    .EQN("(D*(~(A)*B*~(C)*~(E)+A*~(B)*C*~(E)+~(A)*B*C*~(E)+A*B*C*~(E)+A*~(B)*~(C)*E+A*B*~(C)*E+A*~(B)*C*E+A*B*C*E))"),
    .INIT(32'haa00e400))
    _al_u970 (
    .a(_al_u771_o),
    .b(\rfxs[12] [5]),
    .c(\rfxs[13] [5]),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[1]),
    .o(_al_u970_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*(~(A)*B*~(C)*~(E)+A*~(B)*C*~(E)+~(A)*B*C*~(E)+A*B*C*~(E)+A*~(B)*~(C)*E+A*B*~(C)*E+A*~(B)*C*E+A*B*C*E))"),
    .INIT(32'h00aa00e4))
    _al_u971 (
    .a(_al_u770_o),
    .b(\rfxs[4] [5]),
    .c(\rfxs[5] [5]),
    .d(i_rs2idx[3]),
    .e(i_rs2idx[1]),
    .o(_al_u971_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~A*~(E*~C*~B)))"),
    .INIT(32'h00ab00aa))
    _al_u972 (
    .a(_al_u969_o),
    .b(_al_u970_o),
    .c(_al_u971_o),
    .d(i_rs2idx[4]),
    .e(i_rs2idx[2]),
    .o(_al_u972_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u973 (
    .a(n98),
    .b(_al_u965_o),
    .c(_al_u972_o),
    .d(i_rd_wdata[5]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[5]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u974 (
    .a(\rfxs[22] [4]),
    .b(\rfxs[23] [4]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u974_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u975 (
    .a(\rfxs[20] [4]),
    .b(\rfxs[21] [4]),
    .c(_al_u974_o),
    .d(i_rs2idx[1]),
    .o(_al_u975_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u976 (
    .a(\rfxs[18] [4]),
    .b(\rfxs[19] [4]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u976_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u977 (
    .a(\rfxs[16] [4]),
    .b(\rfxs[17] [4]),
    .c(_al_u976_o),
    .d(i_rs2idx[1]),
    .o(_al_u977_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u978 (
    .a(_al_u975_o),
    .b(_al_u977_o),
    .c(i_rs2idx[2]),
    .o(_al_u978_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u979 (
    .a(\rfxs[1] [4]),
    .b(\rfxs[2] [4]),
    .c(\rfxs[3] [4]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u979_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    _al_u98 (
    .a(_al_u79_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n73));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E)"),
    .INIT(32'h0f5533ff))
    _al_u980 (
    .a(\rfxs[5] [4]),
    .b(\rfxs[6] [4]),
    .c(\rfxs[7] [4]),
    .d(i_rs2idx[1]),
    .e(i_rs2idx[0]),
    .o(_al_u980_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~((B*~(D*C)))*~(E)+A*(B*~(D*C))*~(E)+~(A)*(B*~(D*C))*E+A*(B*~(D*C))*E)"),
    .INIT(32'h0cccaaaa))
    _al_u981 (
    .a(_al_u979_o),
    .b(_al_u980_o),
    .c(_al_u776_o),
    .d(\rfxs[4] [4]),
    .e(i_rs2idx[2]),
    .o(_al_u981_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u982 (
    .a(_al_u978_o),
    .b(_al_u981_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u982_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0f35))
    _al_u983 (
    .a(\rfxs[8] [4]),
    .b(\rfxs[10] [4]),
    .c(i_rs2idx[1]),
    .d(i_rs2idx[0]),
    .o(_al_u983_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u984 (
    .a(\rfxs[11] [4]),
    .b(\rfxs[9] [4]),
    .c(_al_u983_o),
    .d(i_rs2idx[0]),
    .o(\mux34_b4/B1_2 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u985 (
    .a(\rfxs[14] [4]),
    .b(\rfxs[15] [4]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u985_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u986 (
    .a(\rfxs[12] [4]),
    .b(\rfxs[13] [4]),
    .c(_al_u985_o),
    .d(i_rs2idx[1]),
    .o(_al_u986_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u987 (
    .a(\mux34_b4/B1_2 ),
    .b(_al_u986_o),
    .c(i_rs2idx[2]),
    .o(_al_u987_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u988 (
    .a(\rfxs[30] [4]),
    .b(\rfxs[31] [4]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u988_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u989 (
    .a(\rfxs[28] [4]),
    .b(\rfxs[29] [4]),
    .c(_al_u988_o),
    .d(i_rs2idx[1]),
    .o(_al_u989_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    _al_u99 (
    .a(_al_u75_o),
    .b(i_rdidx[4]),
    .c(i_rdidx[3]),
    .d(i_rdidx[2]),
    .e(i_rdidx[1]),
    .o(n70));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u990 (
    .a(\rfxs[26] [4]),
    .b(\rfxs[27] [4]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u990_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf053))
    _al_u991 (
    .a(\rfxs[24] [4]),
    .b(\rfxs[25] [4]),
    .c(_al_u990_o),
    .d(i_rs2idx[1]),
    .o(_al_u991_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u992 (
    .a(_al_u989_o),
    .b(_al_u991_o),
    .c(i_rs2idx[2]),
    .o(_al_u992_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C))"),
    .INIT(16'hca00))
    _al_u993 (
    .a(_al_u987_o),
    .b(_al_u992_o),
    .c(i_rs2idx[4]),
    .d(i_rs2idx[3]),
    .o(_al_u993_o));
  AL_MAP_LUT5 #(
    .EQN("(E*((~C*~B)*~(D)*~(A)+(~C*~B)*D*~(A)+~((~C*~B))*D*A+(~C*~B)*D*A))"),
    .INIT(32'hab010000))
    _al_u994 (
    .a(n98),
    .b(_al_u993_o),
    .c(_al_u982_o),
    .d(i_rd_wdata[4]),
    .e(i_rs2ren),
    .o(o_rs2_rdata[4]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u995 (
    .a(\rfxs[26] [31]),
    .b(\rfxs[27] [31]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u995_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u996 (
    .a(\rfxs[24] [31]),
    .b(\rfxs[25] [31]),
    .c(_al_u995_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b31/B1_6 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D)"),
    .INIT(16'h350f))
    _al_u997 (
    .a(\rfxs[30] [31]),
    .b(\rfxs[31] [31]),
    .c(i_rs2idx[0]),
    .d(i_rs2idx[1]),
    .o(_al_u997_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D)"),
    .INIT(16'h0fac))
    _al_u998 (
    .a(\rfxs[28] [31]),
    .b(\rfxs[29] [31]),
    .c(_al_u997_o),
    .d(i_rs2idx[1]),
    .o(\mux34_b31/B1_7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hca0f))
    _al_u999 (
    .a(\mux34_b31/B1_6 ),
    .b(\mux34_b31/B1_7 ),
    .c(i_rs2idx[2]),
    .d(i_rs2idx[3]),
    .o(_al_u999_o));
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b0 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[1] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b1 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[1] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b10 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[1] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b11 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[1] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b12 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[1] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b13 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[1] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b14 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[1] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b15 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[1] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b16 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[1] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b17 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[1] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b18 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[1] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b19 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[1] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b2 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[1] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b20 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[1] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b21 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[1] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b22 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[1] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b23 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[1] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b24 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[1] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b25 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[1] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b26 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[1] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b27 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[1] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b28 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[1] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b29 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[1] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b3 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[1] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b30 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[1] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b31 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[1] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b4 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[1] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b5 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[1] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b6 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[1] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b7 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[1] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b8 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[1] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b9 (
    .ce(n1),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[1] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b0 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[11] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b1 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[11] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b10 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[11] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b11 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[11] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b12 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[11] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b13 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[11] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b14 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[11] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b15 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[11] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b16 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[11] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b17 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[11] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b18 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[11] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b19 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[11] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b2 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[11] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b20 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[11] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b21 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[11] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b22 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[11] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b23 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[11] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b24 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[11] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b25 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[11] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b26 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[11] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b27 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[11] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b28 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[11] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b29 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[11] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b3 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[11] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b30 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[11] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b31 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[11] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b4 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[11] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b5 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[11] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b6 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[11] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b7 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[11] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b8 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[11] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg10_b9 (
    .ce(n31),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[11] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b0 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[12] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b1 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[12] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b10 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[12] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b11 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[12] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b12 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[12] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b13 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[12] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b14 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[12] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b15 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[12] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b16 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[12] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b17 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[12] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b18 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[12] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b19 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[12] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b2 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[12] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b20 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[12] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b21 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[12] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b22 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[12] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b23 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[12] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b24 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[12] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b25 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[12] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b26 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[12] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b27 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[12] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b28 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[12] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b29 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[12] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b3 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[12] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b30 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[12] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b31 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[12] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b4 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[12] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b5 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[12] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b6 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[12] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b7 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[12] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b8 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[12] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg11_b9 (
    .ce(n34),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[12] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b0 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[13] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b1 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[13] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b10 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[13] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b11 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[13] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b12 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[13] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b13 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[13] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b14 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[13] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b15 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[13] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b16 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[13] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b17 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[13] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b18 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[13] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b19 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[13] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b2 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[13] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b20 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[13] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b21 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[13] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b22 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[13] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b23 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[13] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b24 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[13] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b25 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[13] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b26 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[13] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b27 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[13] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b28 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[13] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b29 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[13] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b3 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[13] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b30 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[13] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b31 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[13] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b4 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[13] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b5 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[13] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b6 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[13] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b7 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[13] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b8 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[13] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg12_b9 (
    .ce(n37),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[13] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b0 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[14] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b1 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[14] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b10 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[14] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b11 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[14] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b12 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[14] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b13 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[14] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b14 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[14] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b15 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[14] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b16 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[14] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b17 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[14] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b18 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[14] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b19 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[14] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b2 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[14] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b20 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[14] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b21 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[14] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b22 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[14] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b23 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[14] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b24 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[14] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b25 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[14] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b26 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[14] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b27 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[14] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b28 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[14] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b29 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[14] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b3 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[14] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b30 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[14] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b31 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[14] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b4 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[14] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b5 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[14] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b6 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[14] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b7 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[14] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b8 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[14] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg13_b9 (
    .ce(n40),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[14] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b0 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[15] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b1 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[15] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b10 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[15] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b11 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[15] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b12 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[15] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b13 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[15] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b14 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[15] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b15 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[15] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b16 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[15] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b17 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[15] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b18 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[15] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b19 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[15] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b2 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[15] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b20 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[15] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b21 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[15] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b22 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[15] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b23 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[15] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b24 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[15] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b25 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[15] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b26 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[15] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b27 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[15] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b28 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[15] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b29 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[15] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b3 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[15] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b30 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[15] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b31 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[15] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b4 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[15] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b5 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[15] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b6 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[15] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b7 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[15] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b8 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[15] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg14_b9 (
    .ce(n43),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[15] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b0 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[16] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b1 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[16] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b10 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[16] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b11 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[16] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b12 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[16] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b13 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[16] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b14 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[16] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b15 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[16] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b16 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[16] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b17 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[16] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b18 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[16] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b19 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[16] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b2 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[16] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b20 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[16] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b21 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[16] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b22 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[16] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b23 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[16] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b24 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[16] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b25 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[16] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b26 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[16] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b27 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[16] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b28 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[16] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b29 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[16] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b3 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[16] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b30 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[16] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b31 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[16] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b4 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[16] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b5 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[16] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b6 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[16] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b7 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[16] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b8 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[16] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg15_b9 (
    .ce(n46),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[16] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b0 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[17] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b1 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[17] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b10 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[17] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b11 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[17] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b12 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[17] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b13 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[17] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b14 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[17] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b15 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[17] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b16 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[17] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b17 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[17] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b18 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[17] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b19 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[17] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b2 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[17] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b20 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[17] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b21 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[17] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b22 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[17] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b23 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[17] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b24 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[17] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b25 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[17] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b26 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[17] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b27 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[17] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b28 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[17] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b29 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[17] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b3 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[17] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b30 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[17] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b31 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[17] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b4 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[17] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b5 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[17] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b6 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[17] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b7 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[17] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b8 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[17] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg16_b9 (
    .ce(n49),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[17] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b0 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[18] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b1 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[18] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b10 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[18] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b11 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[18] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b12 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[18] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b13 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[18] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b14 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[18] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b15 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[18] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b16 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[18] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b17 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[18] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b18 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[18] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b19 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[18] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b2 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[18] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b20 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[18] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b21 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[18] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b22 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[18] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b23 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[18] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b24 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[18] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b25 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[18] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b26 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[18] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b27 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[18] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b28 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[18] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b29 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[18] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b3 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[18] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b30 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[18] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b31 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[18] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b4 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[18] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b5 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[18] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b6 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[18] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b7 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[18] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b8 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[18] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg17_b9 (
    .ce(n52),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[18] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b0 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[19] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b1 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[19] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b10 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[19] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b11 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[19] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b12 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[19] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b13 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[19] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b14 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[19] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b15 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[19] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b16 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[19] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b17 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[19] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b18 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[19] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b19 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[19] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b2 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[19] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b20 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[19] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b21 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[19] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b22 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[19] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b23 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[19] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b24 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[19] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b25 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[19] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b26 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[19] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b27 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[19] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b28 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[19] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b29 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[19] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b3 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[19] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b30 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[19] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b31 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[19] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b4 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[19] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b5 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[19] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b6 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[19] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b7 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[19] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b8 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[19] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg18_b9 (
    .ce(n55),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[19] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b0 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[20] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b1 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[20] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b10 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[20] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b11 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[20] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b12 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[20] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b13 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[20] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b14 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[20] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b15 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[20] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b16 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[20] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b17 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[20] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b18 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[20] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b19 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[20] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b2 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[20] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b20 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[20] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b21 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[20] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b22 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[20] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b23 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[20] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b24 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[20] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b25 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[20] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b26 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[20] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b27 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[20] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b28 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[20] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b29 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[20] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b3 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[20] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b30 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[20] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b31 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[20] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b4 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[20] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b5 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[20] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b6 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[20] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b7 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[20] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b8 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[20] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg19_b9 (
    .ce(n58),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[20] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b0 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[2] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b1 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[2] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b10 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[2] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b11 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[2] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b12 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[2] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b13 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[2] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b14 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[2] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b15 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[2] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b16 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[2] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b17 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[2] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b18 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[2] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b19 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[2] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b2 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[2] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b20 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[2] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b21 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[2] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b22 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[2] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b23 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[2] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b24 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[2] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b25 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[2] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b26 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[2] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b27 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[2] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b28 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[2] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b29 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[2] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b3 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[2] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b30 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[2] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b31 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[2] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b4 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[2] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b5 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[2] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b6 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[2] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b7 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[2] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b8 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[2] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b9 (
    .ce(n4),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[2] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b0 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[21] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b1 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[21] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b10 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[21] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b11 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[21] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b12 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[21] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b13 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[21] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b14 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[21] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b15 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[21] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b16 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[21] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b17 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[21] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b18 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[21] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b19 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[21] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b2 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[21] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b20 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[21] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b21 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[21] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b22 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[21] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b23 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[21] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b24 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[21] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b25 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[21] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b26 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[21] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b27 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[21] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b28 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[21] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b29 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[21] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b3 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[21] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b30 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[21] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b31 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[21] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b4 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[21] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b5 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[21] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b6 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[21] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b7 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[21] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b8 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[21] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg20_b9 (
    .ce(n61),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[21] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b0 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[22] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b1 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[22] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b10 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[22] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b11 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[22] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b12 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[22] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b13 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[22] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b14 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[22] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b15 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[22] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b16 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[22] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b17 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[22] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b18 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[22] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b19 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[22] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b2 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[22] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b20 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[22] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b21 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[22] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b22 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[22] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b23 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[22] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b24 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[22] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b25 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[22] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b26 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[22] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b27 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[22] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b28 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[22] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b29 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[22] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b3 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[22] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b30 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[22] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b31 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[22] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b4 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[22] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b5 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[22] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b6 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[22] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b7 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[22] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b8 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[22] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg21_b9 (
    .ce(n64),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[22] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b0 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[23] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b1 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[23] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b10 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[23] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b11 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[23] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b12 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[23] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b13 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[23] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b14 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[23] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b15 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[23] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b16 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[23] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b17 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[23] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b18 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[23] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b19 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[23] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b2 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[23] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b20 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[23] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b21 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[23] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b22 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[23] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b23 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[23] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b24 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[23] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b25 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[23] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b26 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[23] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b27 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[23] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b28 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[23] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b29 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[23] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b3 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[23] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b30 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[23] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b31 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[23] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b4 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[23] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b5 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[23] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b6 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[23] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b7 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[23] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b8 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[23] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg22_b9 (
    .ce(n67),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[23] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b0 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[24] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b1 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[24] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b10 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[24] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b11 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[24] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b12 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[24] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b13 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[24] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b14 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[24] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b15 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[24] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b16 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[24] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b17 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[24] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b18 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[24] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b19 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[24] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b2 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[24] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b20 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[24] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b21 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[24] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b22 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[24] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b23 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[24] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b24 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[24] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b25 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[24] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b26 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[24] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b27 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[24] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b28 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[24] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b29 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[24] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b3 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[24] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b30 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[24] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b31 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[24] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b4 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[24] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b5 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[24] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b6 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[24] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b7 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[24] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b8 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[24] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg23_b9 (
    .ce(n70),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[24] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b0 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[25] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b1 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[25] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b10 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[25] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b11 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[25] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b12 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[25] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b13 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[25] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b14 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[25] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b15 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[25] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b16 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[25] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b17 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[25] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b18 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[25] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b19 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[25] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b2 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[25] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b20 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[25] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b21 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[25] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b22 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[25] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b23 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[25] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b24 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[25] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b25 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[25] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b26 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[25] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b27 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[25] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b28 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[25] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b29 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[25] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b3 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[25] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b30 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[25] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b31 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[25] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b4 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[25] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b5 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[25] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b6 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[25] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b7 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[25] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b8 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[25] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg24_b9 (
    .ce(n73),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[25] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b0 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[26] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b1 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[26] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b10 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[26] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b11 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[26] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b12 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[26] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b13 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[26] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b14 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[26] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b15 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[26] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b16 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[26] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b17 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[26] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b18 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[26] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b19 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[26] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b2 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[26] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b20 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[26] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b21 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[26] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b22 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[26] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b23 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[26] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b24 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[26] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b25 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[26] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b26 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[26] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b27 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[26] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b28 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[26] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b29 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[26] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b3 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[26] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b30 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[26] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b31 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[26] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b4 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[26] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b5 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[26] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b6 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[26] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b7 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[26] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b8 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[26] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg25_b9 (
    .ce(n76),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[26] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b0 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[27] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b1 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[27] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b10 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[27] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b11 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[27] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b12 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[27] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b13 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[27] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b14 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[27] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b15 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[27] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b16 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[27] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b17 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[27] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b18 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[27] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b19 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[27] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b2 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[27] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b20 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[27] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b21 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[27] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b22 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[27] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b23 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[27] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b24 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[27] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b25 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[27] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b26 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[27] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b27 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[27] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b28 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[27] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b29 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[27] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b3 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[27] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b30 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[27] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b31 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[27] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b4 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[27] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b5 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[27] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b6 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[27] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b7 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[27] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b8 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[27] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg26_b9 (
    .ce(n79),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[27] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b0 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[28] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b1 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[28] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b10 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[28] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b11 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[28] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b12 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[28] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b13 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[28] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b14 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[28] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b15 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[28] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b16 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[28] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b17 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[28] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b18 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[28] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b19 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[28] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b2 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[28] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b20 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[28] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b21 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[28] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b22 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[28] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b23 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[28] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b24 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[28] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b25 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[28] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b26 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[28] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b27 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[28] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b28 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[28] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b29 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[28] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b3 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[28] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b30 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[28] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b31 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[28] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b4 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[28] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b5 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[28] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b6 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[28] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b7 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[28] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b8 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[28] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg27_b9 (
    .ce(n82),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[28] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b0 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[29] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b1 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[29] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b10 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[29] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b11 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[29] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b12 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[29] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b13 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[29] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b14 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[29] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b15 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[29] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b16 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[29] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b17 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[29] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b18 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[29] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b19 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[29] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b2 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[29] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b20 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[29] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b21 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[29] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b22 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[29] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b23 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[29] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b24 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[29] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b25 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[29] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b26 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[29] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b27 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[29] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b28 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[29] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b29 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[29] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b3 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[29] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b30 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[29] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b31 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[29] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b4 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[29] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b5 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[29] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b6 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[29] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b7 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[29] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b8 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[29] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg28_b9 (
    .ce(n85),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[29] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b0 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[30] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b1 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[30] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b10 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[30] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b11 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[30] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b12 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[30] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b13 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[30] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b14 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[30] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b15 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[30] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b16 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[30] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b17 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[30] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b18 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[30] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b19 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[30] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b2 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[30] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b20 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[30] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b21 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[30] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b22 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[30] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b23 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[30] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b24 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[30] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b25 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[30] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b26 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[30] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b27 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[30] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b28 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[30] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b29 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[30] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b3 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[30] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b30 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[30] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b31 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[30] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b4 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[30] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b5 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[30] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b6 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[30] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b7 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[30] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b8 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[30] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg29_b9 (
    .ce(n88),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[30] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b0 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[3] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b1 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[3] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b10 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[3] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b11 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[3] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b12 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[3] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b13 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[3] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b14 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[3] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b15 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[3] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b16 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[3] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b17 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[3] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b18 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[3] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b19 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[3] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b2 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[3] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b20 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[3] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b21 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[3] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b22 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[3] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b23 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[3] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b24 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[3] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b25 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[3] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b26 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[3] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b27 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[3] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b28 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[3] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b29 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[3] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b3 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[3] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b30 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[3] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b31 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[3] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b4 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[3] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b5 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[3] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b6 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[3] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b7 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[3] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b8 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[3] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg2_b9 (
    .ce(n7),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[3] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b0 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[31] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b1 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[31] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b10 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[31] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b11 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[31] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b12 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[31] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b13 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[31] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b14 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[31] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b15 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[31] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b16 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[31] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b17 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[31] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b18 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[31] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b19 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[31] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b2 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[31] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b20 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[31] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b21 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[31] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b22 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[31] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b23 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[31] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b24 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[31] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b25 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[31] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b26 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[31] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b27 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[31] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b28 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[31] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b29 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[31] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b3 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[31] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b30 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[31] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b31 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[31] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b4 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[31] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b5 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[31] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b6 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[31] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b7 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[31] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b8 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[31] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg30_b9 (
    .ce(n91),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[31] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b0 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[4] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b1 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[4] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b10 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[4] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b11 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[4] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b12 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[4] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b13 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[4] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b14 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[4] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b15 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[4] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b16 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[4] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b17 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[4] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b18 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[4] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b19 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[4] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b2 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[4] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b20 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[4] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b21 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[4] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b22 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[4] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b23 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[4] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b24 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[4] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b25 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[4] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b26 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[4] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b27 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[4] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b28 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[4] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b29 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[4] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b3 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[4] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b30 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[4] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b31 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[4] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b4 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[4] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b5 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[4] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b6 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[4] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b7 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[4] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b8 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[4] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg3_b9 (
    .ce(n10),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[4] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b0 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[5] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b1 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[5] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b10 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[5] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b11 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[5] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b12 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[5] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b13 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[5] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b14 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[5] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b15 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[5] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b16 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[5] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b17 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[5] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b18 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[5] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b19 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[5] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b2 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[5] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b20 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[5] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b21 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[5] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b22 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[5] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b23 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[5] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b24 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[5] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b25 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[5] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b26 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[5] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b27 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[5] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b28 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[5] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b29 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[5] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b3 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[5] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b30 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[5] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b31 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[5] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b4 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[5] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b5 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[5] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b6 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[5] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b7 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[5] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b8 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[5] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg4_b9 (
    .ce(n13),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[5] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b0 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[6] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b1 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[6] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b10 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[6] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b11 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[6] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b12 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[6] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b13 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[6] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b14 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[6] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b15 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[6] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b16 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[6] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b17 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[6] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b18 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[6] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b19 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[6] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b2 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[6] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b20 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[6] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b21 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[6] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b22 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[6] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b23 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[6] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b24 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[6] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b25 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[6] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b26 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[6] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b27 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[6] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b28 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[6] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b29 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[6] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b3 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[6] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b30 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[6] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b31 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[6] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b4 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[6] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b5 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[6] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b6 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[6] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b7 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[6] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b8 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[6] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg5_b9 (
    .ce(n16),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[6] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b0 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[7] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b1 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[7] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b10 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[7] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b11 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[7] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b12 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[7] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b13 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[7] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b14 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[7] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b15 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[7] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b16 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[7] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b17 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[7] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b18 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[7] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b19 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[7] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b2 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[7] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b20 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[7] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b21 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[7] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b22 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[7] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b23 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[7] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b24 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[7] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b25 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[7] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b26 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[7] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b27 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[7] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b28 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[7] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b29 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[7] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b3 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[7] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b30 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[7] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b31 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[7] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b4 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[7] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b5 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[7] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b6 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[7] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b7 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[7] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b8 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[7] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg6_b9 (
    .ce(n19),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[7] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b0 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[8] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b1 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[8] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b10 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[8] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b11 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[8] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b12 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[8] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b13 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[8] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b14 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[8] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b15 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[8] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b16 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[8] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b17 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[8] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b18 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[8] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b19 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[8] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b2 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[8] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b20 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[8] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b21 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[8] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b22 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[8] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b23 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[8] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b24 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[8] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b25 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[8] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b26 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[8] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b27 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[8] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b28 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[8] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b29 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[8] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b3 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[8] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b30 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[8] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b31 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[8] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b4 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[8] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b5 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[8] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b6 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[8] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b7 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[8] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b8 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[8] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg7_b9 (
    .ce(n22),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[8] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b0 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[9] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b1 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[9] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b10 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[9] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b11 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[9] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b12 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[9] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b13 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[9] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b14 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[9] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b15 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[9] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b16 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[9] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b17 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[9] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b18 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[9] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b19 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[9] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b2 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[9] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b20 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[9] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b21 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[9] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b22 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[9] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b23 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[9] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b24 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[9] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b25 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[9] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b26 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[9] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b27 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[9] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b28 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[9] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b29 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[9] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b3 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[9] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b30 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[9] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b31 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[9] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b4 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[9] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b5 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[9] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b6 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[9] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b7 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[9] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b8 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[9] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg8_b9 (
    .ce(n25),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[9] [9]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b0 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[0]),
    .q(\rfxs[10] [0]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b1 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[1]),
    .q(\rfxs[10] [1]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b10 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[10]),
    .q(\rfxs[10] [10]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b11 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[11]),
    .q(\rfxs[10] [11]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b12 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[12]),
    .q(\rfxs[10] [12]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b13 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[13]),
    .q(\rfxs[10] [13]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b14 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[14]),
    .q(\rfxs[10] [14]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b15 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[15]),
    .q(\rfxs[10] [15]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b16 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[16]),
    .q(\rfxs[10] [16]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b17 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[17]),
    .q(\rfxs[10] [17]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b18 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[18]),
    .q(\rfxs[10] [18]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b19 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[19]),
    .q(\rfxs[10] [19]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b2 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[2]),
    .q(\rfxs[10] [2]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b20 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[20]),
    .q(\rfxs[10] [20]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b21 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[21]),
    .q(\rfxs[10] [21]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b22 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[22]),
    .q(\rfxs[10] [22]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b23 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[23]),
    .q(\rfxs[10] [23]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b24 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[24]),
    .q(\rfxs[10] [24]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b25 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[25]),
    .q(\rfxs[10] [25]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b26 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[26]),
    .q(\rfxs[10] [26]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b27 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[27]),
    .q(\rfxs[10] [27]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b28 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[28]),
    .q(\rfxs[10] [28]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b29 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[29]),
    .q(\rfxs[10] [29]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b3 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[3]),
    .q(\rfxs[10] [3]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b30 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[30]),
    .q(\rfxs[10] [30]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b31 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[31]),
    .q(\rfxs[10] [31]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b4 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[4]),
    .q(\rfxs[10] [4]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b5 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[5]),
    .q(\rfxs[10] [5]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b6 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[6]),
    .q(\rfxs[10] [6]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b7 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[7]),
    .q(\rfxs[10] [7]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b8 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[8]),
    .q(\rfxs[10] [8]));  // ../RTL/core/regfile.v(36)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg9_b9 (
    .ce(n28),
    .clk(i_clk),
    .d(i_rd_wdata[9]),
    .q(\rfxs[10] [9]));  // ../RTL/core/regfile.v(36)

endmodule 

module FPU32  // ../RTL/core/fpu.v(7)
  (
  i_clk,
  i_op1,
  i_op2,
  i_rsn,
  o_addres,
  o_divres,
  o_mulres,
  o_subres
  );

  input i_clk;  // ../RTL/core/fpu.v(8)
  input [31:0] i_op1;  // ../RTL/core/fpu.v(11)
  input [31:0] i_op2;  // ../RTL/core/fpu.v(12)
  input i_rsn;  // ../RTL/core/fpu.v(9)
  output [31:0] o_addres;  // ../RTL/core/fpu.v(15)
  output [31:0] o_divres;  // ../RTL/core/fpu.v(18)
  output [31:0] o_mulres;  // ../RTL/core/fpu.v(17)
  output [31:0] o_subres;  // ../RTL/core/fpu.v(16)

  wire [24:0] n0;
  wire [29:0] n1;
  wire [23:0] \u_mul/normalized_M_mul_result ;  // ../RTL/core/fpu.v(254)
  wire [8:0] \u_mul/sum_E ;  // ../RTL/core/fpu.v(252)
  wire _al_u11_o;
  wire _al_u15_o;
  wire _al_u18_o;
  wire _al_u19_o;
  wire _al_u1_o;
  wire _al_u20_o;
  wire _al_u21_o;
  wire _al_u22_o;
  wire _al_u23_o;
  wire _al_u24_o;
  wire _al_u26_o;
  wire _al_u29_o;
  wire _al_u30_o;
  wire _al_u33_o;
  wire _al_u37_o;
  wire _al_u3_o;
  wire _al_u40_o;
  wire _al_u43_o;
  wire _al_u46_o;
  wire _al_u51_o;
  wire _al_u57_o;
  wire _al_u59_o;
  wire _al_u5_o;
  wire _al_u60_o;
  wire _al_u63_o;
  wire _al_u66_o;
  wire _al_u68_o;
  wire _al_u6_o;
  wire _al_u71_o;
  wire _al_u73_o;
  wire _al_u75_o;
  wire _al_u77_o;
  wire _al_u82_o;
  wire _al_u85_o;
  wire _al_u87_o;
  wire _al_u88_o;
  wire _al_u8_o;
  wire _al_u92_o;
  wire _al_u9_o;
  wire \u1/c1 ;
  wire \u1/c11 ;
  wire \u1/c13 ;
  wire \u1/c15 ;
  wire \u1/c17 ;
  wire \u1/c19 ;
  wire \u1/c21 ;
  wire \u1/c23 ;
  wire \u1/c3 ;
  wire \u1/c5 ;
  wire \u1/c7 ;
  wire \u1/c9 ;
  wire \u2/c11 ;
  wire \u2/c15 ;
  wire \u2/c19 ;
  wire \u2/c23 ;
  wire \u2/c27 ;
  wire \u2/c3 ;
  wire \u2/c7 ;
  wire \u_mul/ADD02/ADD01/ADD01/n17 ;
  wire \u_mul/ADD02/ADD01/ADD02/n11 ;
  wire \u_mul/ADD02/ADD01/ADD02/n7 ;
  wire \u_mul/ADD23/ADD01/ADD01/n17 ;
  wire \u_mul/ADD23/ADD01/ADD01/p0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \u_mul/ADD23/ADD01/ADD02/n10 ;
  wire \u_mul/ADD23/ADD01/ADD02/n21 ;
  wire \u_mul/ADD23/ADD01/ADD02/n3 ;
  wire \u_mul/ADD23/ADD02/ADD01/n20 ;
  wire \u_mul/ADD23/ADD02/ADD01/n3 ;
  wire \u_mul/ADD23/ADD02/ADD02/n10 ;
  wire \u_mul/ADD23/ADD02/ADD02/n20 ;
  wire \u_mul/ADD23/ADD02/ADD02/n3 ;
  wire \u_mul/ADD23/ADD03/ADD01/n10 ;
  wire \u_mul/ADD23/ADD03/ADD01/n20 ;
  wire \u_mul/ADD23/ADD03/ADD01/n3 ;
  wire \u_mul/ADD23/ADD03/ADD02/n3 ;
  wire \u_mul/MUL01/mult0_0_0_0 ;
  wire \u_mul/MUL01/mult0_0_0_1 ;
  wire \u_mul/MUL01/mult0_0_0_10 ;
  wire \u_mul/MUL01/mult0_0_0_11 ;
  wire \u_mul/MUL01/mult0_0_0_12 ;
  wire \u_mul/MUL01/mult0_0_0_13 ;
  wire \u_mul/MUL01/mult0_0_0_14 ;
  wire \u_mul/MUL01/mult0_0_0_15 ;
  wire \u_mul/MUL01/mult0_0_0_16 ;
  wire \u_mul/MUL01/mult0_0_0_17 ;
  wire \u_mul/MUL01/mult0_0_0_18 ;
  wire \u_mul/MUL01/mult0_0_0_19 ;
  wire \u_mul/MUL01/mult0_0_0_2 ;
  wire \u_mul/MUL01/mult0_0_0_20 ;
  wire \u_mul/MUL01/mult0_0_0_21 ;
  wire \u_mul/MUL01/mult0_0_0_22 ;
  wire \u_mul/MUL01/mult0_0_0_23 ;
  wire \u_mul/MUL01/mult0_0_0_24 ;
  wire \u_mul/MUL01/mult0_0_0_25 ;
  wire \u_mul/MUL01/mult0_0_0_26 ;
  wire \u_mul/MUL01/mult0_0_0_27 ;
  wire \u_mul/MUL01/mult0_0_0_28 ;
  wire \u_mul/MUL01/mult0_0_0_29 ;
  wire \u_mul/MUL01/mult0_0_0_3 ;
  wire \u_mul/MUL01/mult0_0_0_30 ;
  wire \u_mul/MUL01/mult0_0_0_31 ;
  wire \u_mul/MUL01/mult0_0_0_32 ;
  wire \u_mul/MUL01/mult0_0_0_33 ;
  wire \u_mul/MUL01/mult0_0_0_34 ;
  wire \u_mul/MUL01/mult0_0_0_35 ;
  wire \u_mul/MUL01/mult0_0_0_4 ;
  wire \u_mul/MUL01/mult0_0_0_5 ;
  wire \u_mul/MUL01/mult0_0_0_6 ;
  wire \u_mul/MUL01/mult0_0_0_7 ;
  wire \u_mul/MUL01/mult0_0_0_8 ;
  wire \u_mul/MUL01/mult0_0_0_9 ;
  wire \u_mul/MUL01/mult0_0_1_0 ;
  wire \u_mul/MUL01/mult0_0_1_1 ;
  wire \u_mul/MUL01/mult0_0_1_10 ;
  wire \u_mul/MUL01/mult0_0_1_11 ;
  wire \u_mul/MUL01/mult0_0_1_12 ;
  wire \u_mul/MUL01/mult0_0_1_13 ;
  wire \u_mul/MUL01/mult0_0_1_14 ;
  wire \u_mul/MUL01/mult0_0_1_15 ;
  wire \u_mul/MUL01/mult0_0_1_16 ;
  wire \u_mul/MUL01/mult0_0_1_17 ;
  wire \u_mul/MUL01/mult0_0_1_18 ;
  wire \u_mul/MUL01/mult0_0_1_19 ;
  wire \u_mul/MUL01/mult0_0_1_2 ;
  wire \u_mul/MUL01/mult0_0_1_20 ;
  wire \u_mul/MUL01/mult0_0_1_21 ;
  wire \u_mul/MUL01/mult0_0_1_22 ;
  wire \u_mul/MUL01/mult0_0_1_23 ;
  wire \u_mul/MUL01/mult0_0_1_3 ;
  wire \u_mul/MUL01/mult0_0_1_4 ;
  wire \u_mul/MUL01/mult0_0_1_5 ;
  wire \u_mul/MUL01/mult0_0_1_6 ;
  wire \u_mul/MUL01/mult0_0_1_7 ;
  wire \u_mul/MUL01/mult0_0_1_8 ;
  wire \u_mul/MUL01/mult0_0_1_9 ;
  wire \u_mul/MUL01/mult0_1_0_0 ;
  wire \u_mul/MUL01/mult0_1_0_1 ;
  wire \u_mul/MUL01/mult0_1_0_10 ;
  wire \u_mul/MUL01/mult0_1_0_11 ;
  wire \u_mul/MUL01/mult0_1_0_12 ;
  wire \u_mul/MUL01/mult0_1_0_13 ;
  wire \u_mul/MUL01/mult0_1_0_14 ;
  wire \u_mul/MUL01/mult0_1_0_15 ;
  wire \u_mul/MUL01/mult0_1_0_16 ;
  wire \u_mul/MUL01/mult0_1_0_17 ;
  wire \u_mul/MUL01/mult0_1_0_18 ;
  wire \u_mul/MUL01/mult0_1_0_19 ;
  wire \u_mul/MUL01/mult0_1_0_2 ;
  wire \u_mul/MUL01/mult0_1_0_20 ;
  wire \u_mul/MUL01/mult0_1_0_21 ;
  wire \u_mul/MUL01/mult0_1_0_22 ;
  wire \u_mul/MUL01/mult0_1_0_23 ;
  wire \u_mul/MUL01/mult0_1_0_3 ;
  wire \u_mul/MUL01/mult0_1_0_4 ;
  wire \u_mul/MUL01/mult0_1_0_5 ;
  wire \u_mul/MUL01/mult0_1_0_6 ;
  wire \u_mul/MUL01/mult0_1_0_7 ;
  wire \u_mul/MUL01/mult0_1_0_8 ;
  wire \u_mul/MUL01/mult0_1_0_9 ;
  wire \u_mul/MUL01/mult0_1_1_0 ;
  wire \u_mul/MUL01/mult0_1_1_1 ;
  wire \u_mul/MUL01/mult0_1_1_10 ;
  wire \u_mul/MUL01/mult0_1_1_11 ;
  wire \u_mul/MUL01/mult0_1_1_2 ;
  wire \u_mul/MUL01/mult0_1_1_3 ;
  wire \u_mul/MUL01/mult0_1_1_4 ;
  wire \u_mul/MUL01/mult0_1_1_5 ;
  wire \u_mul/MUL01/mult0_1_1_6 ;
  wire \u_mul/MUL01/mult0_1_1_7 ;
  wire \u_mul/MUL01/mult0_1_1_8 ;
  wire \u_mul/MUL01/mult0_1_1_9 ;
  wire \u_mul/reduced_or_E1 ;  // ../RTL/core/fpu.v(256)

  assign o_mulres[0] = \u_mul/ADD23/ADD01/ADD01/p0 ;
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u0 (
    .a(i_op1[31]),
    .b(i_op2[31]),
    .o(o_mulres[31]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u1 (
    .a(i_op1[23]),
    .b(i_op2[23]),
    .o(_al_u1_o));
  AL_MAP_LUT5 #(
    .EQN("~(~E*~D*~C*B*A)"),
    .INIT(32'hfffffff7))
    _al_u10 (
    .a(_al_u8_o),
    .b(_al_u9_o),
    .c(i_op1[27]),
    .d(i_op1[26]),
    .e(i_op1[25]),
    .o(\u_mul/reduced_or_E1 ));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*~(B)*~(C)+A*B*~(C)+A*~(B)*C)"),
    .INIT(8'h2b))
    _al_u11 (
    .a(_al_u5_o),
    .b(i_op1[25]),
    .c(i_op2[25]),
    .o(_al_u11_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@B@A)"),
    .INIT(8'h69))
    _al_u12 (
    .a(_al_u11_o),
    .b(i_op1[26]),
    .c(i_op2[26]),
    .o(\u_mul/sum_E [3]));
  AL_MAP_LUT5 #(
    .EQN("(B@(~D*~C*~(~E*~A)))"),
    .INIT(32'hccc3ccc6))
    _al_u13 (
    .a(n1[29]),
    .b(\u_mul/sum_E [3]),
    .c(_al_u6_o),
    .d(_al_u3_o),
    .e(_al_u1_o),
    .o(o_mulres[26]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u14 (
    .a(\u_mul/sum_E [3]),
    .b(_al_u6_o),
    .c(_al_u3_o),
    .o(\u_mul/ADD02/ADD01/ADD01/n17 ));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*~(B)*~(C)+A*B*~(C)+A*~(B)*C)"),
    .INIT(8'h2b))
    _al_u15 (
    .a(_al_u11_o),
    .b(i_op1[26]),
    .c(i_op2[26]),
    .o(_al_u15_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@B@A)"),
    .INIT(8'h69))
    _al_u16 (
    .a(_al_u15_o),
    .b(i_op1[27]),
    .c(i_op2[27]),
    .o(\u_mul/sum_E [4]));
  AL_MAP_LUT4 #(
    .EQN("(C@(B*~(~D*~A)))"),
    .INIT(16'h3c78))
    _al_u17 (
    .a(n1[29]),
    .b(\u_mul/ADD02/ADD01/ADD01/n17 ),
    .c(\u_mul/sum_E [4]),
    .d(_al_u1_o),
    .o(o_mulres[27]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u18 (
    .a(n1[4]),
    .b(n1[2]),
    .c(n1[1]),
    .d(\u_mul/MUL01/mult0_0_0_15 ),
    .o(_al_u18_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u19 (
    .a(n1[3]),
    .b(n1[0]),
    .c(\u_mul/MUL01/mult0_0_0_17 ),
    .d(\u_mul/MUL01/mult0_0_0_16 ),
    .o(_al_u19_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u2 (
    .a(n1[29]),
    .b(_al_u1_o),
    .o(o_mulres[23]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u20 (
    .a(\u_mul/MUL01/mult0_0_0_14 ),
    .b(\u_mul/MUL01/mult0_0_0_13 ),
    .c(\u_mul/MUL01/mult0_0_0_12 ),
    .d(\u_mul/MUL01/mult0_0_0_11 ),
    .o(_al_u20_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u21 (
    .a(_al_u20_o),
    .b(\u_mul/MUL01/mult0_0_0_10 ),
    .c(\u_mul/MUL01/mult0_0_0_9 ),
    .d(\u_mul/MUL01/mult0_0_0_8 ),
    .e(\u_mul/MUL01/mult0_0_0_7 ),
    .o(_al_u21_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u22 (
    .a(\u_mul/MUL01/mult0_0_0_6 ),
    .b(\u_mul/MUL01/mult0_0_0_5 ),
    .c(\u_mul/MUL01/mult0_0_0_4 ),
    .d(\u_mul/MUL01/mult0_0_0_3 ),
    .o(_al_u22_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u23 (
    .a(_al_u22_o),
    .b(\u_mul/MUL01/mult0_0_0_2 ),
    .c(\u_mul/MUL01/mult0_0_0_1 ),
    .d(\u_mul/MUL01/mult0_0_0_0 ),
    .o(_al_u23_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u24 (
    .a(_al_u18_o),
    .b(_al_u19_o),
    .c(_al_u21_o),
    .d(_al_u23_o),
    .o(_al_u24_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h7827))
    _al_u25 (
    .a(n1[29]),
    .b(n1[6]),
    .c(n1[5]),
    .d(_al_u24_o),
    .o(\u_mul/ADD23/ADD01/ADD01/p0 ));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*~(B)*~(C)+A*B*~(C)+A*~(B)*C)"),
    .INIT(8'h2b))
    _al_u26 (
    .a(_al_u15_o),
    .b(i_op1[27]),
    .c(i_op2[27]),
    .o(_al_u26_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@B@A)"),
    .INIT(8'h69))
    _al_u27 (
    .a(_al_u26_o),
    .b(i_op1[28]),
    .c(i_op2[28]),
    .o(\u_mul/sum_E [5]));
  AL_MAP_LUT5 #(
    .EQN("(B@(D*C*~(~E*~A)))"),
    .INIT(32'h3ccc6ccc))
    _al_u28 (
    .a(n1[29]),
    .b(\u_mul/sum_E [5]),
    .c(\u_mul/ADD02/ADD01/ADD01/n17 ),
    .d(\u_mul/sum_E [4]),
    .e(_al_u1_o),
    .o(o_mulres[28]));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*~(B)*~(C)+A*B*~(C)+A*~(B)*C)"),
    .INIT(8'h2b))
    _al_u29 (
    .a(_al_u26_o),
    .b(i_op1[28]),
    .c(i_op2[28]),
    .o(_al_u29_o));
  AL_MAP_LUT4 #(
    .EQN("~(C@A@(D*B))"),
    .INIT(16'h69a5))
    _al_u3 (
    .a(i_op1[24]),
    .b(i_op1[23]),
    .c(i_op2[24]),
    .d(i_op2[23]),
    .o(_al_u3_o));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u30 (
    .a(_al_u29_o),
    .b(i_op1[29]),
    .c(i_op2[29]),
    .o(_al_u30_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u31 (
    .a(_al_u30_o),
    .b(\u_mul/sum_E [5]),
    .o(\u_mul/ADD02/ADD01/ADD02/n7 ));
  AL_MAP_LUT5 #(
    .EQN("(D*C*B*~(~E*~A))"),
    .INIT(32'hc0008000))
    _al_u32 (
    .a(n1[29]),
    .b(\u_mul/ADD02/ADD01/ADD02/n7 ),
    .c(\u_mul/ADD02/ADD01/ADD01/n17 ),
    .d(\u_mul/sum_E [4]),
    .e(_al_u1_o),
    .o(\u_mul/ADD02/ADD01/ADD02/n11 ));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*~(B)*~(C)+A*B*~(C)+A*~(B)*C)"),
    .INIT(8'h2b))
    _al_u33 (
    .a(_al_u29_o),
    .b(i_op1[29]),
    .c(i_op2[29]),
    .o(_al_u33_o));
  AL_MAP_LUT4 #(
    .EQN("(D@C@B@A)"),
    .INIT(16'h6996))
    _al_u34 (
    .a(\u_mul/ADD02/ADD01/ADD02/n11 ),
    .b(_al_u33_o),
    .c(i_op1[30]),
    .d(i_op2[30]),
    .o(o_mulres[30]));
  AL_MAP_LUT3 #(
    .EQN("~(A@(~C*B))"),
    .INIT(8'h59))
    _al_u35 (
    .a(_al_u30_o),
    .b(\u_mul/sum_E [5]),
    .c(o_mulres[28]),
    .o(o_mulres[29]));
  AL_MAP_LUT5 #(
    .EQN("(A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h78d82d78))
    _al_u36 (
    .a(n1[29]),
    .b(n1[7]),
    .c(n1[6]),
    .d(n1[5]),
    .e(_al_u24_o),
    .o(o_mulres[1]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h7f27))
    _al_u37 (
    .a(n1[29]),
    .b(n1[6]),
    .c(n1[5]),
    .d(_al_u24_o),
    .o(_al_u37_o));
  AL_MAP_LUT5 #(
    .EQN("(D*C*(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))"),
    .INIT(32'hd0008000))
    _al_u38 (
    .a(n1[29]),
    .b(n1[9]),
    .c(n1[8]),
    .d(n1[7]),
    .e(n1[6]),
    .o(\u_mul/ADD23/ADD01/ADD01/n17 ));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)@(B*~A))"),
    .INIT(32'hbb4bb444))
    _al_u39 (
    .a(_al_u37_o),
    .b(\u_mul/ADD23/ADD01/ADD01/n17 ),
    .c(n1[29]),
    .d(n1[10]),
    .e(n1[9]),
    .o(o_mulres[4]));
  AL_MAP_LUT3 #(
    .EQN("(B@(~C*~A))"),
    .INIT(8'hc9))
    _al_u4 (
    .a(n1[29]),
    .b(_al_u3_o),
    .c(_al_u1_o),
    .o(o_mulres[24]));
  AL_MAP_LUT5 #(
    .EQN("(B*(A*C*~(D)*~(E)+~(A)*~(C)*D*~(E)+~(A)*C*D*~(E)+A*C*D*~(E)+A*C*D*E))"),
    .INIT(32'h8000c480))
    _al_u40 (
    .a(n1[29]),
    .b(n1[7]),
    .c(n1[6]),
    .d(n1[5]),
    .e(_al_u24_o),
    .o(_al_u40_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h59e27bc0))
    _al_u41 (
    .a(_al_u40_o),
    .b(n1[29]),
    .c(n1[9]),
    .d(n1[8]),
    .e(n1[6]),
    .o(o_mulres[3]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'ha6d1b7c0))
    _al_u42 (
    .a(_al_u37_o),
    .b(n1[29]),
    .c(n1[8]),
    .d(n1[7]),
    .e(n1[6]),
    .o(o_mulres[2]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~(~B*A))"),
    .INIT(16'hd000))
    _al_u43 (
    .a(n1[29]),
    .b(n1[10]),
    .c(n1[9]),
    .d(\u_mul/ADD23/ADD01/ADD01/n17 ),
    .o(_al_u43_o));
  AL_MAP_LUT5 #(
    .EQN("((E*~(D)*~(C)+E*D*~(C)+~(E)*D*C+E*D*C)@(~B*A))"),
    .INIT(32'hdd2dd222))
    _al_u44 (
    .a(_al_u43_o),
    .b(_al_u37_o),
    .c(n1[29]),
    .d(n1[11]),
    .e(n1[10]),
    .o(o_mulres[5]));
  AL_MAP_LUT5 #(
    .EQN("(D*C*(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))"),
    .INIT(32'hd0008000))
    _al_u45 (
    .a(n1[29]),
    .b(n1[12]),
    .c(n1[11]),
    .d(n1[10]),
    .e(n1[9]),
    .o(\u_mul/ADD23/ADD01/ADD02/n10 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u46 (
    .a(n1[29]),
    .b(n1[13]),
    .c(n1[12]),
    .o(_al_u46_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u47 (
    .a(n1[29]),
    .b(n1[14]),
    .c(n1[13]),
    .o(\u_mul/normalized_M_mul_result [8]));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*C*~B*A))"),
    .INIT(32'hffdf0020))
    _al_u48 (
    .a(\u_mul/ADD23/ADD01/ADD02/n10 ),
    .b(_al_u37_o),
    .c(\u_mul/ADD23/ADD01/ADD01/n17 ),
    .d(_al_u46_o),
    .e(\u_mul/normalized_M_mul_result [8]),
    .o(o_mulres[8]));
  AL_MAP_LUT4 #(
    .EQN("~(D@(C*~B*A))"),
    .INIT(16'h20df))
    _al_u49 (
    .a(\u_mul/ADD23/ADD01/ADD02/n10 ),
    .b(_al_u37_o),
    .c(\u_mul/ADD23/ADD01/ADD01/n17 ),
    .d(_al_u46_o),
    .o(o_mulres[7]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(C)*~((D*B))+A*~(C)*~((D*B))+~(A)*C*~((D*B))+~(A)*~(C)*(D*B))"),
    .INIT(16'h175f))
    _al_u5 (
    .a(i_op1[24]),
    .b(i_op1[23]),
    .c(i_op2[24]),
    .d(i_op2[23]),
    .o(_al_u5_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hd080))
    _al_u50 (
    .a(n1[29]),
    .b(n1[11]),
    .c(n1[10]),
    .d(n1[9]),
    .o(\u_mul/ADD23/ADD01/ADD02/n3 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u51 (
    .a(n1[29]),
    .b(n1[12]),
    .c(n1[11]),
    .o(_al_u51_o));
  AL_MAP_LUT4 #(
    .EQN("~(D@(C*B*~A))"),
    .INIT(16'h40bf))
    _al_u52 (
    .a(_al_u37_o),
    .b(\u_mul/ADD23/ADD01/ADD01/n17 ),
    .c(\u_mul/ADD23/ADD01/ADD02/n3 ),
    .d(_al_u51_o),
    .o(o_mulres[6]));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u53 (
    .a(\u_mul/ADD23/ADD01/ADD02/n10 ),
    .b(_al_u37_o),
    .c(\u_mul/ADD23/ADD01/ADD01/n17 ),
    .d(_al_u46_o),
    .o(\u_mul/ADD23/ADD01/ADD02/n21 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*~(B)*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h59e27bc0))
    _al_u54 (
    .a(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .b(n1[29]),
    .c(n1[15]),
    .d(n1[14]),
    .e(n1[13]),
    .o(o_mulres[9]));
  AL_MAP_LUT4 #(
    .EQN("(C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hd080))
    _al_u55 (
    .a(n1[29]),
    .b(n1[15]),
    .c(n1[14]),
    .d(n1[13]),
    .o(\u_mul/ADD23/ADD02/ADD01/n3 ));
  AL_MAP_LUT5 #(
    .EQN("(D*A*(E*~(C)*~(B)+E*C*~(B)+~(E)*C*B+E*C*B))"),
    .INIT(32'ha2008000))
    _al_u56 (
    .a(\u_mul/ADD23/ADD02/ADD01/n3 ),
    .b(n1[29]),
    .c(n1[17]),
    .d(n1[16]),
    .e(n1[15]),
    .o(\u_mul/ADD23/ADD02/ADD01/n20 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u57 (
    .a(n1[29]),
    .b(n1[18]),
    .c(n1[17]),
    .o(_al_u57_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@(B*A))"),
    .INIT(8'h87))
    _al_u58 (
    .a(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .b(\u_mul/ADD23/ADD02/ADD01/n20 ),
    .c(_al_u57_o),
    .o(o_mulres[12]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u59 (
    .a(n1[29]),
    .b(n1[17]),
    .c(n1[16]),
    .o(_al_u59_o));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u6 (
    .a(_al_u5_o),
    .b(i_op1[25]),
    .c(i_op2[25]),
    .o(_al_u6_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u60 (
    .a(n1[29]),
    .b(n1[16]),
    .c(n1[15]),
    .o(_al_u60_o));
  AL_MAP_LUT4 #(
    .EQN("~(C@(~D*B*A))"),
    .INIT(16'h0f87))
    _al_u61 (
    .a(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .b(\u_mul/ADD23/ADD02/ADD01/n3 ),
    .c(_al_u59_o),
    .d(_al_u60_o),
    .o(o_mulres[11]));
  AL_MAP_LUT3 #(
    .EQN("~(C@(B*A))"),
    .INIT(8'h87))
    _al_u62 (
    .a(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .b(\u_mul/ADD23/ADD02/ADD01/n3 ),
    .c(_al_u60_o),
    .o(o_mulres[10]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u63 (
    .a(n1[29]),
    .b(n1[19]),
    .c(n1[18]),
    .o(_al_u63_o));
  AL_MAP_LUT4 #(
    .EQN("~(C@(~D*B*A))"),
    .INIT(16'h0f87))
    _al_u64 (
    .a(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .b(\u_mul/ADD23/ADD02/ADD01/n20 ),
    .c(_al_u63_o),
    .d(_al_u57_o),
    .o(o_mulres[13]));
  AL_MAP_LUT4 #(
    .EQN("(C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hd080))
    _al_u65 (
    .a(n1[29]),
    .b(n1[19]),
    .c(n1[18]),
    .d(n1[17]),
    .o(\u_mul/ADD23/ADD02/ADD02/n3 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u66 (
    .a(n1[29]),
    .b(n1[21]),
    .c(n1[19]),
    .o(_al_u66_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u67 (
    .a(\u_mul/ADD23/ADD02/ADD02/n3 ),
    .b(_al_u66_o),
    .c(n1[20]),
    .o(\u_mul/ADD23/ADD02/ADD02/n20 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u68 (
    .a(n1[29]),
    .b(n1[22]),
    .c(n1[21]),
    .o(_al_u68_o));
  AL_MAP_LUT4 #(
    .EQN("~(D@(C*B*A))"),
    .INIT(16'h807f))
    _al_u69 (
    .a(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .b(\u_mul/ADD23/ADD02/ADD02/n20 ),
    .c(\u_mul/ADD23/ADD02/ADD01/n20 ),
    .d(_al_u68_o),
    .o(o_mulres[16]));
  AL_MAP_LUT4 #(
    .EQN("~(B@(~C*~(~D*~A)))"),
    .INIT(16'h3c39))
    _al_u7 (
    .a(n1[29]),
    .b(_al_u6_o),
    .c(_al_u3_o),
    .d(_al_u1_o),
    .o(o_mulres[25]));
  AL_MAP_LUT5 #(
    .EQN("(D*C*(E*~(B)*~(A)+E*B*~(A)+~(E)*B*A+E*B*A))"),
    .INIT(32'hd0008000))
    _al_u70 (
    .a(n1[29]),
    .b(n1[20]),
    .c(n1[19]),
    .d(n1[18]),
    .e(n1[17]),
    .o(\u_mul/ADD23/ADD02/ADD02/n10 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u71 (
    .a(n1[29]),
    .b(n1[21]),
    .c(n1[20]),
    .o(_al_u71_o));
  AL_MAP_LUT4 #(
    .EQN("~(D@(C*B*A))"),
    .INIT(16'h807f))
    _al_u72 (
    .a(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .b(\u_mul/ADD23/ADD02/ADD01/n20 ),
    .c(\u_mul/ADD23/ADD02/ADD02/n10 ),
    .d(_al_u71_o),
    .o(o_mulres[15]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u73 (
    .a(n1[29]),
    .b(n1[20]),
    .c(n1[19]),
    .o(_al_u73_o));
  AL_MAP_LUT4 #(
    .EQN("~(D@(C*B*A))"),
    .INIT(16'h807f))
    _al_u74 (
    .a(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .b(\u_mul/ADD23/ADD02/ADD01/n20 ),
    .c(\u_mul/ADD23/ADD02/ADD02/n3 ),
    .d(_al_u73_o),
    .o(o_mulres[14]));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u75 (
    .a(n1[29]),
    .b(n1[23]),
    .c(n1[22]),
    .o(_al_u75_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@(~E*C*B*A))"),
    .INIT(32'h00ff807f))
    _al_u76 (
    .a(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .b(\u_mul/ADD23/ADD02/ADD02/n20 ),
    .c(\u_mul/ADD23/ADD02/ADD01/n20 ),
    .d(_al_u75_o),
    .e(_al_u68_o),
    .o(o_mulres[17]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u77 (
    .a(n1[23]),
    .b(n1[22]),
    .o(_al_u77_o));
  AL_MAP_LUT5 #(
    .EQN("(D*A*(E*~(C)*~(B)+E*C*~(B)+~(E)*C*B+E*C*B))"),
    .INIT(32'ha2008000))
    _al_u78 (
    .a(_al_u77_o),
    .b(n1[29]),
    .c(n1[25]),
    .d(n1[24]),
    .e(n1[21]),
    .o(\u_mul/ADD23/ADD03/ADD01/n20 ));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u79 (
    .a(n1[29]),
    .b(n1[26]),
    .c(n1[25]),
    .o(\u_mul/normalized_M_mul_result [20]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u8 (
    .a(i_op1[30]),
    .b(i_op1[29]),
    .c(i_op1[28]),
    .o(_al_u8_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*C*B*A))"),
    .INIT(32'h7fff8000))
    _al_u80 (
    .a(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .b(\u_mul/ADD23/ADD02/ADD02/n20 ),
    .c(\u_mul/ADD23/ADD02/ADD01/n20 ),
    .d(\u_mul/ADD23/ADD03/ADD01/n20 ),
    .e(\u_mul/normalized_M_mul_result [20]),
    .o(o_mulres[20]));
  AL_MAP_LUT4 #(
    .EQN("(A*(D*~(C)*~(B)+D*C*~(B)+~(D)*C*B+D*C*B))"),
    .INIT(16'ha280))
    _al_u81 (
    .a(_al_u77_o),
    .b(n1[29]),
    .c(n1[24]),
    .d(n1[21]),
    .o(\u_mul/ADD23/ADD03/ADD01/n10 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u82 (
    .a(n1[29]),
    .b(n1[25]),
    .c(n1[24]),
    .o(_al_u82_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@(D*C*B*A))"),
    .INIT(32'h80007fff))
    _al_u83 (
    .a(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .b(\u_mul/ADD23/ADD02/ADD02/n20 ),
    .c(\u_mul/ADD23/ADD02/ADD01/n20 ),
    .d(\u_mul/ADD23/ADD03/ADD01/n10 ),
    .e(_al_u82_o),
    .o(o_mulres[19]));
  AL_MAP_LUT4 #(
    .EQN("(C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hd080))
    _al_u84 (
    .a(n1[29]),
    .b(n1[23]),
    .c(n1[22]),
    .d(n1[21]),
    .o(\u_mul/ADD23/ADD03/ADD01/n3 ));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u85 (
    .a(n1[29]),
    .b(n1[24]),
    .c(n1[23]),
    .o(_al_u85_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@(D*C*B*A))"),
    .INIT(32'h80007fff))
    _al_u86 (
    .a(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .b(\u_mul/ADD23/ADD02/ADD02/n20 ),
    .c(\u_mul/ADD23/ADD02/ADD01/n20 ),
    .d(\u_mul/ADD23/ADD03/ADD01/n3 ),
    .e(_al_u85_o),
    .o(o_mulres[18]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u87 (
    .a(n1[24]),
    .b(n1[23]),
    .c(n1[22]),
    .o(_al_u87_o));
  AL_MAP_LUT5 #(
    .EQN("(D*A*(E*~(C)*~(B)+E*C*~(B)+~(E)*C*B+E*C*B))"),
    .INIT(32'ha2008000))
    _al_u88 (
    .a(_al_u87_o),
    .b(n1[29]),
    .c(n1[26]),
    .d(n1[25]),
    .e(n1[21]),
    .o(_al_u88_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u89 (
    .a(n1[29]),
    .b(n1[27]),
    .c(n1[26]),
    .o(\u_mul/normalized_M_mul_result [21]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u9 (
    .a(i_op1[24]),
    .b(i_op1[23]),
    .o(_al_u9_o));
  AL_MAP_LUT4 #(
    .EQN("(C@(~D*B*A))"),
    .INIT(16'hf078))
    _al_u90 (
    .a(\u_mul/ADD23/ADD02/ADD02/n20 ),
    .b(_al_u88_o),
    .c(\u_mul/normalized_M_mul_result [21]),
    .d(o_mulres[12]),
    .o(o_mulres[21]));
  AL_MAP_LUT4 #(
    .EQN("(C*(D*~(B)*~(A)+D*B*~(A)+~(D)*B*A+D*B*A))"),
    .INIT(16'hd080))
    _al_u91 (
    .a(n1[29]),
    .b(n1[27]),
    .c(n1[26]),
    .d(n1[25]),
    .o(\u_mul/ADD23/ADD03/ADD02/n3 ));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*A)"),
    .INIT(32'h00800000))
    _al_u92 (
    .a(\u_mul/ADD23/ADD03/ADD01/n20 ),
    .b(\u_mul/ADD23/ADD03/ADD02/n3 ),
    .c(\u_mul/ADD23/ADD02/ADD02/n3 ),
    .d(_al_u66_o),
    .e(n1[20]),
    .o(_al_u92_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'hd8))
    _al_u93 (
    .a(n1[29]),
    .b(n1[28]),
    .c(n1[27]),
    .o(\u_mul/normalized_M_mul_result [22]));
  AL_MAP_LUT4 #(
    .EQN("(C@(D*B*A))"),
    .INIT(16'h78f0))
    _al_u94 (
    .a(_al_u92_o),
    .b(\u_mul/ADD23/ADD02/ADD01/n20 ),
    .c(\u_mul/normalized_M_mul_result [22]),
    .d(\u_mul/ADD23/ADD01/ADD02/n21 ),
    .o(o_mulres[22]));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u0|u1/ucin  (
    .a({\u_mul/MUL01/mult0_0_1_0 ,1'b0}),
    .b({\u_mul/MUL01/mult0_0_0_18 ,open_n0}),
    .f({n0[0],open_n20}),
    .fco(\u1/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u10|u1/u9  (
    .a({\u_mul/MUL01/mult0_0_1_10 ,\u_mul/MUL01/mult0_0_1_9 }),
    .b({\u_mul/MUL01/mult0_0_0_28 ,\u_mul/MUL01/mult0_0_0_27 }),
    .fci(\u1/c9 ),
    .f(n0[10:9]),
    .fco(\u1/c11 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u12|u1/u11  (
    .a({\u_mul/MUL01/mult0_0_1_12 ,\u_mul/MUL01/mult0_0_1_11 }),
    .b({\u_mul/MUL01/mult0_0_0_30 ,\u_mul/MUL01/mult0_0_0_29 }),
    .fci(\u1/c11 ),
    .f(n0[12:11]),
    .fco(\u1/c13 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u14|u1/u13  (
    .a({\u_mul/MUL01/mult0_0_1_14 ,\u_mul/MUL01/mult0_0_1_13 }),
    .b({\u_mul/MUL01/mult0_0_0_32 ,\u_mul/MUL01/mult0_0_0_31 }),
    .fci(\u1/c13 ),
    .f(n0[14:13]),
    .fco(\u1/c15 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u16|u1/u15  (
    .a({\u_mul/MUL01/mult0_0_1_16 ,\u_mul/MUL01/mult0_0_1_15 }),
    .b({\u_mul/MUL01/mult0_0_0_34 ,\u_mul/MUL01/mult0_0_0_33 }),
    .fci(\u1/c15 ),
    .f(n0[16:15]),
    .fco(\u1/c17 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u18|u1/u17  (
    .a({\u_mul/MUL01/mult0_0_1_18 ,\u_mul/MUL01/mult0_0_1_17 }),
    .b({\u_mul/MUL01/mult0_1_1_0 ,\u_mul/MUL01/mult0_0_0_35 }),
    .fci(\u1/c17 ),
    .f(n0[18:17]),
    .fco(\u1/c19 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u20|u1/u19  (
    .a({\u_mul/MUL01/mult0_0_1_20 ,\u_mul/MUL01/mult0_0_1_19 }),
    .b({\u_mul/MUL01/mult0_1_1_2 ,\u_mul/MUL01/mult0_1_1_1 }),
    .fci(\u1/c19 ),
    .f(n0[20:19]),
    .fco(\u1/c21 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u22|u1/u21  (
    .a({\u_mul/MUL01/mult0_0_1_22 ,\u_mul/MUL01/mult0_0_1_21 }),
    .b({\u_mul/MUL01/mult0_1_1_4 ,\u_mul/MUL01/mult0_1_1_3 }),
    .fci(\u1/c21 ),
    .f(n0[22:21]),
    .fco(\u1/c23 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u2|u1/u1  (
    .a({\u_mul/MUL01/mult0_0_1_2 ,\u_mul/MUL01/mult0_0_1_1 }),
    .b({\u_mul/MUL01/mult0_0_0_20 ,\u_mul/MUL01/mult0_0_0_19 }),
    .fci(\u1/c1 ),
    .f(n0[2:1]),
    .fco(\u1/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u4|u1/u3  (
    .a({\u_mul/MUL01/mult0_0_1_4 ,\u_mul/MUL01/mult0_0_1_3 }),
    .b({\u_mul/MUL01/mult0_0_0_22 ,\u_mul/MUL01/mult0_0_0_21 }),
    .fci(\u1/c3 ),
    .f(n0[4:3]),
    .fco(\u1/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u6|u1/u5  (
    .a({\u_mul/MUL01/mult0_0_1_6 ,\u_mul/MUL01/mult0_0_1_5 }),
    .b({\u_mul/MUL01/mult0_0_0_24 ,\u_mul/MUL01/mult0_0_0_23 }),
    .fci(\u1/c5 ),
    .f(n0[6:5]),
    .fco(\u1/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/u8|u1/u7  (
    .a({\u_mul/MUL01/mult0_0_1_8 ,\u_mul/MUL01/mult0_0_1_7 }),
    .b({\u_mul/MUL01/mult0_0_0_26 ,\u_mul/MUL01/mult0_0_0_25 }),
    .fci(\u1/c7 ),
    .f(n0[8:7]),
    .fco(\u1/c9 ));
  EG_PHY_MSLICE #(
    //.MACRO("u1/u0|u1/ucin"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u1/ucout|u1/u23  (
    .a({open_n267,\u_mul/MUL01/mult0_0_1_23 }),
    .b({open_n268,\u_mul/MUL01/mult0_1_1_5 }),
    .fci(\u1/c23 ),
    .f(n0[24:23]));
  EG_PHY_LSLICE #(
    //.MACRO("u2/ucin_al_u95"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2/u11_al_u98  (
    .a({\u_mul/MUL01/mult0_1_0_13 ,\u_mul/MUL01/mult0_1_0_11 }),
    .b({\u_mul/MUL01/mult0_1_0_14 ,\u_mul/MUL01/mult0_1_0_12 }),
    .c(2'b00),
    .d({n0[13],n0[11]}),
    .e({n0[14],n0[12]}),
    .fci(\u2/c11 ),
    .f({n1[13],n1[11]}),
    .fco(\u2/c15 ),
    .fx({n1[14],n1[12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2/ucin_al_u95"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2/u15_al_u99  (
    .a({\u_mul/MUL01/mult0_1_0_17 ,\u_mul/MUL01/mult0_1_0_15 }),
    .b({\u_mul/MUL01/mult0_1_0_18 ,\u_mul/MUL01/mult0_1_0_16 }),
    .c(2'b00),
    .d({n0[17],n0[15]}),
    .e({n0[18],n0[16]}),
    .fci(\u2/c15 ),
    .f({n1[17],n1[15]}),
    .fco(\u2/c19 ),
    .fx({n1[18],n1[16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2/ucin_al_u95"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2/u19_al_u100  (
    .a({\u_mul/MUL01/mult0_1_0_21 ,\u_mul/MUL01/mult0_1_0_19 }),
    .b({\u_mul/MUL01/mult0_1_0_22 ,\u_mul/MUL01/mult0_1_0_20 }),
    .c(2'b00),
    .d({n0[21],n0[19]}),
    .e({n0[22],n0[20]}),
    .fci(\u2/c19 ),
    .f({n1[21],n1[19]}),
    .fco(\u2/c23 ),
    .fx({n1[22],n1[20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2/ucin_al_u95"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2/u23_al_u101  (
    .a({1'b0,\u_mul/MUL01/mult0_1_0_23 }),
    .b({1'b0,\u_mul/MUL01/mult0_1_1_6 }),
    .c(2'b00),
    .d({\u_mul/MUL01/mult0_1_1_7 ,n0[23]}),
    .e({\u_mul/MUL01/mult0_1_1_8 ,n0[24]}),
    .fci(\u2/c23 ),
    .f({n1[25],n1[23]}),
    .fco(\u2/c27 ),
    .fx({n1[26],n1[24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2/ucin_al_u95"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2/u27_al_u102  (
    .a(2'b00),
    .b({open_n364,1'b0}),
    .c(2'b00),
    .d({\u_mul/MUL01/mult0_1_1_11 ,\u_mul/MUL01/mult0_1_1_9 }),
    .e({open_n367,\u_mul/MUL01/mult0_1_1_10 }),
    .fci(\u2/c27 ),
    .f({n1[29],n1[27]}),
    .fx({open_n383,n1[28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2/ucin_al_u95"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2/u3_al_u96  (
    .a({\u_mul/MUL01/mult0_1_0_5 ,\u_mul/MUL01/mult0_1_0_3 }),
    .b({\u_mul/MUL01/mult0_1_0_6 ,\u_mul/MUL01/mult0_1_0_4 }),
    .c(2'b00),
    .d({n0[5],n0[3]}),
    .e({n0[6],n0[4]}),
    .fci(\u2/c3 ),
    .f({n1[5],n1[3]}),
    .fco(\u2/c7 ),
    .fx({n1[6],n1[4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2/ucin_al_u95"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2/u7_al_u97  (
    .a({\u_mul/MUL01/mult0_1_0_9 ,\u_mul/MUL01/mult0_1_0_7 }),
    .b({\u_mul/MUL01/mult0_1_0_10 ,\u_mul/MUL01/mult0_1_0_8 }),
    .c(2'b00),
    .d({n0[9],n0[7]}),
    .e({n0[10],n0[8]}),
    .fci(\u2/c7 ),
    .f({n1[9],n1[7]}),
    .fco(\u2/c11 ),
    .fx({n1[10],n1[8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u2/ucin_al_u95"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u2/ucin_al_u95  (
    .a({\u_mul/MUL01/mult0_1_0_1 ,1'b0}),
    .b({\u_mul/MUL01/mult0_1_0_2 ,\u_mul/MUL01/mult0_1_0_0 }),
    .c(2'b00),
    .d({n0[1],1'b1}),
    .e({n0[2],n0[0]}),
    .f({n1[1],open_n439}),
    .fco(\u2/c3 ),
    .fx({n1[2],n1[0]}));
  add_sub_1 u_add (
    .n1(i_op1),
    .n2(i_op2),
    .sub(1'b0),
    .result(o_addres));  // ../RTL/core/fpu.v(23)
  EG_PHY_MULT18 #(
    .INPUTREGA("DISABLE"),
    .INPUTREGB("DISABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    \u_mul/MUL01/mult0_0_0_  (
    .a(i_op1[17:0]),
    .b(i_op2[17:0]),
    .p({\u_mul/MUL01/mult0_0_0_35 ,\u_mul/MUL01/mult0_0_0_34 ,\u_mul/MUL01/mult0_0_0_33 ,\u_mul/MUL01/mult0_0_0_32 ,\u_mul/MUL01/mult0_0_0_31 ,\u_mul/MUL01/mult0_0_0_30 ,\u_mul/MUL01/mult0_0_0_29 ,\u_mul/MUL01/mult0_0_0_28 ,\u_mul/MUL01/mult0_0_0_27 ,\u_mul/MUL01/mult0_0_0_26 ,\u_mul/MUL01/mult0_0_0_25 ,\u_mul/MUL01/mult0_0_0_24 ,\u_mul/MUL01/mult0_0_0_23 ,\u_mul/MUL01/mult0_0_0_22 ,\u_mul/MUL01/mult0_0_0_21 ,\u_mul/MUL01/mult0_0_0_20 ,\u_mul/MUL01/mult0_0_0_19 ,\u_mul/MUL01/mult0_0_0_18 ,\u_mul/MUL01/mult0_0_0_17 ,\u_mul/MUL01/mult0_0_0_16 ,\u_mul/MUL01/mult0_0_0_15 ,\u_mul/MUL01/mult0_0_0_14 ,\u_mul/MUL01/mult0_0_0_13 ,\u_mul/MUL01/mult0_0_0_12 ,\u_mul/MUL01/mult0_0_0_11 ,\u_mul/MUL01/mult0_0_0_10 ,\u_mul/MUL01/mult0_0_0_9 ,\u_mul/MUL01/mult0_0_0_8 ,\u_mul/MUL01/mult0_0_0_7 ,\u_mul/MUL01/mult0_0_0_6 ,\u_mul/MUL01/mult0_0_0_5 ,\u_mul/MUL01/mult0_0_0_4 ,\u_mul/MUL01/mult0_0_0_3 ,\u_mul/MUL01/mult0_0_0_2 ,\u_mul/MUL01/mult0_0_0_1 ,\u_mul/MUL01/mult0_0_0_0 }));
  EG_PHY_MULT18 #(
    .INPUTREGA("DISABLE"),
    .INPUTREGB("DISABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    \u_mul/MUL01/mult0_0_1_  (
    .a(i_op1[17:0]),
    .b({12'b000000000000,\u_mul/reduced_or_E1 ,i_op2[22:18]}),
    .p({open_n611,open_n612,open_n613,open_n614,open_n615,open_n616,open_n617,open_n618,open_n619,open_n620,open_n621,open_n622,\u_mul/MUL01/mult0_0_1_23 ,\u_mul/MUL01/mult0_0_1_22 ,\u_mul/MUL01/mult0_0_1_21 ,\u_mul/MUL01/mult0_0_1_20 ,\u_mul/MUL01/mult0_0_1_19 ,\u_mul/MUL01/mult0_0_1_18 ,\u_mul/MUL01/mult0_0_1_17 ,\u_mul/MUL01/mult0_0_1_16 ,\u_mul/MUL01/mult0_0_1_15 ,\u_mul/MUL01/mult0_0_1_14 ,\u_mul/MUL01/mult0_0_1_13 ,\u_mul/MUL01/mult0_0_1_12 ,\u_mul/MUL01/mult0_0_1_11 ,\u_mul/MUL01/mult0_0_1_10 ,\u_mul/MUL01/mult0_0_1_9 ,\u_mul/MUL01/mult0_0_1_8 ,\u_mul/MUL01/mult0_0_1_7 ,\u_mul/MUL01/mult0_0_1_6 ,\u_mul/MUL01/mult0_0_1_5 ,\u_mul/MUL01/mult0_0_1_4 ,\u_mul/MUL01/mult0_0_1_3 ,\u_mul/MUL01/mult0_0_1_2 ,\u_mul/MUL01/mult0_0_1_1 ,\u_mul/MUL01/mult0_0_1_0 }));
  EG_PHY_MULT18 #(
    .INPUTREGA("DISABLE"),
    .INPUTREGB("DISABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    \u_mul/MUL01/mult0_1_0_  (
    .a({12'b000000000000,\u_mul/reduced_or_E1 ,i_op1[22:18]}),
    .b(i_op2[17:0]),
    .p({open_n706,open_n707,open_n708,open_n709,open_n710,open_n711,open_n712,open_n713,open_n714,open_n715,open_n716,open_n717,\u_mul/MUL01/mult0_1_0_23 ,\u_mul/MUL01/mult0_1_0_22 ,\u_mul/MUL01/mult0_1_0_21 ,\u_mul/MUL01/mult0_1_0_20 ,\u_mul/MUL01/mult0_1_0_19 ,\u_mul/MUL01/mult0_1_0_18 ,\u_mul/MUL01/mult0_1_0_17 ,\u_mul/MUL01/mult0_1_0_16 ,\u_mul/MUL01/mult0_1_0_15 ,\u_mul/MUL01/mult0_1_0_14 ,\u_mul/MUL01/mult0_1_0_13 ,\u_mul/MUL01/mult0_1_0_12 ,\u_mul/MUL01/mult0_1_0_11 ,\u_mul/MUL01/mult0_1_0_10 ,\u_mul/MUL01/mult0_1_0_9 ,\u_mul/MUL01/mult0_1_0_8 ,\u_mul/MUL01/mult0_1_0_7 ,\u_mul/MUL01/mult0_1_0_6 ,\u_mul/MUL01/mult0_1_0_5 ,\u_mul/MUL01/mult0_1_0_4 ,\u_mul/MUL01/mult0_1_0_3 ,\u_mul/MUL01/mult0_1_0_2 ,\u_mul/MUL01/mult0_1_0_1 ,\u_mul/MUL01/mult0_1_0_0 }));
  EG_PHY_MULT18 #(
    .INPUTREGA("DISABLE"),
    .INPUTREGB("DISABLE"),
    .MODE("MULT9X9C"),
    .OUTPUTREG("DISABLE"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    \u_mul/MUL01/mult0_1_1_  (
    .a({open_n718,open_n719,open_n720,open_n721,open_n722,open_n723,open_n724,open_n725,open_n726,3'b000,\u_mul/reduced_or_E1 ,i_op1[22:18]}),
    .b({open_n745,open_n746,open_n747,open_n748,open_n749,open_n750,open_n751,open_n752,open_n753,3'b000,\u_mul/reduced_or_E1 ,i_op2[22:18]}),
    .p({open_n819,open_n820,open_n821,open_n822,open_n823,open_n824,open_n825,open_n826,open_n827,open_n828,open_n829,open_n830,open_n831,open_n832,open_n833,open_n834,open_n835,open_n836,open_n837,open_n838,open_n839,open_n840,open_n841,open_n842,\u_mul/MUL01/mult0_1_1_11 ,\u_mul/MUL01/mult0_1_1_10 ,\u_mul/MUL01/mult0_1_1_9 ,\u_mul/MUL01/mult0_1_1_8 ,\u_mul/MUL01/mult0_1_1_7 ,\u_mul/MUL01/mult0_1_1_6 ,\u_mul/MUL01/mult0_1_1_5 ,\u_mul/MUL01/mult0_1_1_4 ,\u_mul/MUL01/mult0_1_1_3 ,\u_mul/MUL01/mult0_1_1_2 ,\u_mul/MUL01/mult0_1_1_1 ,\u_mul/MUL01/mult0_1_1_0 }));
  add_sub u_sub (
    .n1(i_op1),
    .n2(i_op2),
    .sub(1'b1),
    .result(o_subres));  // ../RTL/core/fpu.v(33)

endmodule 

module EXU_MDU  // ../RTL/core/exu_mdu.v(14)
  (
  i_clk,
  i_decinfo_grp,
  i_flush,
  i_mdu_op1,
  i_mdu_op2,
  i_mdu_rdidx,
  i_mdu_rdwen,
  i_mduinfo,
  i_rstn,
  i_vld,
  o_mdu_rdidx,
  o_mdu_rdwdata,
  o_mdu_rdwen,
  o_will_rdidx,
  o_will_rdwen,
  o_working
  );

  input i_clk;  // ../RTL/core/exu_mdu.v(15)
  input [5:0] i_decinfo_grp;  // ../RTL/core/exu_mdu.v(21)
  input i_flush;  // ../RTL/core/exu_mdu.v(19)
  input [31:0] i_mdu_op1;  // ../RTL/core/exu_mdu.v(25)
  input [31:0] i_mdu_op2;  // ../RTL/core/exu_mdu.v(26)
  input [4:0] i_mdu_rdidx;  // ../RTL/core/exu_mdu.v(24)
  input i_mdu_rdwen;  // ../RTL/core/exu_mdu.v(23)
  input [9:0] i_mduinfo;  // ../RTL/core/exu_mdu.v(22)
  input i_rstn;  // ../RTL/core/exu_mdu.v(16)
  input i_vld;  // ../RTL/core/exu_mdu.v(18)
  output [4:0] o_mdu_rdidx;  // ../RTL/core/exu_mdu.v(36)
  output [31:0] o_mdu_rdwdata;  // ../RTL/core/exu_mdu.v(37)
  output o_mdu_rdwen;  // ../RTL/core/exu_mdu.v(35)
  output [4:0] o_will_rdidx;  // ../RTL/core/exu_mdu.v(32)
  output o_will_rdwen;  // ../RTL/core/exu_mdu.v(31)
  output o_working;  // ../RTL/core/exu_mdu.v(29)

  wire [7:0] cnt;  // ../RTL/core/exu_mdu.v(85)
  wire [31:0] div_signed_quo;  // ../RTL/core/exu_mdu.v(125)
  wire [31:0] div_signed_rem;  // ../RTL/core/exu_mdu.v(126)
  wire [31:0] div_unsigned_quo;  // ../RTL/core/exu_mdu.v(140)
  wire [31:0] div_unsigned_rem;  // ../RTL/core/exu_mdu.v(141)
  wire [9:0] mduinfo;  // ../RTL/core/exu_mdu.v(50)
  wire [45:0] n11;
  wire [45:0] n12;
  wire [45:0] n13;
  wire [7:0] n19;
  wire [45:0] n2;
  wire [7:0] n29;
  wire [31:0] n34;
  wire [31:0] n35;
  wire [31:0] n37;
  wire [31:0] n42;
  wire [31:0] n44;
  wire [45:0] n7;
  wire [32:0] n9;
  wire [5:0] \u_DIV_SIGNED/al_00000256AA0CE7C0 ;  // al_ip/div_signed_gate.v(42)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA0CEB40 ;  // al_ip/div_signed_gate.v(58)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA0CF470 ;  // al_ip/div_signed_gate.v(57)
  wire [62:0] \u_DIV_SIGNED/al_00000256AA0D0BA0 ;  // al_ip/div_signed_gate.v(43)
  wire [5:0] \u_DIV_SIGNED/al_00000256AA0D29D0 ;  // al_ip/div_signed_gate.v(48)
  wire [5:0] \u_DIV_SIGNED/al_00000256AA0D38B0 ;  // al_ip/div_signed_gate.v(53)
  wire [62:0] \u_DIV_SIGNED/al_00000256AA0D5590 ;  // al_ip/div_signed_gate.v(54)
  wire [62:0] \u_DIV_SIGNED/al_00000256AA0D7970 ;  // al_ip/div_signed_gate.v(55)
  wire [62:0] \u_DIV_SIGNED/al_00000256AA0D80E0 ;  // al_ip/div_signed_gate.v(56)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA3FF0F0 ;  // al_ip/div_signed_gate.v(44)
  wire [62:0] \u_DIV_SIGNED/al_00000256AA400D60 ;  // al_ip/div_signed_gate.v(45)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA402C70 ;  // al_ip/div_signed_gate.v(47)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA403450 ;  // al_ip/div_signed_gate.v(46)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA4072E0 ;  // al_ip/div_signed_gate.v(49)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA4073C0 ;  // al_ip/div_signed_gate.v(50)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA4098F0 ;  // al_ip/div_signed_gate.v(52)
  wire [31:0] \u_DIV_SIGNED/al_00000256AA40B170 ;  // al_ip/div_signed_gate.v(51)
  wire [5:0] \u_DIV_UNSIGNED/al_00000286E57DB3B0 ;  // al_ip/div_unsigned_gate.v(42)
  wire [31:0] \u_DIV_UNSIGNED/al_00000286E57DBF10 ;  // al_ip/div_unsigned_gate.v(50)
  wire [31:0] \u_DIV_UNSIGNED/al_00000286E57DC290 ;  // al_ip/div_unsigned_gate.v(49)
  wire [62:0] \u_DIV_UNSIGNED/al_00000286E57DE2F0 ;  // al_ip/div_unsigned_gate.v(43)
  wire [62:0] \u_DIV_UNSIGNED/al_00000286E57DEE50 ;  // al_ip/div_unsigned_gate.v(46)
  wire [5:0] \u_DIV_UNSIGNED/al_00000286E57E03C0 ;  // al_ip/div_unsigned_gate.v(44)
  wire [5:0] \u_DIV_UNSIGNED/al_00000286E57E04A0 ;  // al_ip/div_unsigned_gate.v(45)
  wire [62:0] \u_DIV_UNSIGNED/al_00000286E57E1690 ;  // al_ip/div_unsigned_gate.v(47)
  wire [31:0] \u_DIV_UNSIGNED/al_00000286E57E4870 ;  // al_ip/div_unsigned_gate.v(48)
  wire _al_u100_o;
  wire _al_u101_o;
  wire _al_u105_o;
  wire _al_u106_o;
  wire _al_u110_o;
  wire _al_u111_o;
  wire _al_u115_o;
  wire _al_u116_o;
  wire _al_u120_o;
  wire _al_u121_o;
  wire _al_u125_o;
  wire _al_u126_o;
  wire _al_u130_o;
  wire _al_u131_o;
  wire _al_u135_o;
  wire _al_u136_o;
  wire _al_u140_o;
  wire _al_u141_o;
  wire _al_u145_o;
  wire _al_u146_o;
  wire _al_u150_o;
  wire _al_u151_o;
  wire _al_u155_o;
  wire _al_u156_o;
  wire _al_u160_o;
  wire _al_u161_o;
  wire _al_u165_o;
  wire _al_u166_o;
  wire _al_u170_o;
  wire _al_u171_o;
  wire _al_u175_o;
  wire _al_u176_o;
  wire _al_u180_o;
  wire _al_u181_o;
  wire _al_u185_o;
  wire _al_u186_o;
  wire _al_u190_o;
  wire _al_u191_o;
  wire _al_u195_o;
  wire _al_u196_o;
  wire _al_u200_o;
  wire _al_u201_o;
  wire _al_u205_o;
  wire _al_u206_o;
  wire _al_u210_o;
  wire _al_u211_o;
  wire _al_u215_o;
  wire _al_u216_o;
  wire _al_u220_o;
  wire _al_u221_o;
  wire _al_u225_o;
  wire _al_u226_o;
  wire _al_u230_o;
  wire _al_u231_o;
  wire _al_u235_o;
  wire _al_u236_o;
  wire _al_u312_o;
  wire _al_u313_o;
  wire _al_u315_o;
  wire _al_u317_o;
  wire _al_u319_o;
  wire _al_u321_o;
  wire _al_u323_o;
  wire _al_u325_o;
  wire _al_u327_o;
  wire _al_u329_o;
  wire _al_u331_o;
  wire _al_u334_o;
  wire _al_u79_o;
  wire _al_u80_o;
  wire _al_u81_o;
  wire _al_u85_o;
  wire _al_u86_o;
  wire _al_u90_o;
  wire _al_u91_o;
  wire _al_u95_o;
  wire _al_u96_o;
  wire \add0/c1 ;  // ../RTL/core/exu_mdu.v(115)
  wire \add0/c3 ;  // ../RTL/core/exu_mdu.v(115)
  wire \add0/c5 ;  // ../RTL/core/exu_mdu.v(115)
  wire \add0/c7 ;  // ../RTL/core/exu_mdu.v(115)
  wire div_signed_finish;  // ../RTL/core/exu_mdu.v(124)
  wire div_signed_start;  // ../RTL/core/exu_mdu.v(127)
  wire div_unsigned_finish;  // ../RTL/core/exu_mdu.v(139)
  wire div_unsigned_start;  // ../RTL/core/exu_mdu.v(142)
  wire mdu_vld;  // ../RTL/core/exu_mdu.v(47)
  wire mul_finish;  // ../RTL/core/exu_mdu.v(89)
  wire mul_vld;  // ../RTL/core/exu_mdu.v(86)
  wire mult0_0_0_0;
  wire mult0_0_0_1;
  wire mult0_0_0_10;
  wire mult0_0_0_11;
  wire mult0_0_0_12;
  wire mult0_0_0_13;
  wire mult0_0_0_14;
  wire mult0_0_0_15;
  wire mult0_0_0_16;
  wire mult0_0_0_17;
  wire mult0_0_0_18;
  wire mult0_0_0_19;
  wire mult0_0_0_2;
  wire mult0_0_0_20;
  wire mult0_0_0_21;
  wire mult0_0_0_22;
  wire mult0_0_0_23;
  wire mult0_0_0_24;
  wire mult0_0_0_25;
  wire mult0_0_0_26;
  wire mult0_0_0_27;
  wire mult0_0_0_28;
  wire mult0_0_0_29;
  wire mult0_0_0_3;
  wire mult0_0_0_30;
  wire mult0_0_0_31;
  wire mult0_0_0_32;
  wire mult0_0_0_33;
  wire mult0_0_0_34;
  wire mult0_0_0_35;
  wire mult0_0_0_4;
  wire mult0_0_0_5;
  wire mult0_0_0_6;
  wire mult0_0_0_7;
  wire mult0_0_0_8;
  wire mult0_0_0_9;
  wire mult0_0_1_0;
  wire mult0_0_1_1;
  wire mult0_0_1_10;
  wire mult0_0_1_11;
  wire mult0_0_1_12;
  wire mult0_0_1_13;
  wire mult0_0_1_14;
  wire mult0_0_1_15;
  wire mult0_0_1_16;
  wire mult0_0_1_17;
  wire mult0_0_1_18;
  wire mult0_0_1_19;
  wire mult0_0_1_2;
  wire mult0_0_1_20;
  wire mult0_0_1_21;
  wire mult0_0_1_22;
  wire mult0_0_1_23;
  wire mult0_0_1_24;
  wire mult0_0_1_25;
  wire mult0_0_1_26;
  wire mult0_0_1_27;
  wire mult0_0_1_28;
  wire mult0_0_1_29;
  wire mult0_0_1_3;
  wire mult0_0_1_30;
  wire mult0_0_1_31;
  wire mult0_0_1_4;
  wire mult0_0_1_5;
  wire mult0_0_1_6;
  wire mult0_0_1_7;
  wire mult0_0_1_8;
  wire mult0_0_1_9;
  wire mult0_1_0_0;
  wire mult0_1_0_1;
  wire mult0_1_0_10;
  wire mult0_1_0_11;
  wire mult0_1_0_12;
  wire mult0_1_0_13;
  wire mult0_1_0_14;
  wire mult0_1_0_15;
  wire mult0_1_0_16;
  wire mult0_1_0_17;
  wire mult0_1_0_18;
  wire mult0_1_0_19;
  wire mult0_1_0_2;
  wire mult0_1_0_20;
  wire mult0_1_0_21;
  wire mult0_1_0_22;
  wire mult0_1_0_23;
  wire mult0_1_0_24;
  wire mult0_1_0_25;
  wire mult0_1_0_26;
  wire mult0_1_0_27;
  wire mult0_1_0_28;
  wire mult0_1_0_29;
  wire mult0_1_0_3;
  wire mult0_1_0_30;
  wire mult0_1_0_31;
  wire mult0_1_0_4;
  wire mult0_1_0_5;
  wire mult0_1_0_6;
  wire mult0_1_0_7;
  wire mult0_1_0_8;
  wire mult0_1_0_9;
  wire mult0_1_1_0;
  wire mult0_1_1_1;
  wire mult0_1_1_10;
  wire mult0_1_1_11;
  wire mult0_1_1_12;
  wire mult0_1_1_13;
  wire mult0_1_1_14;
  wire mult0_1_1_15;
  wire mult0_1_1_16;
  wire mult0_1_1_17;
  wire mult0_1_1_18;
  wire mult0_1_1_19;
  wire mult0_1_1_2;
  wire mult0_1_1_20;
  wire mult0_1_1_21;
  wire mult0_1_1_22;
  wire mult0_1_1_23;
  wire mult0_1_1_24;
  wire mult0_1_1_25;
  wire mult0_1_1_26;
  wire mult0_1_1_27;
  wire mult0_1_1_3;
  wire mult0_1_1_4;
  wire mult0_1_1_5;
  wire mult0_1_1_6;
  wire mult0_1_1_7;
  wire mult0_1_1_8;
  wire mult0_1_1_9;
  wire mult1_0_1_0;
  wire mult1_0_1_1;
  wire mult1_0_1_10;
  wire mult1_0_1_11;
  wire mult1_0_1_12;
  wire mult1_0_1_13;
  wire mult1_0_1_14;
  wire mult1_0_1_15;
  wire mult1_0_1_16;
  wire mult1_0_1_17;
  wire mult1_0_1_18;
  wire mult1_0_1_19;
  wire mult1_0_1_2;
  wire mult1_0_1_20;
  wire mult1_0_1_21;
  wire mult1_0_1_22;
  wire mult1_0_1_23;
  wire mult1_0_1_24;
  wire mult1_0_1_25;
  wire mult1_0_1_26;
  wire mult1_0_1_27;
  wire mult1_0_1_28;
  wire mult1_0_1_29;
  wire mult1_0_1_3;
  wire mult1_0_1_30;
  wire mult1_0_1_31;
  wire mult1_0_1_4;
  wire mult1_0_1_5;
  wire mult1_0_1_6;
  wire mult1_0_1_7;
  wire mult1_0_1_8;
  wire mult1_0_1_9;
  wire mult1_1_0_0;
  wire mult1_1_0_1;
  wire mult1_1_0_10;
  wire mult1_1_0_11;
  wire mult1_1_0_12;
  wire mult1_1_0_13;
  wire mult1_1_0_14;
  wire mult1_1_0_15;
  wire mult1_1_0_16;
  wire mult1_1_0_17;
  wire mult1_1_0_18;
  wire mult1_1_0_19;
  wire mult1_1_0_2;
  wire mult1_1_0_20;
  wire mult1_1_0_21;
  wire mult1_1_0_22;
  wire mult1_1_0_23;
  wire mult1_1_0_24;
  wire mult1_1_0_25;
  wire mult1_1_0_26;
  wire mult1_1_0_27;
  wire mult1_1_0_28;
  wire mult1_1_0_29;
  wire mult1_1_0_3;
  wire mult1_1_0_30;
  wire mult1_1_0_31;
  wire mult1_1_0_4;
  wire mult1_1_0_5;
  wire mult1_1_0_6;
  wire mult1_1_0_7;
  wire mult1_1_0_8;
  wire mult1_1_0_9;
  wire mult1_1_1_0;
  wire mult1_1_1_1;
  wire mult1_1_1_10;
  wire mult1_1_1_11;
  wire mult1_1_1_12;
  wire mult1_1_1_13;
  wire mult1_1_1_14;
  wire mult1_1_1_15;
  wire mult1_1_1_16;
  wire mult1_1_1_17;
  wire mult1_1_1_18;
  wire mult1_1_1_19;
  wire mult1_1_1_2;
  wire mult1_1_1_20;
  wire mult1_1_1_21;
  wire mult1_1_1_22;
  wire mult1_1_1_23;
  wire mult1_1_1_24;
  wire mult1_1_1_25;
  wire mult1_1_1_26;
  wire mult1_1_1_27;
  wire mult1_1_1_3;
  wire mult1_1_1_4;
  wire mult1_1_1_5;
  wire mult1_1_1_6;
  wire mult1_1_1_7;
  wire mult1_1_1_8;
  wire mult1_1_1_9;
  wire mult2_0_1_0;
  wire mult2_0_1_1;
  wire mult2_0_1_10;
  wire mult2_0_1_11;
  wire mult2_0_1_12;
  wire mult2_0_1_13;
  wire mult2_0_1_14;
  wire mult2_0_1_15;
  wire mult2_0_1_16;
  wire mult2_0_1_17;
  wire mult2_0_1_18;
  wire mult2_0_1_19;
  wire mult2_0_1_2;
  wire mult2_0_1_20;
  wire mult2_0_1_21;
  wire mult2_0_1_22;
  wire mult2_0_1_23;
  wire mult2_0_1_24;
  wire mult2_0_1_25;
  wire mult2_0_1_26;
  wire mult2_0_1_27;
  wire mult2_0_1_28;
  wire mult2_0_1_29;
  wire mult2_0_1_3;
  wire mult2_0_1_30;
  wire mult2_0_1_31;
  wire mult2_0_1_32;
  wire mult2_0_1_4;
  wire mult2_0_1_5;
  wire mult2_0_1_6;
  wire mult2_0_1_7;
  wire mult2_0_1_8;
  wire mult2_0_1_9;
  wire mult2_1_1_0;
  wire mult2_1_1_1;
  wire mult2_1_1_10;
  wire mult2_1_1_11;
  wire mult2_1_1_12;
  wire mult2_1_1_13;
  wire mult2_1_1_14;
  wire mult2_1_1_15;
  wire mult2_1_1_16;
  wire mult2_1_1_17;
  wire mult2_1_1_18;
  wire mult2_1_1_19;
  wire mult2_1_1_2;
  wire mult2_1_1_20;
  wire mult2_1_1_21;
  wire mult2_1_1_22;
  wire mult2_1_1_23;
  wire mult2_1_1_24;
  wire mult2_1_1_25;
  wire mult2_1_1_26;
  wire mult2_1_1_27;
  wire mult2_1_1_3;
  wire mult2_1_1_4;
  wire mult2_1_1_5;
  wire mult2_1_1_6;
  wire mult2_1_1_7;
  wire mult2_1_1_8;
  wire mult2_1_1_9;
  wire mux10_b0_sel_is_2_o;
  wire mux2_b0_sel_is_2_o;
  wire n10;
  wire n24_lutinv;
  wire n26;
  wire n30;
  wire n3_lutinv;
  wire n5_lutinv;
  wire n6;
  wire n8;
  wire \neg0/c11 ;  // ../RTL/core/exu_mdu.v(165)
  wire \neg0/c15 ;  // ../RTL/core/exu_mdu.v(165)
  wire \neg0/c19 ;  // ../RTL/core/exu_mdu.v(165)
  wire \neg0/c23 ;  // ../RTL/core/exu_mdu.v(165)
  wire \neg0/c27 ;  // ../RTL/core/exu_mdu.v(165)
  wire \neg0/c3 ;  // ../RTL/core/exu_mdu.v(165)
  wire \neg0/c31 ;  // ../RTL/core/exu_mdu.v(165)
  wire \neg0/c7 ;  // ../RTL/core/exu_mdu.v(165)
  wire rem_op1_sym;  // ../RTL/core/exu_mdu.v(45)
  wire \u1/c11 ;
  wire \u1/c15 ;
  wire \u1/c19 ;
  wire \u1/c23 ;
  wire \u1/c27 ;
  wire \u1/c3 ;
  wire \u1/c31 ;
  wire \u1/c35 ;
  wire \u1/c39 ;
  wire \u1/c43 ;
  wire \u1/c7 ;
  wire \u15/c11 ;
  wire \u15/c15 ;
  wire \u15/c19 ;
  wire \u15/c23 ;
  wire \u15/c27 ;
  wire \u15/c3 ;
  wire \u15/c31 ;
  wire \u15/c35 ;
  wire \u15/c39 ;
  wire \u15/c43 ;
  wire \u15/c7 ;
  wire \u5/c11 ;
  wire \u5/c15 ;
  wire \u5/c19 ;
  wire \u5/c23 ;
  wire \u5/c27 ;
  wire \u5/c3 ;
  wire \u5/c31 ;
  wire \u5/c35 ;
  wire \u5/c39 ;
  wire \u5/c43 ;
  wire \u5/c7 ;
  wire \u6/c11 ;
  wire \u6/c15 ;
  wire \u6/c19 ;
  wire \u6/c23 ;
  wire \u6/c27 ;
  wire \u6/c3 ;
  wire \u6/c31 ;
  wire \u6/c7 ;
  wire \u7/c11 ;
  wire \u7/c15 ;
  wire \u7/c19 ;
  wire \u7/c23 ;
  wire \u7/c27 ;
  wire \u7/c3 ;
  wire \u7/c31 ;
  wire \u7/c35 ;
  wire \u7/c39 ;
  wire \u7/c43 ;
  wire \u7/c7 ;
  wire \u8/c11 ;
  wire \u8/c15 ;
  wire \u8/c19 ;
  wire \u8/c23 ;
  wire \u8/c27 ;
  wire \u8/c3 ;
  wire \u8/c31 ;
  wire \u8/c35 ;
  wire \u8/c39 ;
  wire \u8/c43 ;
  wire \u8/c7 ;
  wire \u_DIV_SIGNED/al_00000256AA3DB110 ;  // al_ip/div_signed_gate.v(103)
  wire \u_DIV_SIGNED/al_00000256AA3DB320 ;  // al_ip/div_signed_gate.v(120)
  wire \u_DIV_SIGNED/al_00000256AA3DB3D0 ;  // al_ip/div_signed_gate.v(127)
  wire \u_DIV_SIGNED/al_00000256AA3DB480 ;  // al_ip/div_signed_gate.v(129)
  wire \u_DIV_SIGNED/al_00000256AA3DB5E0 ;  // al_ip/div_signed_gate.v(116)
  wire \u_DIV_SIGNED/al_00000256AA3DB7F0 ;  // al_ip/div_signed_gate.v(196)
  wire \u_DIV_SIGNED/al_00000256AA3DC030 ;  // al_ip/div_signed_gate.v(263)
  wire \u_DIV_SIGNED/al_00000256AA3DC450 ;  // al_ip/div_signed_gate.v(107)
  wire \u_DIV_SIGNED/al_00000256AA3DC5B0 ;  // al_ip/div_signed_gate.v(264)
  wire \u_DIV_SIGNED/al_00000256AA3DC870 ;  // al_ip/div_signed_gate.v(105)
  wire \u_DIV_SIGNED/al_00000256AA3DC9D0 ;  // al_ip/div_signed_gate.v(122)
  wire \u_DIV_SIGNED/al_00000256AA3DCC90 ;  // al_ip/div_signed_gate.v(114)
  wire \u_DIV_SIGNED/al_00000256AA3DD2C0 ;  // al_ip/div_signed_gate.v(101)
  wire \u_DIV_SIGNED/al_00000256AA3DD420 ;  // al_ip/div_signed_gate.v(111)
  wire \u_DIV_SIGNED/al_00000256AA3DD580 ;  // al_ip/div_signed_gate.v(118)
  wire \u_DIV_SIGNED/al_00000256AA3DD840 ;  // al_ip/div_signed_gate.v(123)
  wire \u_DIV_SIGNED/al_00000256AA3DD9A0 ;  // al_ip/div_signed_gate.v(261)
  wire \u_DIV_SIGNED/al_00000256AA3DDA50 ;  // al_ip/div_signed_gate.v(109)
  wire \u_DIV_SIGNED/al_00000256AA3DDB00 ;  // al_ip/div_signed_gate.v(125)
  wire \u_DIV_SIGNED/al_00000256AA3DEA20 ;  // al_ip/div_signed_gate.v(131)
  wire \u_DIV_SIGNED/al_00000256AA3E0300 ;  // al_ip/div_signed_gate.v(163)
  wire \u_DIV_SIGNED/al_00000256AA421080 ;  // al_ip/div_signed_gate.v(77)
  wire \u_DIV_SIGNED/al_00000256AA421130 ;  // al_ip/div_signed_gate.v(79)
  wire \u_DIV_SIGNED/al_00000256AA421550 ;  // al_ip/div_signed_gate.v(82)
  wire \u_DIV_SIGNED/al_00000256AA421600 ;  // al_ip/div_signed_gate.v(93)
  wire \u_DIV_SIGNED/al_00000256AA4216B0 ;  // al_ip/div_signed_gate.v(90)
  wire \u_DIV_SIGNED/al_00000256AA4218C0 ;  // al_ip/div_signed_gate.v(91)
  wire \u_DIV_SIGNED/al_00000256AA421C30 ;  // al_ip/div_signed_gate.v(95)
  wire \u_DIV_SIGNED/al_00000256AA421CE0 ;  // al_ip/div_signed_gate.v(88)
  wire \u_DIV_SIGNED/al_00000256AA422310 ;  // al_ip/div_signed_gate.v(86)
  wire \u_DIV_SIGNED/al_00000256AA422470 ;  // al_ip/div_signed_gate.v(97)
  wire \u_DIV_SIGNED/al_00000256AA422680 ;  // al_ip/div_signed_gate.v(262)
  wire \u_DIV_SIGNED/al_00000256AA422940 ;  // al_ip/div_signed_gate.v(75)
  wire \u_DIV_SIGNED/al_00000256AA422E10 ;  // al_ip/div_signed_gate.v(73)
  wire \u_DIV_SIGNED/al_00000256AA4232E0 ;  // al_ip/div_signed_gate.v(99)
  wire \u_DIV_SIGNED/al_00000256AA423390 ;  // al_ip/div_signed_gate.v(71)
  wire \u_DIV_SIGNED/al_00000256AA423700 ;  // al_ip/div_signed_gate.v(84)
  wire \u_DIV_SIGNED/al_00000256AA423B20 ;  // al_ip/div_signed_gate.v(69)
  wire \u_DIV_SIGNED/al_00000256AA443130 ;  // al_ip/div_signed_gate.v(150)
  wire \u_DIV_SIGNED/al_00000256AA4436B0 ;  // al_ip/div_signed_gate.v(135)
  wire \u_DIV_SIGNED/al_00000256AA443760 ;  // al_ip/div_signed_gate.v(141)
  wire \u_DIV_SIGNED/al_00000256AA443810 ;  // al_ip/div_signed_gate.v(143)
  wire \u_DIV_SIGNED/al_00000256AA443CE0 ;  // al_ip/div_signed_gate.v(137)
  wire \u_DIV_SIGNED/al_00000256AA443E40 ;  // al_ip/div_signed_gate.v(139)
  wire \u_DIV_SIGNED/al_00000256AA444100 ;  // al_ip/div_signed_gate.v(148)
  wire \u_DIV_SIGNED/al_00000256AA444260 ;  // al_ip/div_signed_gate.v(154)
  wire \u_DIV_SIGNED/al_00000256AA4445D0 ;  // al_ip/div_signed_gate.v(157)
  wire \u_DIV_SIGNED/al_00000256AA444680 ;  // al_ip/div_signed_gate.v(146)
  wire \u_DIV_SIGNED/al_00000256AA444940 ;  // al_ip/div_signed_gate.v(159)
  wire \u_DIV_SIGNED/al_00000256AA444B50 ;  // al_ip/div_signed_gate.v(152)
  wire \u_DIV_SIGNED/al_00000256AA444CB0 ;  // al_ip/div_signed_gate.v(155)
  wire \u_DIV_SIGNED/al_00000256AA444E10 ;  // al_ip/div_signed_gate.v(161)
  wire \u_DIV_SIGNED/al_00000256AA445230 ;  // al_ip/div_signed_gate.v(133)
  wire \u_DIV_SIGNED/al_00000256AA653890 ;  // al_ip/div_signed_gate.v(65)
  wire \u_DIV_SIGNED/al_00000256AA653E10 ;  // al_ip/div_signed_gate.v(67)
  wire \u_DIV_SIGNED/al_00000256AA6547B0 ;  // al_ip/div_signed_gate.v(63)
  wire \u_DIV_SIGNED/al_00000256AA88A8D0 ;  // al_ip/div_signed_gate.v(202)
  wire \u_DIV_SIGNED/al_00000256AA88A980 ;  // al_ip/div_signed_gate.v(260)
  wire \u_DIV_SIGNED/al_00000256AA88AC40 ;  // al_ip/div_signed_gate.v(187)
  wire \u_DIV_SIGNED/al_00000256AA88ADA0 ;  // al_ip/div_signed_gate.v(242)
  wire \u_DIV_SIGNED/al_00000256AA88AF00 ;  // al_ip/div_signed_gate.v(195)
  wire \u_DIV_SIGNED/al_00000256AA88B060 ;  // al_ip/div_signed_gate.v(186)
  wire \u_DIV_SIGNED/al_00000256AA88B110 ;  // al_ip/div_signed_gate.v(206)
  wire \u_DIV_SIGNED/al_00000256AA88B270 ;  // al_ip/div_signed_gate.v(191)
  wire \u_DIV_SIGNED/al_00000256AA88B480 ;  // al_ip/div_signed_gate.v(208)
  wire \u_DIV_SIGNED/al_00000256AA88B530 ;  // al_ip/div_signed_gate.v(193)
  wire \u_DIV_SIGNED/al_00000256AA88B950 ;  // al_ip/div_signed_gate.v(184)
  wire \u_DIV_SIGNED/al_00000256AA88BA00 ;  // al_ip/div_signed_gate.v(211)
  wire \u_DIV_SIGNED/al_00000256AA88BAB0 ;  // al_ip/div_signed_gate.v(213)
  wire \u_DIV_SIGNED/al_00000256AA88BC10 ;  // al_ip/div_signed_gate.v(215)
  wire \u_DIV_SIGNED/al_00000256AA88BCC0 ;  // al_ip/div_signed_gate.v(200)
  wire \u_DIV_SIGNED/al_00000256AA88BE20 ;  // al_ip/div_signed_gate.v(217)
  wire \u_DIV_SIGNED/al_00000256AA88BED0 ;  // al_ip/div_signed_gate.v(173)
  wire \u_DIV_SIGNED/al_00000256AA88C030 ;  // al_ip/div_signed_gate.v(219)
  wire \u_DIV_SIGNED/al_00000256AA88C190 ;  // al_ip/div_signed_gate.v(165)
  wire \u_DIV_SIGNED/al_00000256AA88C240 ;  // al_ip/div_signed_gate.v(169)
  wire \u_DIV_SIGNED/al_00000256AA88C3A0 ;  // al_ip/div_signed_gate.v(204)
  wire \u_DIV_SIGNED/al_00000256AA88C450 ;  // al_ip/div_signed_gate.v(220)
  wire \u_DIV_SIGNED/al_00000256AA88C500 ;  // al_ip/div_signed_gate.v(198)
  wire \u_DIV_SIGNED/al_00000256AA88C5B0 ;  // al_ip/div_signed_gate.v(180)
  wire \u_DIV_SIGNED/al_00000256AA88C660 ;  // al_ip/div_signed_gate.v(171)
  wire \u_DIV_SIGNED/al_00000256AA88C710 ;  // al_ip/div_signed_gate.v(189)
  wire \u_DIV_SIGNED/al_00000256AA88CA80 ;  // al_ip/div_signed_gate.v(182)
  wire \u_DIV_SIGNED/al_00000256AA88CBE0 ;  // al_ip/div_signed_gate.v(178)
  wire \u_DIV_SIGNED/al_00000256AA88CEA0 ;  // al_ip/div_signed_gate.v(175)
  wire \u_DIV_SIGNED/al_00000256AA88D0B0 ;  // al_ip/div_signed_gate.v(258)
  wire \u_DIV_SIGNED/al_00000256AA88D420 ;  // al_ip/div_signed_gate.v(167)
  wire \u_DIV_SIGNED/al_00000256AA88D630 ;  // al_ip/div_signed_gate.v(257)
  wire \u_DIV_SIGNED/al_00000256AA88DB00 ;  // al_ip/div_signed_gate.v(224)
  wire \u_DIV_SIGNED/al_00000256AA88DE70 ;  // al_ip/div_signed_gate.v(237)
  wire \u_DIV_SIGNED/al_00000256AA88DF20 ;  // al_ip/div_signed_gate.v(241)
  wire \u_DIV_SIGNED/al_00000256AA88DFD0 ;  // al_ip/div_signed_gate.v(248)
  wire \u_DIV_SIGNED/al_00000256AA88E130 ;  // al_ip/div_signed_gate.v(235)
  wire \u_DIV_SIGNED/al_00000256AA88E1E0 ;  // al_ip/div_signed_gate.v(239)
  wire \u_DIV_SIGNED/al_00000256AA88E340 ;  // al_ip/div_signed_gate.v(252)
  wire \u_DIV_SIGNED/al_00000256AA88EE40 ;  // al_ip/div_signed_gate.v(226)
  wire \u_DIV_SIGNED/al_00000256AA88F3C0 ;  // al_ip/div_signed_gate.v(230)
  wire \u_DIV_SIGNED/al_00000256AA88F470 ;  // al_ip/div_signed_gate.v(228)
  wire \u_DIV_SIGNED/al_00000256AA88F520 ;  // al_ip/div_signed_gate.v(244)
  wire \u_DIV_SIGNED/al_00000256AA88F680 ;  // al_ip/div_signed_gate.v(250)
  wire \u_DIV_SIGNED/al_00000256AA88F730 ;  // al_ip/div_signed_gate.v(255)
  wire \u_DIV_SIGNED/al_00000256AA88F890 ;  // al_ip/div_signed_gate.v(233)
  wire \u_DIV_SIGNED/al_00000256AA88F9F0 ;  // al_ip/div_signed_gate.v(246)
  wire \u_DIV_SIGNED/al_00000256AA88FC00 ;  // al_ip/div_signed_gate.v(222)
  wire \u_DIV_SIGNED/al_00000256AA893670 ;  // al_ip/div_signed_gate.v(59)
  wire \u_DIV_SIGNED/al_00000256AA8940C0 ;  // al_ip/div_signed_gate.v(61)
  wire \u_DIV_SIGNED/al_00000256AA895350 ;  // al_ip/div_signed_gate.v(60)
  wire \u_DIV_SIGNED/al_00000256AA898630 ;  // al_ip/div_signed_gate.v(285)
  wire \u_DIV_SIGNED/al_00000256AA898DC0 ;  // al_ip/div_signed_gate.v(276)
  wire \u_DIV_SIGNED/al_00000256AA898E70 ;  // al_ip/div_signed_gate.v(281)
  wire \u_DIV_SIGNED/al_00000256AA898FD0 ;  // al_ip/div_signed_gate.v(288)
  wire \u_DIV_SIGNED/al_00000256AA899130 ;  // al_ip/div_signed_gate.v(272)
  wire \u_DIV_SIGNED/al_00000256AA899290 ;  // al_ip/div_signed_gate.v(268)
  wire \u_DIV_SIGNED/al_00000256AA899810 ;  // al_ip/div_signed_gate.v(290)
  wire \u_DIV_SIGNED/al_00000256AA89AEC0 ;  // al_ip/div_signed_gate.v(294)
  wire \u_DIV_UNSIGNED/al_00000286E447F350 ;  // al_ip/div_unsigned_gate.v(126)
  wire \u_DIV_UNSIGNED/al_00000286E447FE50 ;  // al_ip/div_unsigned_gate.v(139)
  wire \u_DIV_UNSIGNED/al_00000286E447FF00 ;  // al_ip/div_unsigned_gate.v(143)
  wire \u_DIV_UNSIGNED/al_00000286E4480480 ;  // al_ip/div_unsigned_gate.v(136)
  wire \u_DIV_UNSIGNED/al_00000286E4480530 ;  // al_ip/div_unsigned_gate.v(145)
  wire \u_DIV_UNSIGNED/al_00000286E44805E0 ;  // al_ip/div_unsigned_gate.v(148)
  wire \u_DIV_UNSIGNED/al_00000286E44808A0 ;  // al_ip/div_unsigned_gate.v(132)
  wire \u_DIV_UNSIGNED/al_00000286E4480B60 ;  // al_ip/div_unsigned_gate.v(150)
  wire \u_DIV_UNSIGNED/al_00000286E4480CC0 ;  // al_ip/div_unsigned_gate.v(141)
  wire \u_DIV_UNSIGNED/al_00000286E44810E0 ;  // al_ip/div_unsigned_gate.v(130)
  wire \u_DIV_UNSIGNED/al_00000286E44812F0 ;  // al_ip/div_unsigned_gate.v(147)
  wire \u_DIV_UNSIGNED/al_00000286E44815B0 ;  // al_ip/div_unsigned_gate.v(152)
  wire \u_DIV_UNSIGNED/al_00000286E4481710 ;  // al_ip/div_unsigned_gate.v(154)
  wire \u_DIV_UNSIGNED/al_00000286E44819D0 ;  // al_ip/div_unsigned_gate.v(134)
  wire \u_DIV_UNSIGNED/al_00000286E4481B30 ;  // al_ip/div_unsigned_gate.v(128)
  wire \u_DIV_UNSIGNED/al_00000286E44833F0 ;  // al_ip/div_unsigned_gate.v(156)
  wire \u_DIV_UNSIGNED/al_00000286E4688A90 ;  // al_ip/div_unsigned_gate.v(51)
  wire \u_DIV_UNSIGNED/al_00000286E468A980 ;  // al_ip/div_unsigned_gate.v(52)
  wire \u_DIV_UNSIGNED/al_00000286E4A23D20 ;  // al_ip/div_unsigned_gate.v(83)
  wire \u_DIV_UNSIGNED/al_00000286E4A23F30 ;  // al_ip/div_unsigned_gate.v(65)
  wire \u_DIV_UNSIGNED/al_00000286E4A23FE0 ;  // al_ip/div_unsigned_gate.v(67)
  wire \u_DIV_UNSIGNED/al_00000286E4A24560 ;  // al_ip/div_unsigned_gate.v(54)
  wire \u_DIV_UNSIGNED/al_00000286E4A24820 ;  // al_ip/div_unsigned_gate.v(123)
  wire \u_DIV_UNSIGNED/al_00000286E4A24A30 ;  // al_ip/div_unsigned_gate.v(58)
  wire \u_DIV_UNSIGNED/al_00000286E4A24E50 ;  // al_ip/div_unsigned_gate.v(56)
  wire \u_DIV_UNSIGNED/al_00000286E4A24FB0 ;  // al_ip/div_unsigned_gate.v(121)
  wire \u_DIV_UNSIGNED/al_00000286E4A25060 ;  // al_ip/div_unsigned_gate.v(69)
  wire \u_DIV_UNSIGNED/al_00000286E4A25530 ;  // al_ip/div_unsigned_gate.v(61)
  wire \u_DIV_UNSIGNED/al_00000286E4A25690 ;  // al_ip/div_unsigned_gate.v(105)
  wire \u_DIV_UNSIGNED/al_00000286E4A25740 ;  // al_ip/div_unsigned_gate.v(63)
  wire \u_DIV_UNSIGNED/al_00000286E4A258A0 ;  // al_ip/div_unsigned_gate.v(71)
  wire \u_DIV_UNSIGNED/al_00000286E4A25950 ;  // al_ip/div_unsigned_gate.v(74)
  wire \u_DIV_UNSIGNED/al_00000286E4A25A00 ;  // al_ip/div_unsigned_gate.v(78)
  wire \u_DIV_UNSIGNED/al_00000286E4A25C10 ;  // al_ip/div_unsigned_gate.v(80)
  wire \u_DIV_UNSIGNED/al_00000286E4A25ED0 ;  // al_ip/div_unsigned_gate.v(76)
  wire \u_DIV_UNSIGNED/al_00000286E4A25F80 ;  // al_ip/div_unsigned_gate.v(82)
  wire \u_DIV_UNSIGNED/al_00000286E4A260E0 ;  // al_ip/div_unsigned_gate.v(85)
  wire \u_DIV_UNSIGNED/al_00000286E4A26A80 ;  // al_ip/div_unsigned_gate.v(91)
  wire \u_DIV_UNSIGNED/al_00000286E4A26BE0 ;  // al_ip/div_unsigned_gate.v(109)
  wire \u_DIV_UNSIGNED/al_00000286E4A26D40 ;  // al_ip/div_unsigned_gate.v(120)
  wire \u_DIV_UNSIGNED/al_00000286E4A26F50 ;  // al_ip/div_unsigned_gate.v(93)
  wire \u_DIV_UNSIGNED/al_00000286E4A270B0 ;  // al_ip/div_unsigned_gate.v(98)
  wire \u_DIV_UNSIGNED/al_00000286E4A27160 ;  // al_ip/div_unsigned_gate.v(118)
  wire \u_DIV_UNSIGNED/al_00000286E4A27210 ;  // al_ip/div_unsigned_gate.v(104)
  wire \u_DIV_UNSIGNED/al_00000286E4A272C0 ;  // al_ip/div_unsigned_gate.v(113)
  wire \u_DIV_UNSIGNED/al_00000286E4A27370 ;  // al_ip/div_unsigned_gate.v(102)
  wire \u_DIV_UNSIGNED/al_00000286E4A276E0 ;  // al_ip/div_unsigned_gate.v(96)
  wire \u_DIV_UNSIGNED/al_00000286E4A27B00 ;  // al_ip/div_unsigned_gate.v(111)
  wire \u_DIV_UNSIGNED/al_00000286E4A27BB0 ;  // al_ip/div_unsigned_gate.v(87)
  wire \u_DIV_UNSIGNED/al_00000286E4A27C60 ;  // al_ip/div_unsigned_gate.v(100)
  wire \u_DIV_UNSIGNED/al_00000286E4A28810 ;  // al_ip/div_unsigned_gate.v(89)
  wire \u_DIV_UNSIGNED/al_00000286E4A28B80 ;  // al_ip/div_unsigned_gate.v(107)
  wire \u_DIV_UNSIGNED/al_00000286E4A28E40 ;  // al_ip/div_unsigned_gate.v(115)
  wire \u_DIV_UNSIGNED/al_00000286E5A5D8C0 ;  // al_ip/div_unsigned_gate.v(59)
  wire \u_DIV_UNSIGNED/al_00000286E5A5E1B0 ;  // al_ip/div_unsigned_gate.v(124)
  wire working;  // ../RTL/core/exu_mdu.v(46)

  assign o_mdu_rdidx[4] = o_will_rdidx[4];
  assign o_mdu_rdidx[3] = o_will_rdidx[3];
  assign o_mdu_rdidx[0] = o_will_rdidx[0];
  assign o_will_rdidx[2] = o_mdu_rdidx[2];
  assign o_will_rdidx[1] = o_mdu_rdidx[1];
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u100 (
    .a(n37[4]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[4]),
    .o(_al_u100_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u101 (
    .a(_al_u100_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[4]),
    .o(_al_u101_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u102 (
    .a(_al_u101_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[4]),
    .e(div_unsigned_quo[4]),
    .o(n42[4]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u103 (
    .a(n13[18]),
    .b(n11[18]),
    .c(n42[4]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[4]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u104 (
    .a(n44[4]),
    .b(n7[18]),
    .c(mult0_0_0_4),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[4]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u105 (
    .a(n37[5]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[5]),
    .o(_al_u105_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u106 (
    .a(_al_u105_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[5]),
    .o(_al_u106_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u107 (
    .a(_al_u106_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[5]),
    .e(div_unsigned_quo[5]),
    .o(n42[5]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u108 (
    .a(n13[19]),
    .b(n11[19]),
    .c(n42[5]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[5]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u109 (
    .a(n44[5]),
    .b(n7[19]),
    .c(mult0_0_0_5),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u110 (
    .a(n37[6]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[6]),
    .o(_al_u110_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u111 (
    .a(_al_u110_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[6]),
    .o(_al_u111_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u112 (
    .a(_al_u111_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[6]),
    .e(div_unsigned_quo[6]),
    .o(n42[6]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u113 (
    .a(n13[20]),
    .b(n11[20]),
    .c(n42[6]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[6]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u114 (
    .a(n44[6]),
    .b(n7[20]),
    .c(mult0_0_0_6),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[6]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u115 (
    .a(n37[1]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[1]),
    .o(_al_u115_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u116 (
    .a(_al_u115_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[1]),
    .o(_al_u116_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u117 (
    .a(_al_u116_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[1]),
    .e(div_unsigned_quo[1]),
    .o(n42[1]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u118 (
    .a(n13[15]),
    .b(n11[15]),
    .c(n42[1]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[1]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u119 (
    .a(n44[1]),
    .b(n7[15]),
    .c(mult0_0_0_1),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[1]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u120 (
    .a(n37[11]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[11]),
    .o(_al_u120_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u121 (
    .a(_al_u120_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[11]),
    .o(_al_u121_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u122 (
    .a(_al_u121_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[11]),
    .e(div_unsigned_quo[11]),
    .o(n42[11]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u123 (
    .a(n13[25]),
    .b(n11[25]),
    .c(n42[11]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[11]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u124 (
    .a(n44[11]),
    .b(n7[25]),
    .c(mult0_0_0_11),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[11]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u125 (
    .a(n37[25]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[25]),
    .o(_al_u125_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u126 (
    .a(_al_u125_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[25]),
    .o(_al_u126_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u127 (
    .a(_al_u126_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[25]),
    .e(div_unsigned_quo[25]),
    .o(n42[25]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u128 (
    .a(n13[39]),
    .b(n11[39]),
    .c(n42[25]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[25]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u129 (
    .a(n44[25]),
    .b(n7[39]),
    .c(n7[7]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[25]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u130 (
    .a(n37[9]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[9]),
    .o(_al_u130_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u131 (
    .a(_al_u130_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[9]),
    .o(_al_u131_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u132 (
    .a(_al_u131_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[9]),
    .e(div_unsigned_quo[9]),
    .o(n42[9]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u133 (
    .a(n13[23]),
    .b(n11[23]),
    .c(n42[9]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[9]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u134 (
    .a(n44[9]),
    .b(n7[23]),
    .c(mult0_0_0_9),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[9]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u135 (
    .a(n37[20]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[20]),
    .o(_al_u135_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u136 (
    .a(_al_u135_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[20]),
    .o(_al_u136_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u137 (
    .a(_al_u136_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[20]),
    .e(div_unsigned_quo[20]),
    .o(n42[20]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u138 (
    .a(n13[34]),
    .b(n11[34]),
    .c(n42[20]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[20]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u139 (
    .a(n44[20]),
    .b(n7[34]),
    .c(n7[2]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[20]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u140 (
    .a(n37[18]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[18]),
    .o(_al_u140_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u141 (
    .a(_al_u140_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[18]),
    .o(_al_u141_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u142 (
    .a(_al_u141_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[18]),
    .e(div_unsigned_quo[18]),
    .o(n42[18]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u143 (
    .a(n13[32]),
    .b(n11[32]),
    .c(n42[18]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[18]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u144 (
    .a(n44[18]),
    .b(n7[32]),
    .c(n7[0]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[18]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u145 (
    .a(n37[23]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[23]),
    .o(_al_u145_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u146 (
    .a(_al_u145_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[23]),
    .o(_al_u146_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u147 (
    .a(_al_u146_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[23]),
    .e(div_unsigned_quo[23]),
    .o(n42[23]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u148 (
    .a(n13[37]),
    .b(n11[37]),
    .c(n42[23]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[23]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u149 (
    .a(n44[23]),
    .b(n7[37]),
    .c(n7[5]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[23]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u150 (
    .a(n37[17]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[17]),
    .o(_al_u150_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u151 (
    .a(_al_u150_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[17]),
    .o(_al_u151_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u152 (
    .a(_al_u151_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[17]),
    .e(div_unsigned_quo[17]),
    .o(n42[17]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u153 (
    .a(n13[31]),
    .b(n11[31]),
    .c(n42[17]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[17]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u154 (
    .a(n44[17]),
    .b(n7[31]),
    .c(mult0_0_0_17),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[17]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u155 (
    .a(n37[29]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[29]),
    .o(_al_u155_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u156 (
    .a(_al_u155_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[29]),
    .o(_al_u156_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u157 (
    .a(_al_u156_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[29]),
    .e(div_unsigned_quo[29]),
    .o(n42[29]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u158 (
    .a(n13[43]),
    .b(n11[43]),
    .c(n42[29]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[29]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u159 (
    .a(n44[29]),
    .b(n7[43]),
    .c(n7[11]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[29]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u160 (
    .a(n37[8]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[8]),
    .o(_al_u160_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u161 (
    .a(_al_u160_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[8]),
    .o(_al_u161_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u162 (
    .a(_al_u161_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[8]),
    .e(div_unsigned_quo[8]),
    .o(n42[8]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u163 (
    .a(n13[22]),
    .b(n11[22]),
    .c(n42[8]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[8]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u164 (
    .a(n44[8]),
    .b(n7[22]),
    .c(mult0_0_0_8),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[8]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u165 (
    .a(n37[16]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[16]),
    .o(_al_u165_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u166 (
    .a(_al_u165_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[16]),
    .o(_al_u166_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u167 (
    .a(_al_u166_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[16]),
    .e(div_unsigned_quo[16]),
    .o(n42[16]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u168 (
    .a(n13[30]),
    .b(n11[30]),
    .c(n42[16]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[16]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u169 (
    .a(n44[16]),
    .b(n7[30]),
    .c(mult0_0_0_16),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[16]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u170 (
    .a(n37[19]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[19]),
    .o(_al_u170_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u171 (
    .a(_al_u170_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[19]),
    .o(_al_u171_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u172 (
    .a(_al_u171_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[19]),
    .e(div_unsigned_quo[19]),
    .o(n42[19]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u173 (
    .a(n13[33]),
    .b(n11[33]),
    .c(n42[19]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[19]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u174 (
    .a(n44[19]),
    .b(n7[33]),
    .c(n7[1]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[19]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u175 (
    .a(n37[13]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[13]),
    .o(_al_u175_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u176 (
    .a(_al_u175_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[13]),
    .o(_al_u176_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u177 (
    .a(_al_u176_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[13]),
    .e(div_unsigned_quo[13]),
    .o(n42[13]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u178 (
    .a(n13[27]),
    .b(n11[27]),
    .c(n42[13]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[13]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u179 (
    .a(n44[13]),
    .b(n7[27]),
    .c(mult0_0_0_13),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[13]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u180 (
    .a(n37[10]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[10]),
    .o(_al_u180_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u181 (
    .a(_al_u180_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[10]),
    .o(_al_u181_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u182 (
    .a(_al_u181_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[10]),
    .e(div_unsigned_quo[10]),
    .o(n42[10]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u183 (
    .a(n13[24]),
    .b(n11[24]),
    .c(n42[10]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[10]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u184 (
    .a(n44[10]),
    .b(n7[24]),
    .c(mult0_0_0_10),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[10]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u185 (
    .a(n37[12]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[12]),
    .o(_al_u185_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u186 (
    .a(_al_u185_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[12]),
    .o(_al_u186_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u187 (
    .a(_al_u186_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[12]),
    .e(div_unsigned_quo[12]),
    .o(n42[12]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u188 (
    .a(n13[26]),
    .b(n11[26]),
    .c(n42[12]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[12]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u189 (
    .a(n44[12]),
    .b(n7[26]),
    .c(mult0_0_0_12),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[12]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u190 (
    .a(n37[15]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[15]),
    .o(_al_u190_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u191 (
    .a(_al_u190_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[15]),
    .o(_al_u191_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u192 (
    .a(_al_u191_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[15]),
    .e(div_unsigned_quo[15]),
    .o(n42[15]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u193 (
    .a(n13[29]),
    .b(n11[29]),
    .c(n42[15]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[15]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u194 (
    .a(n44[15]),
    .b(n7[29]),
    .c(mult0_0_0_15),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[15]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u195 (
    .a(n37[14]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[14]),
    .o(_al_u195_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u196 (
    .a(_al_u195_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[14]),
    .o(_al_u196_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u197 (
    .a(_al_u196_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[14]),
    .e(div_unsigned_quo[14]),
    .o(n42[14]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u198 (
    .a(n13[28]),
    .b(n11[28]),
    .c(n42[14]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[14]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u199 (
    .a(n44[14]),
    .b(n7[28]),
    .c(mult0_0_0_14),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[14]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u200 (
    .a(n37[21]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[21]),
    .o(_al_u200_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u201 (
    .a(_al_u200_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[21]),
    .o(_al_u201_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u202 (
    .a(_al_u201_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[21]),
    .e(div_unsigned_quo[21]),
    .o(n42[21]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u203 (
    .a(n13[35]),
    .b(n11[35]),
    .c(n42[21]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[21]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u204 (
    .a(n44[21]),
    .b(n7[35]),
    .c(n7[3]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[21]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u205 (
    .a(n37[22]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[22]),
    .o(_al_u205_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u206 (
    .a(_al_u205_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[22]),
    .o(_al_u206_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u207 (
    .a(_al_u206_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[22]),
    .e(div_unsigned_quo[22]),
    .o(n42[22]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u208 (
    .a(n13[36]),
    .b(n11[36]),
    .c(n42[22]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[22]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u209 (
    .a(n44[22]),
    .b(n7[36]),
    .c(n7[4]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[22]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u210 (
    .a(n37[26]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[26]),
    .o(_al_u210_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u211 (
    .a(_al_u210_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[26]),
    .o(_al_u211_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u212 (
    .a(_al_u211_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[26]),
    .e(div_unsigned_quo[26]),
    .o(n42[26]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u213 (
    .a(n13[40]),
    .b(n11[40]),
    .c(n42[26]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[26]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u214 (
    .a(n44[26]),
    .b(n7[40]),
    .c(n7[8]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[26]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u215 (
    .a(n37[28]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[28]),
    .o(_al_u215_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u216 (
    .a(_al_u215_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[28]),
    .o(_al_u216_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u217 (
    .a(_al_u216_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[28]),
    .e(div_unsigned_quo[28]),
    .o(n42[28]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u218 (
    .a(n13[42]),
    .b(n11[42]),
    .c(n42[28]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[28]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u219 (
    .a(n44[28]),
    .b(n7[42]),
    .c(n7[10]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[28]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u220 (
    .a(n37[30]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[30]),
    .o(_al_u220_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u221 (
    .a(_al_u220_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[30]),
    .o(_al_u221_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u222 (
    .a(_al_u221_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[30]),
    .e(div_unsigned_quo[30]),
    .o(n42[30]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u223 (
    .a(n13[44]),
    .b(n11[44]),
    .c(n42[30]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[30]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u224 (
    .a(n44[30]),
    .b(n7[44]),
    .c(n7[12]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[30]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u225 (
    .a(n37[24]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[24]),
    .o(_al_u225_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u226 (
    .a(_al_u225_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[24]),
    .o(_al_u226_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u227 (
    .a(_al_u226_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[24]),
    .e(div_unsigned_quo[24]),
    .o(n42[24]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u228 (
    .a(n13[38]),
    .b(n11[38]),
    .c(n42[24]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[24]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u229 (
    .a(n44[24]),
    .b(n7[38]),
    .c(n7[6]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[24]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u230 (
    .a(n37[31]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[31]),
    .o(_al_u230_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u231 (
    .a(_al_u230_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[31]),
    .o(_al_u231_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u232 (
    .a(_al_u231_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[31]),
    .e(div_unsigned_quo[31]),
    .o(n42[31]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u233 (
    .a(n13[45]),
    .b(n11[45]),
    .c(n42[31]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[31]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u234 (
    .a(n44[31]),
    .b(n7[45]),
    .c(n7[13]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[31]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u235 (
    .a(n37[27]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[27]),
    .o(_al_u235_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u236 (
    .a(_al_u235_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[27]),
    .o(_al_u236_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u237 (
    .a(_al_u236_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[27]),
    .e(div_unsigned_quo[27]),
    .o(n42[27]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u238 (
    .a(n13[41]),
    .b(n11[41]),
    .c(n42[27]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[27]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u239 (
    .a(n44[27]),
    .b(n7[41]),
    .c(n7[9]),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[27]));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*A*~(~E*~D))"),
    .INIT(32'h20202000))
    _al_u240 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mduinfo[8]),
    .e(i_mduinfo[6]),
    .o(div_unsigned_start));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*A*~(~E*~D))"),
    .INIT(32'h20202000))
    _al_u241 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mduinfo[7]),
    .e(i_mduinfo[5]),
    .o(div_signed_start));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u242 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[31]),
    .o(n35[31]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u243 (
    .a(mul_finish),
    .b(rem_op1_sym),
    .c(div_signed_finish),
    .d(div_unsigned_finish),
    .o(n5_lutinv));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E)*~((D*~B*A))+C*E*~((D*~B*A))+~(C)*E*(D*~B*A)+C*E*(D*~B*A))"),
    .INIT(32'hf2f0d0f0))
    _al_u244 (
    .a(i_vld),
    .b(o_working),
    .c(n5_lutinv),
    .d(i_decinfo_grp[3]),
    .e(i_mdu_op1[31]),
    .o(n10));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C*A))"),
    .INIT(8'hec))
    _al_u245 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .o(n8));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*~A)"),
    .INIT(32'h00000010))
    _al_u246 (
    .a(i_flush),
    .b(mul_finish),
    .c(o_will_rdwen),
    .d(div_signed_finish),
    .e(div_unsigned_finish),
    .o(n3_lutinv));
  AL_MAP_LUT5 #(
    .EQN("(B*~(E)*~((D*~C*A))+B*E*~((D*~C*A))+~(B)*E*(D*~C*A)+B*E*(D*~C*A))"),
    .INIT(32'hceccc4cc))
    _al_u247 (
    .a(i_vld),
    .b(n3_lutinv),
    .c(o_working),
    .d(i_decinfo_grp[3]),
    .e(i_mdu_rdwen),
    .o(n6));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u248 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_rstn),
    .o(mux2_b0_sel_is_2_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u249 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[9]),
    .o(n35[9]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u250 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[8]),
    .o(n35[8]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u251 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[7]),
    .o(n35[7]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u252 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[6]),
    .o(n35[6]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u253 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[5]),
    .o(n35[5]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u254 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[4]),
    .o(n35[4]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u255 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[30]),
    .o(n35[30]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u256 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[3]),
    .o(n35[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u257 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[29]),
    .o(n35[29]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u258 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[28]),
    .o(n35[28]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u259 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[27]),
    .o(n35[27]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u260 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[26]),
    .o(n35[26]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u261 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[25]),
    .o(n35[25]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u262 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[24]),
    .o(n35[24]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u263 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[23]),
    .o(n35[23]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u264 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[22]),
    .o(n35[22]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u265 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[21]),
    .o(n35[21]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u266 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[20]),
    .o(n35[20]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u267 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[2]),
    .o(n35[2]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u268 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[19]),
    .o(n35[19]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u269 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[18]),
    .o(n35[18]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u270 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[17]),
    .o(n35[17]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u271 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[16]),
    .o(n35[16]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u272 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[15]),
    .o(n35[15]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u273 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[14]),
    .o(n35[14]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u274 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[13]),
    .o(n35[13]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u275 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[12]),
    .o(n35[12]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u276 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[11]),
    .o(n35[11]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u277 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[10]),
    .o(n35[10]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u278 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[1]),
    .o(n35[1]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u279 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op1[0]),
    .o(n35[0]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u280 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[9]),
    .o(n34[9]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u281 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[8]),
    .o(n34[8]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u282 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[7]),
    .o(n34[7]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u283 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[6]),
    .o(n34[6]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u284 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[5]),
    .o(n34[5]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u285 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[4]),
    .o(n34[4]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u286 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[31]),
    .o(n34[31]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u287 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[30]),
    .o(n34[30]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u288 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[3]),
    .o(n34[3]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u289 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[29]),
    .o(n34[29]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u290 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[28]),
    .o(n34[28]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u291 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[27]),
    .o(n34[27]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u292 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[26]),
    .o(n34[26]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u293 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[25]),
    .o(n34[25]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u294 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[24]),
    .o(n34[24]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u295 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[23]),
    .o(n34[23]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u296 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[22]),
    .o(n34[22]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u297 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[21]),
    .o(n34[21]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u298 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[20]),
    .o(n34[20]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u299 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[2]),
    .o(n34[2]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u300 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[19]),
    .o(n34[19]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u301 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[18]),
    .o(n34[18]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u302 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[17]),
    .o(n34[17]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u303 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[16]),
    .o(n34[16]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u304 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[15]),
    .o(n34[15]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u305 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[14]),
    .o(n34[14]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u306 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[13]),
    .o(n34[13]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u307 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[12]),
    .o(n34[12]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u308 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[11]),
    .o(n34[11]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u309 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[10]),
    .o(n34[10]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u310 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[1]),
    .o(n34[1]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u311 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .d(i_mdu_op2[0]),
    .o(n34[0]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u312 (
    .a(cnt[4]),
    .b(cnt[5]),
    .c(cnt[6]),
    .d(cnt[7]),
    .o(_al_u312_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    _al_u313 (
    .a(_al_u312_o),
    .b(cnt[0]),
    .c(cnt[1]),
    .d(cnt[2]),
    .e(cnt[3]),
    .o(_al_u313_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u314 (
    .a(_al_u313_o),
    .b(mul_vld),
    .o(n24_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u315 (
    .a(i_mduinfo[4]),
    .b(i_mduinfo[3]),
    .c(i_mduinfo[2]),
    .d(i_mduinfo[1]),
    .o(_al_u315_o));
  AL_MAP_LUT5 #(
    .EQN("~(~B*~(E*~D*~C*A))"),
    .INIT(32'hcccecccc))
    _al_u316 (
    .a(i_vld),
    .b(n24_lutinv),
    .c(_al_u315_o),
    .d(o_working),
    .e(i_decinfo_grp[3]),
    .o(n26));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((B*~A))*~(C)+D*(B*~A)*~(C)+~(D)*(B*~A)*C+D*(B*~A)*C)"),
    .INIT(16'hb0bf))
    _al_u317 (
    .a(_al_u313_o),
    .b(n19[7]),
    .c(mul_vld),
    .d(cnt[7]),
    .o(_al_u317_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~D*~C*A))"),
    .INIT(32'h33313333))
    _al_u318 (
    .a(i_vld),
    .b(_al_u317_o),
    .c(_al_u315_o),
    .d(o_working),
    .e(i_decinfo_grp[3]),
    .o(n29[7]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((B*~A))*~(C)+D*(B*~A)*~(C)+~(D)*(B*~A)*C+D*(B*~A)*C)"),
    .INIT(16'hb0bf))
    _al_u319 (
    .a(_al_u313_o),
    .b(n19[6]),
    .c(mul_vld),
    .d(cnt[6]),
    .o(_al_u319_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~D*~C*A))"),
    .INIT(32'h33313333))
    _al_u320 (
    .a(i_vld),
    .b(_al_u319_o),
    .c(_al_u315_o),
    .d(o_working),
    .e(i_decinfo_grp[3]),
    .o(n29[6]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((B*~A))*~(C)+D*(B*~A)*~(C)+~(D)*(B*~A)*C+D*(B*~A)*C)"),
    .INIT(16'hb0bf))
    _al_u321 (
    .a(_al_u313_o),
    .b(n19[5]),
    .c(mul_vld),
    .d(cnt[5]),
    .o(_al_u321_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~D*~C*A))"),
    .INIT(32'h33313333))
    _al_u322 (
    .a(i_vld),
    .b(_al_u321_o),
    .c(_al_u315_o),
    .d(o_working),
    .e(i_decinfo_grp[3]),
    .o(n29[5]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((B*~A))*~(C)+D*(B*~A)*~(C)+~(D)*(B*~A)*C+D*(B*~A)*C)"),
    .INIT(16'hb0bf))
    _al_u323 (
    .a(_al_u313_o),
    .b(n19[4]),
    .c(mul_vld),
    .d(cnt[4]),
    .o(_al_u323_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~D*~C*A))"),
    .INIT(32'h33313333))
    _al_u324 (
    .a(i_vld),
    .b(_al_u323_o),
    .c(_al_u315_o),
    .d(o_working),
    .e(i_decinfo_grp[3]),
    .o(n29[4]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((B*~A))*~(C)+D*(B*~A)*~(C)+~(D)*(B*~A)*C+D*(B*~A)*C)"),
    .INIT(16'hb0bf))
    _al_u325 (
    .a(_al_u313_o),
    .b(n19[3]),
    .c(mul_vld),
    .d(cnt[3]),
    .o(_al_u325_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~D*~C*A))"),
    .INIT(32'h33313333))
    _al_u326 (
    .a(i_vld),
    .b(_al_u325_o),
    .c(_al_u315_o),
    .d(o_working),
    .e(i_decinfo_grp[3]),
    .o(n29[3]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((B*~A))*~(C)+D*(B*~A)*~(C)+~(D)*(B*~A)*C+D*(B*~A)*C)"),
    .INIT(16'hb0bf))
    _al_u327 (
    .a(_al_u313_o),
    .b(n19[2]),
    .c(mul_vld),
    .d(cnt[2]),
    .o(_al_u327_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~D*~C*A))"),
    .INIT(32'h33313333))
    _al_u328 (
    .a(i_vld),
    .b(_al_u327_o),
    .c(_al_u315_o),
    .d(o_working),
    .e(i_decinfo_grp[3]),
    .o(n29[2]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((B*~A))*~(C)+D*(B*~A)*~(C)+~(D)*(B*~A)*C+D*(B*~A)*C)"),
    .INIT(16'hb0bf))
    _al_u329 (
    .a(_al_u313_o),
    .b(n19[1]),
    .c(mul_vld),
    .d(cnt[1]),
    .o(_al_u329_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~D*~C*A))"),
    .INIT(32'h33313333))
    _al_u330 (
    .a(i_vld),
    .b(_al_u329_o),
    .c(_al_u315_o),
    .d(o_working),
    .e(i_decinfo_grp[3]),
    .o(n29[1]));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((B*~A))*~(C)+D*(B*~A)*~(C)+~(D)*(B*~A)*C+D*(B*~A)*C)"),
    .INIT(16'hb0bf))
    _al_u331 (
    .a(_al_u313_o),
    .b(n19[0]),
    .c(mul_vld),
    .d(cnt[0]),
    .o(_al_u331_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~D*~C*A))"),
    .INIT(32'h33313333))
    _al_u332 (
    .a(i_vld),
    .b(_al_u331_o),
    .c(_al_u315_o),
    .d(o_working),
    .e(i_decinfo_grp[3]),
    .o(n29[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u333 (
    .a(mux2_b0_sel_is_2_o),
    .b(_al_u315_o),
    .o(mux10_b0_sel_is_2_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u334 (
    .a(_al_u313_o),
    .b(mul_finish),
    .c(mul_vld),
    .o(_al_u334_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(E*~D*~C*A))"),
    .INIT(32'hccc4cccc))
    _al_u335 (
    .a(i_vld),
    .b(_al_u334_o),
    .c(_al_u315_o),
    .d(o_working),
    .e(i_decinfo_grp[3]),
    .o(n30));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~C*~A))"),
    .INIT(16'hccc8))
    _al_u76 (
    .a(mul_finish),
    .b(o_will_rdwen),
    .c(div_signed_finish),
    .d(div_unsigned_finish),
    .o(o_mdu_rdwen));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u77 (
    .a(mul_finish),
    .b(div_signed_finish),
    .c(div_unsigned_finish),
    .d(working),
    .o(o_working));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u78 (
    .a(i_vld),
    .b(o_working),
    .c(i_decinfo_grp[3]),
    .o(mdu_vld));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u79 (
    .a(n37[2]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[2]),
    .o(_al_u79_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u80 (
    .a(mduinfo[7]),
    .b(mduinfo[8]),
    .o(_al_u80_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u81 (
    .a(_al_u79_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[2]),
    .o(_al_u81_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u82 (
    .a(_al_u81_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[2]),
    .e(div_unsigned_quo[2]),
    .o(n42[2]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u83 (
    .a(n13[16]),
    .b(n11[16]),
    .c(n42[2]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[2]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u84 (
    .a(n44[2]),
    .b(n7[16]),
    .c(mult0_0_0_2),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[2]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u85 (
    .a(n37[0]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[0]),
    .o(_al_u85_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u86 (
    .a(_al_u85_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[0]),
    .o(_al_u86_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u87 (
    .a(_al_u86_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[0]),
    .e(div_unsigned_quo[0]),
    .o(n42[0]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u88 (
    .a(n13[14]),
    .b(n11[14]),
    .c(n42[0]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[0]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u89 (
    .a(n44[0]),
    .b(n7[14]),
    .c(mult0_0_0_0),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[0]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u90 (
    .a(n37[7]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[7]),
    .o(_al_u90_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u91 (
    .a(_al_u90_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[7]),
    .o(_al_u91_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u92 (
    .a(_al_u91_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[7]),
    .e(div_unsigned_quo[7]),
    .o(n42[7]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u93 (
    .a(n13[21]),
    .b(n11[21]),
    .c(n42[7]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[7]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u94 (
    .a(n44[7]),
    .b(n7[21]),
    .c(mult0_0_0_7),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[7]));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(A)*~(C)+D*A*~(C)+~(D)*A*C+D*A*C))"),
    .INIT(16'h8c80))
    _al_u95 (
    .a(n37[3]),
    .b(mduinfo[7]),
    .c(rem_op1_sym),
    .d(div_signed_rem[3]),
    .o(_al_u95_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u96 (
    .a(_al_u95_o),
    .b(_al_u80_o),
    .c(div_unsigned_rem[3]),
    .o(_al_u96_o));
  AL_MAP_LUT5 #(
    .EQN("((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*~(D)*~(B)+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*~(B)+~((~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C))*D*B+(~A*~(E)*~(C)+~A*E*~(C)+~(~A)*E*C+~A*E*C)*D*B)"),
    .INIT(32'hfd31cd01))
    _al_u97 (
    .a(_al_u96_o),
    .b(mduinfo[5]),
    .c(mduinfo[6]),
    .d(div_signed_quo[3]),
    .e(div_unsigned_quo[3]),
    .o(n42[3]));
  AL_MAP_LUT5 #(
    .EQN("((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*~(B)*~(E)+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*~(E)+~((C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))*B*E+(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D)*B*E)"),
    .INIT(32'hccccaaf0))
    _al_u98 (
    .a(n13[17]),
    .b(n11[17]),
    .c(n42[3]),
    .d(mduinfo[3]),
    .e(mduinfo[4]),
    .o(n44[3]));
  AL_MAP_LUT5 #(
    .EQN("((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*~(C)*~(D)+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*~(D)+~((A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E))*C*D+(A*~(B)*~(E)+A*B*~(E)+~(A)*B*E+A*B*E)*C*D)"),
    .INIT(32'hf0ccf0aa))
    _al_u99 (
    .a(n44[3]),
    .b(n7[17]),
    .c(mult0_0_0_3),
    .d(mduinfo[1]),
    .e(mduinfo[2]),
    .o(o_mdu_rdwdata[3]));
  EG_PHY_MSLICE #(
    //.MACRO("add0/u0|add0/ucin"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \add0/u0|add0/ucin  (
    .a({cnt[0],1'b0}),
    .b({1'b1,open_n0}),
    .f({n19[0],open_n20}),
    .fco(\add0/c1 ));
  EG_PHY_MSLICE #(
    //.MACRO("add0/u0|add0/ucin"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \add0/u2|add0/u1  (
    .a(cnt[2:1]),
    .b(2'b00),
    .fci(\add0/c1 ),
    .f(n19[2:1]),
    .fco(\add0/c3 ));
  EG_PHY_MSLICE #(
    //.MACRO("add0/u0|add0/ucin"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \add0/u4|add0/u3  (
    .a(cnt[4:3]),
    .b(2'b00),
    .fci(\add0/c3 ),
    .f(n19[4:3]),
    .fco(\add0/c5 ));
  EG_PHY_MSLICE #(
    //.MACRO("add0/u0|add0/ucin"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \add0/u6|add0/u5  (
    .a(cnt[6:5]),
    .b(2'b00),
    .fci(\add0/c5 ),
    .f(n19[6:5]),
    .fco(\add0/c7 ));
  EG_PHY_MSLICE #(
    //.MACRO("add0/u0|add0/ucin"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \add0/u7_al_u423  (
    .a({open_n91,cnt[7]}),
    .b({open_n92,1'b0}),
    .fci(\add0/c7 ),
    .f({open_n111,n19[7]}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    mul_finish_reg (
    .clk(i_clk),
    .d(n30),
    .sr(i_rstn),
    .q(mul_finish));  // ../RTL/core/exu_mdu.v(96)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    mul_vld_reg (
    .clk(i_clk),
    .d(n26),
    .sr(i_rstn),
    .q(mul_vld));  // ../RTL/core/exu_mdu.v(96)
  EG_PHY_MULT18 #(
    .CEAMUX("SIG"),
    .CEBMUX("SIG"),
    .CLKMUX("SIG"),
    .INPUTREGA("ENABLE"),
    .INPUTREGB("ENABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .RSTANMUX("1"),
    .RSTBNMUX("1"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    mult0_0_0_ (
    .a(i_mdu_op1[17:0]),
    .b(i_mdu_op2[17:0]),
    .cea(mux10_b0_sel_is_2_o),
    .ceb(mux10_b0_sel_is_2_o),
    .clk(i_clk),
    .p({mult0_0_0_35,mult0_0_0_34,mult0_0_0_33,mult0_0_0_32,mult0_0_0_31,mult0_0_0_30,mult0_0_0_29,mult0_0_0_28,mult0_0_0_27,mult0_0_0_26,mult0_0_0_25,mult0_0_0_24,mult0_0_0_23,mult0_0_0_22,mult0_0_0_21,mult0_0_0_20,mult0_0_0_19,mult0_0_0_18,mult0_0_0_17,mult0_0_0_16,mult0_0_0_15,mult0_0_0_14,mult0_0_0_13,mult0_0_0_12,mult0_0_0_11,mult0_0_0_10,mult0_0_0_9,mult0_0_0_8,mult0_0_0_7,mult0_0_0_6,mult0_0_0_5,mult0_0_0_4,mult0_0_0_3,mult0_0_0_2,mult0_0_0_1,mult0_0_0_0}));
  EG_PHY_MULT18 #(
    .CEAMUX("SIG"),
    .CEBMUX("SIG"),
    .CLKMUX("SIG"),
    .INPUTREGA("ENABLE"),
    .INPUTREGB("ENABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .RSTANMUX("1"),
    .RSTBNMUX("1"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("1"))
    mult0_0_1_ (
    .a(i_mdu_op1[17:0]),
    .b({i_mdu_op2[31],i_mdu_op2[31],i_mdu_op2[31],i_mdu_op2[31],i_mdu_op2[31:18]}),
    .cea(mux10_b0_sel_is_2_o),
    .ceb(mux10_b0_sel_is_2_o),
    .clk(i_clk),
    .p({open_n279,open_n280,open_n281,open_n282,mult0_0_1_31,mult0_0_1_30,mult0_0_1_29,mult0_0_1_28,mult0_0_1_27,mult0_0_1_26,mult0_0_1_25,mult0_0_1_24,mult0_0_1_23,mult0_0_1_22,mult0_0_1_21,mult0_0_1_20,mult0_0_1_19,mult0_0_1_18,mult0_0_1_17,mult0_0_1_16,mult0_0_1_15,mult0_0_1_14,mult0_0_1_13,mult0_0_1_12,mult0_0_1_11,mult0_0_1_10,mult0_0_1_9,mult0_0_1_8,mult0_0_1_7,mult0_0_1_6,mult0_0_1_5,mult0_0_1_4,mult0_0_1_3,mult0_0_1_2,mult0_0_1_1,mult0_0_1_0}));
  EG_PHY_MULT18 #(
    .CEAMUX("SIG"),
    .CEBMUX("SIG"),
    .CLKMUX("SIG"),
    .INPUTREGA("ENABLE"),
    .INPUTREGB("ENABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .RSTANMUX("1"),
    .RSTBNMUX("1"),
    .SIGNEDAMUX("1"),
    .SIGNEDBMUX("0"))
    mult0_1_0_ (
    .a({i_mdu_op1[31],i_mdu_op1[31],i_mdu_op1[31],i_mdu_op1[31],i_mdu_op1[31:18]}),
    .b(i_mdu_op2[17:0]),
    .cea(mux10_b0_sel_is_2_o),
    .ceb(mux10_b0_sel_is_2_o),
    .clk(i_clk),
    .p({open_n363,open_n364,open_n365,open_n366,mult0_1_0_31,mult0_1_0_30,mult0_1_0_29,mult0_1_0_28,mult0_1_0_27,mult0_1_0_26,mult0_1_0_25,mult0_1_0_24,mult0_1_0_23,mult0_1_0_22,mult0_1_0_21,mult0_1_0_20,mult0_1_0_19,mult0_1_0_18,mult0_1_0_17,mult0_1_0_16,mult0_1_0_15,mult0_1_0_14,mult0_1_0_13,mult0_1_0_12,mult0_1_0_11,mult0_1_0_10,mult0_1_0_9,mult0_1_0_8,mult0_1_0_7,mult0_1_0_6,mult0_1_0_5,mult0_1_0_4,mult0_1_0_3,mult0_1_0_2,mult0_1_0_1,mult0_1_0_0}));
  EG_PHY_MULT18 #(
    .CEAMUX("SIG"),
    .CEBMUX("SIG"),
    .CLKMUX("SIG"),
    .INPUTREGA("ENABLE"),
    .INPUTREGB("ENABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .RSTANMUX("1"),
    .RSTBNMUX("1"),
    .SIGNEDAMUX("1"),
    .SIGNEDBMUX("1"))
    mult0_1_1_ (
    .a({i_mdu_op1[31],i_mdu_op1[31],i_mdu_op1[31],i_mdu_op1[31],i_mdu_op1[31:18]}),
    .b({i_mdu_op2[31],i_mdu_op2[31],i_mdu_op2[31],i_mdu_op2[31],i_mdu_op2[31:18]}),
    .cea(mux10_b0_sel_is_2_o),
    .ceb(mux10_b0_sel_is_2_o),
    .clk(i_clk),
    .p({open_n447,open_n448,open_n449,open_n450,open_n451,open_n452,open_n453,open_n454,mult0_1_1_27,mult0_1_1_26,mult0_1_1_25,mult0_1_1_24,mult0_1_1_23,mult0_1_1_22,mult0_1_1_21,mult0_1_1_20,mult0_1_1_19,mult0_1_1_18,mult0_1_1_17,mult0_1_1_16,mult0_1_1_15,mult0_1_1_14,mult0_1_1_13,mult0_1_1_12,mult0_1_1_11,mult0_1_1_10,mult0_1_1_9,mult0_1_1_8,mult0_1_1_7,mult0_1_1_6,mult0_1_1_5,mult0_1_1_4,mult0_1_1_3,mult0_1_1_2,mult0_1_1_1,mult0_1_1_0}));
  EG_PHY_MULT18 #(
    .CEAMUX("SIG"),
    .CEBMUX("SIG"),
    .CLKMUX("SIG"),
    .INPUTREGA("ENABLE"),
    .INPUTREGB("ENABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .RSTANMUX("1"),
    .RSTBNMUX("1"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    mult1_0_1_ (
    .a(i_mdu_op1[17:0]),
    .b({4'b0000,i_mdu_op2[31:18]}),
    .cea(mux10_b0_sel_is_2_o),
    .ceb(mux10_b0_sel_is_2_o),
    .clk(i_clk),
    .p({open_n535,open_n536,open_n537,open_n538,mult1_0_1_31,mult1_0_1_30,mult1_0_1_29,mult1_0_1_28,mult1_0_1_27,mult1_0_1_26,mult1_0_1_25,mult1_0_1_24,mult1_0_1_23,mult1_0_1_22,mult1_0_1_21,mult1_0_1_20,mult1_0_1_19,mult1_0_1_18,mult1_0_1_17,mult1_0_1_16,mult1_0_1_15,mult1_0_1_14,mult1_0_1_13,mult1_0_1_12,mult1_0_1_11,mult1_0_1_10,mult1_0_1_9,mult1_0_1_8,mult1_0_1_7,mult1_0_1_6,mult1_0_1_5,mult1_0_1_4,mult1_0_1_3,mult1_0_1_2,mult1_0_1_1,mult1_0_1_0}));
  EG_PHY_MULT18 #(
    .CEAMUX("SIG"),
    .CEBMUX("SIG"),
    .CLKMUX("SIG"),
    .INPUTREGA("ENABLE"),
    .INPUTREGB("ENABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .RSTANMUX("1"),
    .RSTBNMUX("1"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    mult1_1_0_ (
    .a({4'b0000,i_mdu_op1[31:18]}),
    .b(i_mdu_op2[17:0]),
    .cea(mux10_b0_sel_is_2_o),
    .ceb(mux10_b0_sel_is_2_o),
    .clk(i_clk),
    .p({open_n619,open_n620,open_n621,open_n622,mult1_1_0_31,mult1_1_0_30,mult1_1_0_29,mult1_1_0_28,mult1_1_0_27,mult1_1_0_26,mult1_1_0_25,mult1_1_0_24,mult1_1_0_23,mult1_1_0_22,mult1_1_0_21,mult1_1_0_20,mult1_1_0_19,mult1_1_0_18,mult1_1_0_17,mult1_1_0_16,mult1_1_0_15,mult1_1_0_14,mult1_1_0_13,mult1_1_0_12,mult1_1_0_11,mult1_1_0_10,mult1_1_0_9,mult1_1_0_8,mult1_1_0_7,mult1_1_0_6,mult1_1_0_5,mult1_1_0_4,mult1_1_0_3,mult1_1_0_2,mult1_1_0_1,mult1_1_0_0}));
  EG_PHY_MULT18 #(
    .CEAMUX("SIG"),
    .CEBMUX("SIG"),
    .CLKMUX("SIG"),
    .INPUTREGA("ENABLE"),
    .INPUTREGB("ENABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .RSTANMUX("1"),
    .RSTBNMUX("1"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("0"))
    mult1_1_1_ (
    .a({4'b0000,i_mdu_op1[31:18]}),
    .b({4'b0000,i_mdu_op2[31:18]}),
    .cea(mux10_b0_sel_is_2_o),
    .ceb(mux10_b0_sel_is_2_o),
    .clk(i_clk),
    .p({open_n703,open_n704,open_n705,open_n706,open_n707,open_n708,open_n709,open_n710,mult1_1_1_27,mult1_1_1_26,mult1_1_1_25,mult1_1_1_24,mult1_1_1_23,mult1_1_1_22,mult1_1_1_21,mult1_1_1_20,mult1_1_1_19,mult1_1_1_18,mult1_1_1_17,mult1_1_1_16,mult1_1_1_15,mult1_1_1_14,mult1_1_1_13,mult1_1_1_12,mult1_1_1_11,mult1_1_1_10,mult1_1_1_9,mult1_1_1_8,mult1_1_1_7,mult1_1_1_6,mult1_1_1_5,mult1_1_1_4,mult1_1_1_3,mult1_1_1_2,mult1_1_1_1,mult1_1_1_0}));
  EG_PHY_MULT18 #(
    .CEAMUX("SIG"),
    .CEBMUX("SIG"),
    .CLKMUX("SIG"),
    .INPUTREGA("ENABLE"),
    .INPUTREGB("ENABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .RSTANMUX("1"),
    .RSTBNMUX("1"),
    .SIGNEDAMUX("0"),
    .SIGNEDBMUX("1"))
    mult2_0_1_ (
    .a(i_mdu_op1[17:0]),
    .b({4'b0000,i_mdu_op2[31:18]}),
    .cea(mux10_b0_sel_is_2_o),
    .ceb(mux10_b0_sel_is_2_o),
    .clk(i_clk),
    .p({open_n791,open_n792,open_n793,mult2_0_1_32,mult2_0_1_31,mult2_0_1_30,mult2_0_1_29,mult2_0_1_28,mult2_0_1_27,mult2_0_1_26,mult2_0_1_25,mult2_0_1_24,mult2_0_1_23,mult2_0_1_22,mult2_0_1_21,mult2_0_1_20,mult2_0_1_19,mult2_0_1_18,mult2_0_1_17,mult2_0_1_16,mult2_0_1_15,mult2_0_1_14,mult2_0_1_13,mult2_0_1_12,mult2_0_1_11,mult2_0_1_10,mult2_0_1_9,mult2_0_1_8,mult2_0_1_7,mult2_0_1_6,mult2_0_1_5,mult2_0_1_4,mult2_0_1_3,mult2_0_1_2,mult2_0_1_1,mult2_0_1_0}));
  EG_PHY_MULT18 #(
    .CEAMUX("SIG"),
    .CEBMUX("SIG"),
    .CLKMUX("SIG"),
    .INPUTREGA("ENABLE"),
    .INPUTREGB("ENABLE"),
    .MODE("MULT18X18C"),
    .OUTPUTREG("DISABLE"),
    .RSTANMUX("1"),
    .RSTBNMUX("1"),
    .SIGNEDAMUX("1"),
    .SIGNEDBMUX("1"))
    mult2_1_1_ (
    .a({i_mdu_op1[31],i_mdu_op1[31],i_mdu_op1[31],i_mdu_op1[31],i_mdu_op1[31:18]}),
    .b({4'b0000,i_mdu_op2[31:18]}),
    .cea(mux10_b0_sel_is_2_o),
    .ceb(mux10_b0_sel_is_2_o),
    .clk(i_clk),
    .p({open_n874,open_n875,open_n876,open_n877,open_n878,open_n879,open_n880,open_n881,mult2_1_1_27,mult2_1_1_26,mult2_1_1_25,mult2_1_1_24,mult2_1_1_23,mult2_1_1_22,mult2_1_1_21,mult2_1_1_20,mult2_1_1_19,mult2_1_1_18,mult2_1_1_17,mult2_1_1_16,mult2_1_1_15,mult2_1_1_14,mult2_1_1_13,mult2_1_1_12,mult2_1_1_11,mult2_1_1_10,mult2_1_1_9,mult2_1_1_8,mult2_1_1_7,mult2_1_1_6,mult2_1_1_5,mult2_1_1_4,mult2_1_1_3,mult2_1_1_2,mult2_1_1_1,mult2_1_1_0}));
  EG_PHY_LSLICE #(
    //.MACRO("neg0/ucin_al_u405"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \neg0/u11_al_u408  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({div_signed_rem[13],div_signed_rem[11]}),
    .e({div_signed_rem[14],div_signed_rem[12]}),
    .fci(\neg0/c11 ),
    .f({n37[13],n37[11]}),
    .fco(\neg0/c15 ),
    .fx({n37[14],n37[12]}));
  EG_PHY_LSLICE #(
    //.MACRO("neg0/ucin_al_u405"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \neg0/u15_al_u409  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({div_signed_rem[17],div_signed_rem[15]}),
    .e({div_signed_rem[18],div_signed_rem[16]}),
    .fci(\neg0/c15 ),
    .f({n37[17],n37[15]}),
    .fco(\neg0/c19 ),
    .fx({n37[18],n37[16]}));
  EG_PHY_LSLICE #(
    //.MACRO("neg0/ucin_al_u405"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \neg0/u19_al_u410  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({div_signed_rem[21],div_signed_rem[19]}),
    .e({div_signed_rem[22],div_signed_rem[20]}),
    .fci(\neg0/c19 ),
    .f({n37[21],n37[19]}),
    .fco(\neg0/c23 ),
    .fx({n37[22],n37[20]}));
  EG_PHY_LSLICE #(
    //.MACRO("neg0/ucin_al_u405"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \neg0/u23_al_u411  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({div_signed_rem[25],div_signed_rem[23]}),
    .e({div_signed_rem[26],div_signed_rem[24]}),
    .fci(\neg0/c23 ),
    .f({n37[25],n37[23]}),
    .fco(\neg0/c27 ),
    .fx({n37[26],n37[24]}));
  EG_PHY_LSLICE #(
    //.MACRO("neg0/ucin_al_u405"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \neg0/u27_al_u412  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({div_signed_rem[29],div_signed_rem[27]}),
    .e({div_signed_rem[30],div_signed_rem[28]}),
    .fci(\neg0/c27 ),
    .f({n37[29],n37[27]}),
    .fco(\neg0/c31 ),
    .fx({n37[30],n37[28]}));
  EG_PHY_LSLICE #(
    //.MACRO("neg0/ucin_al_u405"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \neg0/u31_al_u413  (
    .a({open_n972,1'b0}),
    .c(2'b11),
    .d({open_n977,div_signed_rem[31]}),
    .fci(\neg0/c31 ),
    .f({open_n994,n37[31]}));
  EG_PHY_LSLICE #(
    //.MACRO("neg0/ucin_al_u405"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \neg0/u3_al_u406  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({div_signed_rem[5],div_signed_rem[3]}),
    .e({div_signed_rem[6],div_signed_rem[4]}),
    .fci(\neg0/c3 ),
    .f({n37[5],n37[3]}),
    .fco(\neg0/c7 ),
    .fx({n37[6],n37[4]}));
  EG_PHY_LSLICE #(
    //.MACRO("neg0/ucin_al_u405"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \neg0/u7_al_u407  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({div_signed_rem[9],div_signed_rem[7]}),
    .e({div_signed_rem[10],div_signed_rem[8]}),
    .fci(\neg0/c7 ),
    .f({n37[9],n37[7]}),
    .fco(\neg0/c11 ),
    .fx({n37[10],n37[8]}));
  EG_PHY_LSLICE #(
    //.MACRO("neg0/ucin_al_u405"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \neg0/ucin_al_u405  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b11),
    .d({div_signed_rem[1],1'b1}),
    .e({div_signed_rem[2],div_signed_rem[0]}),
    .f({n37[1],open_n1053}),
    .fco(\neg0/c3 ),
    .fx({n37[2],n37[0]}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    rdwen_reg (
    .clk(i_clk),
    .d(n6),
    .sr(i_rstn),
    .q(o_will_rdwen));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b0 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mdu_rdidx[0]),
    .q(o_will_rdidx[0]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b1 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mdu_rdidx[1]),
    .q(o_mdu_rdidx[1]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b2 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mdu_rdidx[2]),
    .q(o_mdu_rdidx[2]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b3 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mdu_rdidx[3]),
    .q(o_will_rdidx[3]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg0_b4 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mdu_rdidx[4]),
    .q(o_will_rdidx[4]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b1 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mduinfo[1]),
    .q(mduinfo[1]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b2 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mduinfo[2]),
    .q(mduinfo[2]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b3 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mduinfo[3]),
    .q(mduinfo[3]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b4 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mduinfo[4]),
    .q(mduinfo[4]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b5 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mduinfo[5]),
    .q(mduinfo[5]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b6 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mduinfo[6]),
    .q(mduinfo[6]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b7 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mduinfo[7]),
    .q(mduinfo[7]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    reg1_b8 (
    .ce(mux2_b0_sel_is_2_o),
    .clk(i_clk),
    .d(i_mduinfo[8]),
    .q(mduinfo[8]));  // ../RTL/core/exu_mdu.v(52)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b0 (
    .clk(i_clk),
    .d(n29[0]),
    .sr(i_rstn),
    .q(cnt[0]));  // ../RTL/core/exu_mdu.v(96)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b1 (
    .clk(i_clk),
    .d(n29[1]),
    .sr(i_rstn),
    .q(cnt[1]));  // ../RTL/core/exu_mdu.v(96)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b2 (
    .clk(i_clk),
    .d(n29[2]),
    .sr(i_rstn),
    .q(cnt[2]));  // ../RTL/core/exu_mdu.v(96)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b3 (
    .clk(i_clk),
    .d(n29[3]),
    .sr(i_rstn),
    .q(cnt[3]));  // ../RTL/core/exu_mdu.v(96)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b4 (
    .clk(i_clk),
    .d(n29[4]),
    .sr(i_rstn),
    .q(cnt[4]));  // ../RTL/core/exu_mdu.v(96)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b5 (
    .clk(i_clk),
    .d(n29[5]),
    .sr(i_rstn),
    .q(cnt[5]));  // ../RTL/core/exu_mdu.v(96)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b6 (
    .clk(i_clk),
    .d(n29[6]),
    .sr(i_rstn),
    .q(cnt[6]));  // ../RTL/core/exu_mdu.v(96)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    reg2_b7 (
    .clk(i_clk),
    .d(n29[7]),
    .sr(i_rstn),
    .q(cnt[7]));  // ../RTL/core/exu_mdu.v(96)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    rem_op1_sym_reg (
    .clk(i_clk),
    .d(n10),
    .sr(i_rstn),
    .q(rem_op1_sym));  // ../RTL/core/exu_mdu.v(52)
  EG_PHY_LSLICE #(
    //.MACRO("u1/ucin_al_u336"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1/u11_al_u339  (
    .a({mult0_1_0_13,mult0_1_0_11}),
    .b({mult0_1_0_14,mult0_1_0_12}),
    .c(2'b00),
    .d({mult0_0_0_31,mult0_0_0_29}),
    .e({mult0_0_0_32,mult0_0_0_30}),
    .fci(\u1/c11 ),
    .f({n2[13],n2[11]}),
    .fco(\u1/c15 ),
    .fx({n2[14],n2[12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1/ucin_al_u336"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1/u15_al_u340  (
    .a({mult0_1_0_17,mult0_1_0_15}),
    .b({mult0_1_0_18,mult0_1_0_16}),
    .c(2'b00),
    .d({mult0_0_0_35,mult0_0_0_33}),
    .e({mult0_1_1_0,mult0_0_0_34}),
    .fci(\u1/c15 ),
    .f({n2[17],n2[15]}),
    .fco(\u1/c19 ),
    .fx({n2[18],n2[16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1/ucin_al_u336"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1/u19_al_u341  (
    .a({mult0_1_0_21,mult0_1_0_19}),
    .b({mult0_1_0_22,mult0_1_0_20}),
    .c(2'b00),
    .d({mult0_1_1_3,mult0_1_1_1}),
    .e({mult0_1_1_4,mult0_1_1_2}),
    .fci(\u1/c19 ),
    .f({n2[21],n2[19]}),
    .fco(\u1/c23 ),
    .fx({n2[22],n2[20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1/ucin_al_u336"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1/u23_al_u342  (
    .a({mult0_1_0_25,mult0_1_0_23}),
    .b({mult0_1_0_26,mult0_1_0_24}),
    .c(2'b00),
    .d({mult0_1_1_7,mult0_1_1_5}),
    .e({mult0_1_1_8,mult0_1_1_6}),
    .fci(\u1/c23 ),
    .f({n2[25],n2[23]}),
    .fco(\u1/c27 ),
    .fx({n2[26],n2[24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1/ucin_al_u336"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1/u27_al_u343  (
    .a({mult0_1_0_29,mult0_1_0_27}),
    .b({mult0_1_0_30,mult0_1_0_28}),
    .c(2'b00),
    .d({mult0_1_1_11,mult0_1_1_9}),
    .e({mult0_1_1_12,mult0_1_1_10}),
    .fci(\u1/c27 ),
    .f({n2[29],n2[27]}),
    .fco(\u1/c31 ),
    .fx({n2[30],n2[28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1/ucin_al_u336"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1/u31_al_u344  (
    .a({mult0_1_0_31,mult0_1_0_31}),
    .b({mult0_1_0_31,mult0_1_0_31}),
    .c(2'b00),
    .d({mult0_1_1_15,mult0_1_1_13}),
    .e({mult0_1_1_16,mult0_1_1_14}),
    .fci(\u1/c31 ),
    .f({n2[33],n2[31]}),
    .fco(\u1/c35 ),
    .fx({n2[34],n2[32]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1/ucin_al_u336"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1/u35_al_u345  (
    .a({mult0_1_0_31,mult0_1_0_31}),
    .b({mult0_1_0_31,mult0_1_0_31}),
    .c(2'b00),
    .d({mult0_1_1_19,mult0_1_1_17}),
    .e({mult0_1_1_20,mult0_1_1_18}),
    .fci(\u1/c35 ),
    .f({n2[37],n2[35]}),
    .fco(\u1/c39 ),
    .fx({n2[38],n2[36]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1/ucin_al_u336"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1/u39_al_u346  (
    .a({mult0_1_0_31,mult0_1_0_31}),
    .b({mult0_1_0_31,mult0_1_0_31}),
    .c(2'b00),
    .d({mult0_1_1_23,mult0_1_1_21}),
    .e({mult0_1_1_24,mult0_1_1_22}),
    .fci(\u1/c39 ),
    .f({n2[41],n2[39]}),
    .fco(\u1/c43 ),
    .fx({n2[42],n2[40]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1/ucin_al_u336"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1/u3_al_u337  (
    .a({mult0_1_0_5,mult0_1_0_3}),
    .b({mult0_1_0_6,mult0_1_0_4}),
    .c(2'b00),
    .d({mult0_0_0_23,mult0_0_0_21}),
    .e({mult0_0_0_24,mult0_0_0_22}),
    .fci(\u1/c3 ),
    .f({n2[5],n2[3]}),
    .fco(\u1/c7 ),
    .fx({n2[6],n2[4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1/ucin_al_u336"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1/u43_al_u347  (
    .a({mult0_1_0_31,mult0_1_0_31}),
    .b({open_n1241,mult0_1_0_31}),
    .c(2'b00),
    .d({mult0_1_1_27,mult0_1_1_25}),
    .e({open_n1244,mult0_1_1_26}),
    .fci(\u1/c43 ),
    .f({n2[45],n2[43]}),
    .fx({open_n1260,n2[44]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1/ucin_al_u336"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1/u7_al_u338  (
    .a({mult0_1_0_9,mult0_1_0_7}),
    .b({mult0_1_0_10,mult0_1_0_8}),
    .c(2'b00),
    .d({mult0_0_0_27,mult0_0_0_25}),
    .e({mult0_0_0_28,mult0_0_0_26}),
    .fci(\u1/c7 ),
    .f({n2[9],n2[7]}),
    .fco(\u1/c11 ),
    .fx({n2[10],n2[8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u1/ucin_al_u336"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u1/ucin_al_u336  (
    .a({mult0_1_0_1,1'b0}),
    .b({mult0_1_0_2,mult0_1_0_0}),
    .c(2'b00),
    .d({mult0_0_0_19,1'b1}),
    .e({mult0_0_0_20,mult0_0_0_18}),
    .f({n2[1],open_n1298}),
    .fco(\u1/c3 ),
    .fx({n2[2],n2[0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u15/ucin_al_u348"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u15/u11_al_u351  (
    .a({mult2_0_1_13,mult2_0_1_11}),
    .b({mult2_0_1_14,mult2_0_1_12}),
    .c(2'b00),
    .d({n12[13],n12[11]}),
    .e({n12[14],n12[12]}),
    .fci(\u15/c11 ),
    .fco(\u15/c15 ),
    .fx({n13[14],open_n1319}));
  EG_PHY_LSLICE #(
    //.MACRO("u15/ucin_al_u348"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u15/u15_al_u352  (
    .a({mult2_0_1_17,mult2_0_1_15}),
    .b({mult2_0_1_18,mult2_0_1_16}),
    .c(2'b00),
    .d({n12[17],n12[15]}),
    .e({n12[18],n12[16]}),
    .fci(\u15/c15 ),
    .f({n13[17],n13[15]}),
    .fco(\u15/c19 ),
    .fx({n13[18],n13[16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u15/ucin_al_u348"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u15/u19_al_u353  (
    .a({mult2_0_1_21,mult2_0_1_19}),
    .b({mult2_0_1_22,mult2_0_1_20}),
    .c(2'b00),
    .d({n12[21],n12[19]}),
    .e({n12[22],n12[20]}),
    .fci(\u15/c19 ),
    .f({n13[21],n13[19]}),
    .fco(\u15/c23 ),
    .fx({n13[22],n13[20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u15/ucin_al_u348"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u15/u23_al_u354  (
    .a({mult2_0_1_25,mult2_0_1_23}),
    .b({mult2_0_1_26,mult2_0_1_24}),
    .c(2'b00),
    .d({n12[25],n12[23]}),
    .e({n12[26],n12[24]}),
    .fci(\u15/c23 ),
    .f({n13[25],n13[23]}),
    .fco(\u15/c27 ),
    .fx({n13[26],n13[24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u15/ucin_al_u348"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u15/u27_al_u355  (
    .a({mult2_0_1_29,mult2_0_1_27}),
    .b({mult2_0_1_30,mult2_0_1_28}),
    .c(2'b00),
    .d({n12[29],n12[27]}),
    .e({n12[30],n12[28]}),
    .fci(\u15/c27 ),
    .f({n13[29],n13[27]}),
    .fco(\u15/c31 ),
    .fx({n13[30],n13[28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u15/ucin_al_u348"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u15/u31_al_u356  (
    .a({mult2_0_1_32,mult2_0_1_31}),
    .b({mult2_0_1_32,mult2_0_1_32}),
    .c(2'b00),
    .d({n12[33],n12[31]}),
    .e({n12[34],n12[32]}),
    .fci(\u15/c31 ),
    .f({n13[33],n13[31]}),
    .fco(\u15/c35 ),
    .fx({n13[34],n13[32]}));
  EG_PHY_LSLICE #(
    //.MACRO("u15/ucin_al_u348"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u15/u35_al_u357  (
    .a({mult2_0_1_32,mult2_0_1_32}),
    .b({mult2_0_1_32,mult2_0_1_32}),
    .c(2'b00),
    .d({n12[37],n12[35]}),
    .e({n12[38],n12[36]}),
    .fci(\u15/c35 ),
    .f({n13[37],n13[35]}),
    .fco(\u15/c39 ),
    .fx({n13[38],n13[36]}));
  EG_PHY_LSLICE #(
    //.MACRO("u15/ucin_al_u348"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u15/u39_al_u358  (
    .a({mult2_0_1_32,mult2_0_1_32}),
    .b({mult2_0_1_32,mult2_0_1_32}),
    .c(2'b00),
    .d({n12[41],n12[39]}),
    .e({n12[42],n12[40]}),
    .fci(\u15/c39 ),
    .f({n13[41],n13[39]}),
    .fco(\u15/c43 ),
    .fx({n13[42],n13[40]}));
  EG_PHY_LSLICE #(
    //.MACRO("u15/ucin_al_u348"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u15/u3_al_u349  (
    .a({mult2_0_1_5,mult2_0_1_3}),
    .b({mult2_0_1_6,mult2_0_1_4}),
    .c(2'b00),
    .d({n12[5],n12[3]}),
    .e({n12[6],n12[4]}),
    .fci(\u15/c3 ),
    .fco(\u15/c7 ));
  EG_PHY_LSLICE #(
    //.MACRO("u15/ucin_al_u348"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u15/u43_al_u359  (
    .a({mult2_0_1_32,mult2_0_1_32}),
    .b({open_n1470,mult2_0_1_32}),
    .c(2'b00),
    .d({n12[45],n12[43]}),
    .e({open_n1473,n12[44]}),
    .fci(\u15/c43 ),
    .f({n13[45],n13[43]}),
    .fx({open_n1489,n13[44]}));
  EG_PHY_LSLICE #(
    //.MACRO("u15/ucin_al_u348"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u15/u7_al_u350  (
    .a({mult2_0_1_9,mult2_0_1_7}),
    .b({mult2_0_1_10,mult2_0_1_8}),
    .c(2'b00),
    .d({n12[9],n12[7]}),
    .e({n12[10],n12[8]}),
    .fci(\u15/c7 ),
    .fco(\u15/c11 ));
  EG_PHY_LSLICE #(
    //.MACRO("u15/ucin_al_u348"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u15/ucin_al_u348  (
    .a({mult2_0_1_1,1'b0}),
    .b({mult2_0_1_2,mult2_0_1_0}),
    .c(2'b00),
    .d({n12[1],1'b1}),
    .e({n12[2],n12[0]}),
    .fco(\u15/c3 ));
  EG_PHY_LSLICE #(
    //.MACRO("u5/ucin_al_u360"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u5/u11_al_u363  (
    .a({mult0_0_1_13,mult0_0_1_11}),
    .b({mult0_0_1_14,mult0_0_1_12}),
    .c(2'b00),
    .d({n2[13],n2[11]}),
    .e({n2[14],n2[12]}),
    .fci(\u5/c11 ),
    .f({n7[13],n7[11]}),
    .fco(\u5/c15 ),
    .fx({n7[14],n7[12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u5/ucin_al_u360"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u5/u15_al_u364  (
    .a({mult0_0_1_17,mult0_0_1_15}),
    .b({mult0_0_1_18,mult0_0_1_16}),
    .c(2'b00),
    .d({n2[17],n2[15]}),
    .e({n2[18],n2[16]}),
    .fci(\u5/c15 ),
    .f({n7[17],n7[15]}),
    .fco(\u5/c19 ),
    .fx({n7[18],n7[16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u5/ucin_al_u360"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u5/u19_al_u365  (
    .a({mult0_0_1_21,mult0_0_1_19}),
    .b({mult0_0_1_22,mult0_0_1_20}),
    .c(2'b00),
    .d({n2[21],n2[19]}),
    .e({n2[22],n2[20]}),
    .fci(\u5/c19 ),
    .f({n7[21],n7[19]}),
    .fco(\u5/c23 ),
    .fx({n7[22],n7[20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u5/ucin_al_u360"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u5/u23_al_u366  (
    .a({mult0_0_1_25,mult0_0_1_23}),
    .b({mult0_0_1_26,mult0_0_1_24}),
    .c(2'b00),
    .d({n2[25],n2[23]}),
    .e({n2[26],n2[24]}),
    .fci(\u5/c23 ),
    .f({n7[25],n7[23]}),
    .fco(\u5/c27 ),
    .fx({n7[26],n7[24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u5/ucin_al_u360"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u5/u27_al_u367  (
    .a({mult0_0_1_29,mult0_0_1_27}),
    .b({mult0_0_1_30,mult0_0_1_28}),
    .c(2'b00),
    .d({n2[29],n2[27]}),
    .e({n2[30],n2[28]}),
    .fci(\u5/c27 ),
    .f({n7[29],n7[27]}),
    .fco(\u5/c31 ),
    .fx({n7[30],n7[28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u5/ucin_al_u360"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u5/u31_al_u368  (
    .a({mult0_0_1_31,mult0_0_1_31}),
    .b({mult0_0_1_31,mult0_0_1_31}),
    .c(2'b00),
    .d({n2[33],n2[31]}),
    .e({n2[34],n2[32]}),
    .fci(\u5/c31 ),
    .f({n7[33],n7[31]}),
    .fco(\u5/c35 ),
    .fx({n7[34],n7[32]}));
  EG_PHY_LSLICE #(
    //.MACRO("u5/ucin_al_u360"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u5/u35_al_u369  (
    .a({mult0_0_1_31,mult0_0_1_31}),
    .b({mult0_0_1_31,mult0_0_1_31}),
    .c(2'b00),
    .d({n2[37],n2[35]}),
    .e({n2[38],n2[36]}),
    .fci(\u5/c35 ),
    .f({n7[37],n7[35]}),
    .fco(\u5/c39 ),
    .fx({n7[38],n7[36]}));
  EG_PHY_LSLICE #(
    //.MACRO("u5/ucin_al_u360"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u5/u39_al_u370  (
    .a({mult0_0_1_31,mult0_0_1_31}),
    .b({mult0_0_1_31,mult0_0_1_31}),
    .c(2'b00),
    .d({n2[41],n2[39]}),
    .e({n2[42],n2[40]}),
    .fci(\u5/c39 ),
    .f({n7[41],n7[39]}),
    .fco(\u5/c43 ),
    .fx({n7[42],n7[40]}));
  EG_PHY_LSLICE #(
    //.MACRO("u5/ucin_al_u360"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u5/u3_al_u361  (
    .a({mult0_0_1_5,mult0_0_1_3}),
    .b({mult0_0_1_6,mult0_0_1_4}),
    .c(2'b00),
    .d({n2[5],n2[3]}),
    .e({n2[6],n2[4]}),
    .fci(\u5/c3 ),
    .f({n7[5],n7[3]}),
    .fco(\u5/c7 ),
    .fx({n7[6],n7[4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u5/ucin_al_u360"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u5/u43_al_u371  (
    .a({mult0_0_1_31,mult0_0_1_31}),
    .b({open_n1699,mult0_0_1_31}),
    .c(2'b00),
    .d({n2[45],n2[43]}),
    .e({open_n1702,n2[44]}),
    .fci(\u5/c43 ),
    .f({n7[45],n7[43]}),
    .fx({open_n1718,n7[44]}));
  EG_PHY_LSLICE #(
    //.MACRO("u5/ucin_al_u360"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u5/u7_al_u362  (
    .a({mult0_0_1_9,mult0_0_1_7}),
    .b({mult0_0_1_10,mult0_0_1_8}),
    .c(2'b00),
    .d({n2[9],n2[7]}),
    .e({n2[10],n2[8]}),
    .fci(\u5/c7 ),
    .f({n7[9],n7[7]}),
    .fco(\u5/c11 ),
    .fx({n7[10],n7[8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u5/ucin_al_u360"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u5/ucin_al_u360  (
    .a({mult0_0_1_1,1'b0}),
    .b({mult0_0_1_2,mult0_0_1_0}),
    .c(2'b00),
    .d({n2[1],1'b1}),
    .e({n2[2],n2[0]}),
    .f({n7[1],open_n1756}),
    .fco(\u5/c3 ),
    .fx({n7[2],n7[0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u6/ucin_al_u396"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u6/u11_al_u399  (
    .a({mult1_0_1_13,mult1_0_1_11}),
    .b({mult1_0_1_14,mult1_0_1_12}),
    .c(2'b00),
    .d({mult0_0_0_31,mult0_0_0_29}),
    .e({mult0_0_0_32,mult0_0_0_30}),
    .fci(\u6/c11 ),
    .f({n9[13],n9[11]}),
    .fco(\u6/c15 ),
    .fx({n9[14],n9[12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u6/ucin_al_u396"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u6/u15_al_u400  (
    .a({mult1_0_1_17,mult1_0_1_15}),
    .b({mult1_0_1_18,mult1_0_1_16}),
    .c(2'b00),
    .d({mult0_0_0_35,mult0_0_0_33}),
    .e({mult1_1_1_0,mult0_0_0_34}),
    .fci(\u6/c15 ),
    .f({n9[17],n9[15]}),
    .fco(\u6/c19 ),
    .fx({n9[18],n9[16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u6/ucin_al_u396"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u6/u19_al_u401  (
    .a({mult1_0_1_21,mult1_0_1_19}),
    .b({mult1_0_1_22,mult1_0_1_20}),
    .c(2'b00),
    .d({mult1_1_1_3,mult1_1_1_1}),
    .e({mult1_1_1_4,mult1_1_1_2}),
    .fci(\u6/c19 ),
    .f({n9[21],n9[19]}),
    .fco(\u6/c23 ),
    .fx({n9[22],n9[20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u6/ucin_al_u396"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u6/u23_al_u402  (
    .a({mult1_0_1_25,mult1_0_1_23}),
    .b({mult1_0_1_26,mult1_0_1_24}),
    .c(2'b00),
    .d({mult1_1_1_7,mult1_1_1_5}),
    .e({mult1_1_1_8,mult1_1_1_6}),
    .fci(\u6/c23 ),
    .f({n9[25],n9[23]}),
    .fco(\u6/c27 ),
    .fx({n9[26],n9[24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u6/ucin_al_u396"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u6/u27_al_u403  (
    .a({mult1_0_1_29,mult1_0_1_27}),
    .b({mult1_0_1_30,mult1_0_1_28}),
    .c(2'b00),
    .d({mult1_1_1_11,mult1_1_1_9}),
    .e({mult1_1_1_12,mult1_1_1_10}),
    .fci(\u6/c27 ),
    .f({n9[29],n9[27]}),
    .fco(\u6/c31 ),
    .fx({n9[30],n9[28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u6/ucin_al_u396"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u6/u31_al_u404  (
    .a({open_n1849,mult1_0_1_31}),
    .c(2'b00),
    .d({open_n1854,mult1_1_1_13}),
    .fci(\u6/c31 ),
    .f({open_n1871,n9[31]}),
    .fx({open_n1873,n9[32]}));
  EG_PHY_LSLICE #(
    //.MACRO("u6/ucin_al_u396"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u6/u3_al_u397  (
    .a({mult1_0_1_5,mult1_0_1_3}),
    .b({mult1_0_1_6,mult1_0_1_4}),
    .c(2'b00),
    .d({mult0_0_0_23,mult0_0_0_21}),
    .e({mult0_0_0_24,mult0_0_0_22}),
    .fci(\u6/c3 ),
    .f({n9[5],n9[3]}),
    .fco(\u6/c7 ),
    .fx({n9[6],n9[4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u6/ucin_al_u396"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u6/u7_al_u398  (
    .a({mult1_0_1_9,mult1_0_1_7}),
    .b({mult1_0_1_10,mult1_0_1_8}),
    .c(2'b00),
    .d({mult0_0_0_27,mult0_0_0_25}),
    .e({mult0_0_0_28,mult0_0_0_26}),
    .fci(\u6/c7 ),
    .f({n9[9],n9[7]}),
    .fco(\u6/c11 ),
    .fx({n9[10],n9[8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u6/ucin_al_u396"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u6/ucin_al_u396  (
    .a({mult1_0_1_1,1'b0}),
    .b({mult1_0_1_2,mult1_0_1_0}),
    .c(2'b00),
    .d({mult0_0_0_19,1'b1}),
    .e({mult0_0_0_20,mult0_0_0_18}),
    .f({n9[1],open_n1929}),
    .fco(\u6/c3 ),
    .fx({n9[2],n9[0]}));
  EG_PHY_LSLICE #(
    //.MACRO("u7/ucin_al_u372"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u7/u11_al_u375  (
    .a({mult1_1_0_13,mult1_1_0_11}),
    .b({mult1_1_0_14,mult1_1_0_12}),
    .c(2'b00),
    .d({n9[13],n9[11]}),
    .e({n9[14],n9[12]}),
    .fci(\u7/c11 ),
    .fco(\u7/c15 ),
    .fx({n11[14],open_n1950}));
  EG_PHY_LSLICE #(
    //.MACRO("u7/ucin_al_u372"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u7/u15_al_u376  (
    .a({mult1_1_0_17,mult1_1_0_15}),
    .b({mult1_1_0_18,mult1_1_0_16}),
    .c(2'b00),
    .d({n9[17],n9[15]}),
    .e({n9[18],n9[16]}),
    .fci(\u7/c15 ),
    .f({n11[17],n11[15]}),
    .fco(\u7/c19 ),
    .fx({n11[18],n11[16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u7/ucin_al_u372"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u7/u19_al_u377  (
    .a({mult1_1_0_21,mult1_1_0_19}),
    .b({mult1_1_0_22,mult1_1_0_20}),
    .c(2'b00),
    .d({n9[21],n9[19]}),
    .e({n9[22],n9[20]}),
    .fci(\u7/c19 ),
    .f({n11[21],n11[19]}),
    .fco(\u7/c23 ),
    .fx({n11[22],n11[20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u7/ucin_al_u372"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u7/u23_al_u378  (
    .a({mult1_1_0_25,mult1_1_0_23}),
    .b({mult1_1_0_26,mult1_1_0_24}),
    .c(2'b00),
    .d({n9[25],n9[23]}),
    .e({n9[26],n9[24]}),
    .fci(\u7/c23 ),
    .f({n11[25],n11[23]}),
    .fco(\u7/c27 ),
    .fx({n11[26],n11[24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u7/ucin_al_u372"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u7/u27_al_u379  (
    .a({mult1_1_0_29,mult1_1_0_27}),
    .b({mult1_1_0_30,mult1_1_0_28}),
    .c(2'b00),
    .d({n9[29],n9[27]}),
    .e({n9[30],n9[28]}),
    .fci(\u7/c27 ),
    .f({n11[29],n11[27]}),
    .fco(\u7/c31 ),
    .fx({n11[30],n11[28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u7/ucin_al_u372"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u7/u31_al_u380  (
    .a({1'b0,mult1_1_0_31}),
    .b({1'b0,mult1_1_1_14}),
    .c(2'b00),
    .d({mult1_1_1_15,n9[31]}),
    .e({mult1_1_1_16,n9[32]}),
    .fci(\u7/c31 ),
    .f({n11[33],n11[31]}),
    .fco(\u7/c35 ),
    .fx({n11[34],n11[32]}));
  EG_PHY_LSLICE #(
    //.MACRO("u7/ucin_al_u372"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u7/u35_al_u381  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b00),
    .d({mult1_1_1_19,mult1_1_1_17}),
    .e({mult1_1_1_20,mult1_1_1_18}),
    .fci(\u7/c35 ),
    .f({n11[37],n11[35]}),
    .fco(\u7/c39 ),
    .fx({n11[38],n11[36]}));
  EG_PHY_LSLICE #(
    //.MACRO("u7/ucin_al_u372"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u7/u39_al_u382  (
    .a(2'b00),
    .b(2'b00),
    .c(2'b00),
    .d({mult1_1_1_23,mult1_1_1_21}),
    .e({mult1_1_1_24,mult1_1_1_22}),
    .fci(\u7/c39 ),
    .f({n11[41],n11[39]}),
    .fco(\u7/c43 ),
    .fx({n11[42],n11[40]}));
  EG_PHY_LSLICE #(
    //.MACRO("u7/ucin_al_u372"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u7/u3_al_u373  (
    .a({mult1_1_0_5,mult1_1_0_3}),
    .b({mult1_1_0_6,mult1_1_0_4}),
    .c(2'b00),
    .d({n9[5],n9[3]}),
    .e({n9[6],n9[4]}),
    .fci(\u7/c3 ),
    .fco(\u7/c7 ));
  EG_PHY_LSLICE #(
    //.MACRO("u7/ucin_al_u372"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u7/u43_al_u383  (
    .a(2'b00),
    .b({open_n2101,1'b0}),
    .c(2'b00),
    .d({mult1_1_1_27,mult1_1_1_25}),
    .e({open_n2104,mult1_1_1_26}),
    .fci(\u7/c43 ),
    .f({n11[45],n11[43]}),
    .fx({open_n2120,n11[44]}));
  EG_PHY_LSLICE #(
    //.MACRO("u7/ucin_al_u372"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u7/u7_al_u374  (
    .a({mult1_1_0_9,mult1_1_0_7}),
    .b({mult1_1_0_10,mult1_1_0_8}),
    .c(2'b00),
    .d({n9[9],n9[7]}),
    .e({n9[10],n9[8]}),
    .fci(\u7/c7 ),
    .fco(\u7/c11 ));
  EG_PHY_LSLICE #(
    //.MACRO("u7/ucin_al_u372"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u7/ucin_al_u372  (
    .a({mult1_1_0_1,1'b0}),
    .b({mult1_1_0_2,mult1_1_0_0}),
    .c(2'b00),
    .d({n9[1],1'b1}),
    .e({n9[2],n9[0]}),
    .fco(\u7/c3 ));
  EG_PHY_LSLICE #(
    //.MACRO("u8/ucin_al_u384"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u8/u11_al_u387  (
    .a({mult0_1_0_13,mult0_1_0_11}),
    .b({mult0_1_0_14,mult0_1_0_12}),
    .c(2'b00),
    .d({mult0_0_0_31,mult0_0_0_29}),
    .e({mult0_0_0_32,mult0_0_0_30}),
    .fci(\u8/c11 ),
    .f({n12[13],n12[11]}),
    .fco(\u8/c15 ),
    .fx({n12[14],n12[12]}));
  EG_PHY_LSLICE #(
    //.MACRO("u8/ucin_al_u384"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u8/u15_al_u388  (
    .a({mult0_1_0_17,mult0_1_0_15}),
    .b({mult0_1_0_18,mult0_1_0_16}),
    .c(2'b00),
    .d({mult0_0_0_35,mult0_0_0_33}),
    .e({mult2_1_1_0,mult0_0_0_34}),
    .fci(\u8/c15 ),
    .f({n12[17],n12[15]}),
    .fco(\u8/c19 ),
    .fx({n12[18],n12[16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u8/ucin_al_u384"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u8/u19_al_u389  (
    .a({mult0_1_0_21,mult0_1_0_19}),
    .b({mult0_1_0_22,mult0_1_0_20}),
    .c(2'b00),
    .d({mult2_1_1_3,mult2_1_1_1}),
    .e({mult2_1_1_4,mult2_1_1_2}),
    .fci(\u8/c19 ),
    .f({n12[21],n12[19]}),
    .fco(\u8/c23 ),
    .fx({n12[22],n12[20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u8/ucin_al_u384"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u8/u23_al_u390  (
    .a({mult0_1_0_25,mult0_1_0_23}),
    .b({mult0_1_0_26,mult0_1_0_24}),
    .c(2'b00),
    .d({mult2_1_1_7,mult2_1_1_5}),
    .e({mult2_1_1_8,mult2_1_1_6}),
    .fci(\u8/c23 ),
    .f({n12[25],n12[23]}),
    .fco(\u8/c27 ),
    .fx({n12[26],n12[24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u8/ucin_al_u384"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u8/u27_al_u391  (
    .a({mult0_1_0_29,mult0_1_0_27}),
    .b({mult0_1_0_30,mult0_1_0_28}),
    .c(2'b00),
    .d({mult2_1_1_11,mult2_1_1_9}),
    .e({mult2_1_1_12,mult2_1_1_10}),
    .fci(\u8/c27 ),
    .f({n12[29],n12[27]}),
    .fco(\u8/c31 ),
    .fx({n12[30],n12[28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u8/ucin_al_u384"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u8/u31_al_u392  (
    .a({mult0_1_0_31,mult0_1_0_31}),
    .b({mult0_1_0_31,mult0_1_0_31}),
    .c(2'b00),
    .d({mult2_1_1_15,mult2_1_1_13}),
    .e({mult2_1_1_16,mult2_1_1_14}),
    .fci(\u8/c31 ),
    .f({n12[33],n12[31]}),
    .fco(\u8/c35 ),
    .fx({n12[34],n12[32]}));
  EG_PHY_LSLICE #(
    //.MACRO("u8/ucin_al_u384"),
    //.R_POSITION("X0Y4Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u8/u35_al_u393  (
    .a({mult0_1_0_31,mult0_1_0_31}),
    .b({mult0_1_0_31,mult0_1_0_31}),
    .c(2'b00),
    .d({mult2_1_1_19,mult2_1_1_17}),
    .e({mult2_1_1_20,mult2_1_1_18}),
    .fci(\u8/c35 ),
    .f({n12[37],n12[35]}),
    .fco(\u8/c39 ),
    .fx({n12[38],n12[36]}));
  EG_PHY_LSLICE #(
    //.MACRO("u8/ucin_al_u384"),
    //.R_POSITION("X0Y5Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u8/u39_al_u394  (
    .a({mult0_1_0_31,mult0_1_0_31}),
    .b({mult0_1_0_31,mult0_1_0_31}),
    .c(2'b00),
    .d({mult2_1_1_23,mult2_1_1_21}),
    .e({mult2_1_1_24,mult2_1_1_22}),
    .fci(\u8/c39 ),
    .f({n12[41],n12[39]}),
    .fco(\u8/c43 ),
    .fx({n12[42],n12[40]}));
  EG_PHY_LSLICE #(
    //.MACRO("u8/ucin_al_u384"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u8/u3_al_u385  (
    .a({mult0_1_0_5,mult0_1_0_3}),
    .b({mult0_1_0_6,mult0_1_0_4}),
    .c(2'b00),
    .d({mult0_0_0_23,mult0_0_0_21}),
    .e({mult0_0_0_24,mult0_0_0_22}),
    .fci(\u8/c3 ),
    .f({n12[5],n12[3]}),
    .fco(\u8/c7 ),
    .fx({n12[6],n12[4]}));
  EG_PHY_LSLICE #(
    //.MACRO("u8/ucin_al_u384"),
    //.R_POSITION("X0Y5Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u8/u43_al_u395  (
    .a({mult0_1_0_31,mult0_1_0_31}),
    .b({open_n2330,mult0_1_0_31}),
    .c(2'b00),
    .d({mult2_1_1_27,mult2_1_1_25}),
    .e({open_n2333,mult2_1_1_26}),
    .fci(\u8/c43 ),
    .f({n12[45],n12[43]}),
    .fx({open_n2349,n12[44]}));
  EG_PHY_LSLICE #(
    //.MACRO("u8/ucin_al_u384"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u8/u7_al_u386  (
    .a({mult0_1_0_9,mult0_1_0_7}),
    .b({mult0_1_0_10,mult0_1_0_8}),
    .c(2'b00),
    .d({mult0_0_0_27,mult0_0_0_25}),
    .e({mult0_0_0_28,mult0_0_0_26}),
    .fci(\u8/c7 ),
    .f({n12[9],n12[7]}),
    .fco(\u8/c11 ),
    .fx({n12[10],n12[8]}));
  EG_PHY_LSLICE #(
    //.MACRO("u8/ucin_al_u384"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u8/ucin_al_u384  (
    .a({mult0_1_0_1,1'b0}),
    .b({mult0_1_0_2,mult0_1_0_0}),
    .c(2'b00),
    .d({mult0_0_0_19,1'b1}),
    .e({mult0_0_0_20,mult0_0_0_18}),
    .f({n12[1],open_n2387}),
    .fco(\u8/c3 ),
    .fx({n12[2],n12[0]}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F8880  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [8]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [9]));  // al_ip/div_signed_gate.v(4358)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F8990  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [14]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [15]));  // al_ip/div_signed_gate.v(4142)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F8AA0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [19]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [20]));  // al_ip/div_signed_gate.v(4196)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F8CC0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [20]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [21]));  // al_ip/div_signed_gate.v(4205)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F8DD0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [22]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [23]));  // al_ip/div_signed_gate.v(4223)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F8FF0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [18]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [19]));  // al_ip/div_signed_gate.v(4178)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256A66F9210  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [0]),
    .sr(i_rstn),
    .q(div_signed_quo[0]));  // al_ip/div_signed_gate.v(4367)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F9430  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [11]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [12]));  // al_ip/div_signed_gate.v(4115)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F9540  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [23]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [24]));  // al_ip/div_signed_gate.v(4232)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F9650  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [15]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [16]));  // al_ip/div_signed_gate.v(4151)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F9760  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [24]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [25]));  // al_ip/div_signed_gate.v(4241)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66F9BA0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [26]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [26]));  // al_ip/div_signed_gate.v(3962)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256A66F9CB0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [1]),
    .sr(i_rstn),
    .q(div_signed_quo[1]));  // al_ip/div_signed_gate.v(4376)
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y16Z0"),
    .ALUTYPE("A_LE_B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F9DC0_al_u424  (
    .a({open_n2402,1'b0}),
    .b({open_n2403,1'b1}),
    .clk(i_clk),
    .fci(\u_DIV_SIGNED/al_00000256AA88D630 ),
    .sr(div_signed_start),
    .f({open_n2420,\u_DIV_SIGNED/al_00000256AA3DB7F0 }),
    .q({open_n2424,\u_DIV_SIGNED/al_00000256AA0CEB40 [0]}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F9ED0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [0]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [1]));  // al_ip/div_signed_gate.v(4088)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66F9FE0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [3]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [4]));  // al_ip/div_signed_gate.v(4313)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FA0F0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [4]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [5]));  // al_ip/div_signed_gate.v(4322)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FA200  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [6]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [7]));  // al_ip/div_signed_gate.v(4340)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256A66FA310  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [2]),
    .sr(i_rstn),
    .q(div_signed_quo[2]));  // al_ip/div_signed_gate.v(4475)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FA420  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [25]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [25]));  // al_ip/div_signed_gate.v(3953)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FA530  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [10]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [11]));  // al_ip/div_signed_gate.v(4106)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FA640  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [12]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [13]));  // al_ip/div_signed_gate.v(4124)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FA860  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [2]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [3]));  // al_ip/div_signed_gate.v(4286)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FAB90  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [27]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [27]));  // al_ip/div_signed_gate.v(3971)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FACA0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [5]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [6]));  // al_ip/div_signed_gate.v(4331)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FAFD0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [28]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [28]));  // al_ip/div_signed_gate.v(3980)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FB1F0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [9]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [10]));  // al_ip/div_signed_gate.v(4097)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FB300  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [13]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [14]));  // al_ip/div_signed_gate.v(4133)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FB410  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [16]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [17]));  // al_ip/div_signed_gate.v(4160)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FB630  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [17]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [18]));  // al_ip/div_signed_gate.v(4169)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FB740  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [21]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [22]));  // al_ip/div_signed_gate.v(4214)
  EG_PHY_LSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256A66FB850_al_u414"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h0005),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256A66FB850_al_u414  (
    .a({\u_DIV_SIGNED/al_00000256AA0CF470 [1],1'b0}),
    .b({\u_DIV_SIGNED/al_00000256AA0CF470 [2],\u_DIV_SIGNED/al_00000256AA0CF470 [0]}),
    .c(2'b11),
    .d({\u_DIV_SIGNED/al_00000256AA0D0BA0 [1],1'b1}),
    .e({\u_DIV_SIGNED/al_00000256AA0D0BA0 [2],\u_DIV_SIGNED/al_00000256AA0D0BA0 [0]}),
    .f({\u_DIV_SIGNED/al_00000256AA400D60 [1],open_n2461}),
    .fco(\u_DIV_SIGNED/al_00000256AA898FD0 ),
    .fx({\u_DIV_SIGNED/al_00000256AA400D60 [2],\u_DIV_SIGNED/al_00000256AA400D60 [0]}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FBA70  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [31]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [31]));  // al_ip/div_signed_gate.v(4016)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FC2F0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [23]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [23]));  // al_ip/div_signed_gate.v(3935)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FC400  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [30]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [30]));  // al_ip/div_signed_gate.v(4007)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FC620  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [29]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [29]));  // al_ip/div_signed_gate.v(3989)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FC840  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [24]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [24]));  // al_ip/div_signed_gate.v(3944)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FCA60  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [1]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [2]));  // al_ip/div_signed_gate.v(4187)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256A66FCB70  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [7]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [8]));  // al_ip/div_signed_gate.v(4349)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FE0B0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [15]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [15]));  // al_ip/div_signed_gate.v(3854)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FE3E0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [16]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [16]));  // al_ip/div_signed_gate.v(3863)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FE820  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [17]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [17]));  // al_ip/div_signed_gate.v(3872)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FEE80  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [18]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [18]));  // al_ip/div_signed_gate.v(3881)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FEF90  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [19]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [19]));  // al_ip/div_signed_gate.v(3890)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FF1B0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [20]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [20]));  // al_ip/div_signed_gate.v(3908)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FF700  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [21]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [21]));  // al_ip/div_signed_gate.v(3917)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FF810  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [22]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [22]));  // al_ip/div_signed_gate.v(3926)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FFB40  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [13]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [13]));  // al_ip/div_signed_gate.v(3836)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256A66FFD60  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [14]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [14]));  // al_ip/div_signed_gate.v(3845)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA39D160  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [25]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [26]));  // al_ip/div_signed_gate.v(4250)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A1780  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [26]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [27]));  // al_ip/div_signed_gate.v(4259)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A1AB0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [11]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [10]));  // al_ip/div_signed_gate.v(3242)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A1CD0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [12]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [11]));  // al_ip/div_signed_gate.v(3251)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A2110  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [17]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [16]));  // al_ip/div_signed_gate.v(3296)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A2550  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [1]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [0]));  // al_ip/div_signed_gate.v(3224)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A2990  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [14]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [13]));  // al_ip/div_signed_gate.v(3269)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A2AA0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [13]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [12]));  // al_ip/div_signed_gate.v(3260)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A2BB0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [18]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [17]));  // al_ip/div_signed_gate.v(3305)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A2CC0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [20]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [19]));  // al_ip/div_signed_gate.v(3323)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A2EE0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [3]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [2]));  // al_ip/div_signed_gate.v(3332)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A3100  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [21]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [20]));  // al_ip/div_signed_gate.v(3341)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A3210  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [4]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [3]));  // al_ip/div_signed_gate.v(3431)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A3320  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [8]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [7]));  // al_ip/div_signed_gate.v(3764)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A3540  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [15]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [14]));  // al_ip/div_signed_gate.v(3278)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A3650  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [22]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [21]));  // al_ip/div_signed_gate.v(3350)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A3760  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [23]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [22]));  // al_ip/div_signed_gate.v(3359)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A3870  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [25]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [24]));  // al_ip/div_signed_gate.v(3377)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A3980  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [9]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [8]));  // al_ip/div_signed_gate.v(3773)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A3ED0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [19]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [18]));  // al_ip/div_signed_gate.v(3314)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A3FE0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [26]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [25]));  // al_ip/div_signed_gate.v(3386)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A40F0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [27]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [26]));  // al_ip/div_signed_gate.v(3395)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A4200  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [28]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [27]));  // al_ip/div_signed_gate.v(3404)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A4310  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [29]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [28]));  // al_ip/div_signed_gate.v(3413)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A4420  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [6]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [5]));  // al_ip/div_signed_gate.v(3629)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A4530  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [30]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [29]));  // al_ip/div_signed_gate.v(3422)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A4640  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [31]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [30]));  // al_ip/div_signed_gate.v(3440)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A4750  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [31]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [31]));  // al_ip/div_signed_gate.v(3449)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A4860  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [7]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [6]));  // al_ip/div_signed_gate.v(3728)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A4970  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [16]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [15]));  // al_ip/div_signed_gate.v(3287)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A4A80  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [24]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [23]));  // al_ip/div_signed_gate.v(3368)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A4CA0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [32]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [32]));  // al_ip/div_signed_gate.v(3458)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A4DB0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [33]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [33]));  // al_ip/div_signed_gate.v(3467)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A50E0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [2]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [1]));  // al_ip/div_signed_gate.v(3233)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A5520  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [10]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [9]));  // al_ip/div_signed_gate.v(3782)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A5850  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D0BA0 [5]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [4]));  // al_ip/div_signed_gate.v(3530)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A5C90  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [29]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [30]));  // al_ip/div_signed_gate.v(4295)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A5DA0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [30]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [31]));  // al_ip/div_signed_gate.v(4304)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A5FC0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [3]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [3]));  // al_ip/div_signed_gate.v(3998)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A60D0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [7]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [7]));  // al_ip/div_signed_gate.v(4052)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A61E0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [39]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [39]));  // al_ip/div_signed_gate.v(3521)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A62F0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [61]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [61]));  // al_ip/div_signed_gate.v(3746)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A6510  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [10]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [10]));  // al_ip/div_signed_gate.v(3809)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A6620  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [11]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [11]));  // al_ip/div_signed_gate.v(3818)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A6730  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [55]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [55]));  // al_ip/div_signed_gate.v(3683)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A6840  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [56]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [56]));  // al_ip/div_signed_gate.v(3692)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A6950  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [43]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [43]));  // al_ip/div_signed_gate.v(3566)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A6A60  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [5]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [5]));  // al_ip/div_signed_gate.v(4034)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A6B70  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [8]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [8]));  // al_ip/div_signed_gate.v(4061)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A6C80  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [46]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [46]));  // al_ip/div_signed_gate.v(3593)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A6D90  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [12]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [12]));  // al_ip/div_signed_gate.v(3827)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A6EA0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [42]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [42]));  // al_ip/div_signed_gate.v(3557)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A6FB0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [41]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [41]));  // al_ip/div_signed_gate.v(3548)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A70C0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [60]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [60]));  // al_ip/div_signed_gate.v(3737)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A71D0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [48]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [48]));  // al_ip/div_signed_gate.v(3611)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A72E0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [36]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [36]));  // al_ip/div_signed_gate.v(3494)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A73F0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [47]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [47]));  // al_ip/div_signed_gate.v(3602)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A7500  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [54]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [54]));  // al_ip/div_signed_gate.v(3674)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA3A7610  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D7970 [62]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [62]));  // al_ip/div_signed_gate.v(3755)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A7720  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [27]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [28]));  // al_ip/div_signed_gate.v(4268)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A7830  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [0]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [0]));  // al_ip/div_signed_gate.v(3791)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A7940  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [38]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [38]));  // al_ip/div_signed_gate.v(3512)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A7A50  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [57]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [57]));  // al_ip/div_signed_gate.v(3701)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A7B60  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [1]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [1]));  // al_ip/div_signed_gate.v(3800)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A7C70  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [45]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [45]));  // al_ip/div_signed_gate.v(3584)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A7D80  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [40]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [40]));  // al_ip/div_signed_gate.v(3539)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A7E90  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [50]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [50]));  // al_ip/div_signed_gate.v(3638)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A7FA0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [59]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [59]));  // al_ip/div_signed_gate.v(3719)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A80B0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [4]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [4]));  // al_ip/div_signed_gate.v(4025)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A81C0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [34]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [34]));  // al_ip/div_signed_gate.v(3476)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A82D0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [2]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [2]));  // al_ip/div_signed_gate.v(3899)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A83E0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [6]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [6]));  // al_ip/div_signed_gate.v(4043)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A84F0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA402C70 [9]),
    .q(\u_DIV_SIGNED/al_00000256AA0CF470 [9]));  // al_ip/div_signed_gate.v(4070)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A8600  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [49]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [49]));  // al_ip/div_signed_gate.v(3620)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A8710  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [58]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [58]));  // al_ip/div_signed_gate.v(3710)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A8820  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [51]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [51]));  // al_ip/div_signed_gate.v(3647)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A8930  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [37]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [37]));  // al_ip/div_signed_gate.v(3503)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A8A40  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [52]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [52]));  // al_ip/div_signed_gate.v(3656)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_SIGNED/al_00000256AA3A8B50  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0CEB40 [28]),
    .sr(div_signed_start),
    .q(\u_DIV_SIGNED/al_00000256AA0CEB40 [29]));  // al_ip/div_signed_gate.v(4277)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A8C60  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [44]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [44]));  // al_ip/div_signed_gate.v(3575)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A8D70  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [35]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [35]));  // al_ip/div_signed_gate.v(3485)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA3A8E80  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D80E0 [53]),
    .q(\u_DIV_SIGNED/al_00000256AA0D0BA0 [53]));  // al_ip/div_signed_gate.v(3665)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47F090  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [0]),
    .sr(i_rstn),
    .q(div_signed_rem[0]));  // al_ip/div_signed_gate.v(4655)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47F1A0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [3]),
    .sr(i_rstn),
    .q(div_signed_rem[3]));  // al_ip/div_signed_gate.v(4862)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47F2B0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [9]),
    .sr(i_rstn),
    .q(div_signed_quo[9]));  // al_ip/div_signed_gate.v(4646)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47F3C0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [17]),
    .sr(i_rstn),
    .q(div_signed_rem[17]));  // al_ip/div_signed_gate.v(4736)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47F4D0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [19]),
    .sr(i_rstn),
    .q(div_signed_rem[19]));  // al_ip/div_signed_gate.v(4754)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47F5E0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [6]),
    .sr(i_rstn),
    .q(div_signed_quo[6]));  // al_ip/div_signed_gate.v(4619)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47F6F0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D38B0 [1]),
    .sr(i_rstn),
    .q(\u_DIV_SIGNED/al_00000256AA0CE7C0 [1]));  // al_ip/div_signed_gate.v(4952)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47F800  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [13]),
    .sr(i_rstn),
    .q(div_signed_quo[13]));  // al_ip/div_signed_gate.v(4412)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47F910  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [6]),
    .sr(i_rstn),
    .q(div_signed_rem[6]));  // al_ip/div_signed_gate.v(4907)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47FA20  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [26]),
    .sr(i_rstn),
    .q(div_signed_rem[26]));  // al_ip/div_signed_gate.v(4826)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47FB30  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [27]),
    .sr(i_rstn),
    .q(div_signed_quo[27]));  // al_ip/div_signed_gate.v(4547)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47FC40  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [30]),
    .sr(i_rstn),
    .q(div_signed_quo[30]));  // al_ip/div_signed_gate.v(4583)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47FD50  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [11]),
    .sr(i_rstn),
    .q(div_signed_rem[11]));  // al_ip/div_signed_gate.v(4682)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47FE60  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [12]),
    .sr(i_rstn),
    .q(div_signed_rem[12]));  // al_ip/div_signed_gate.v(4691)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA47FF70  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [20]),
    .sr(i_rstn),
    .q(div_signed_rem[20]));  // al_ip/div_signed_gate.v(4772)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA480080  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [5]),
    .sr(i_rstn),
    .q(div_signed_quo[5]));  // al_ip/div_signed_gate.v(4610)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA480190  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [14]),
    .sr(i_rstn),
    .q(div_signed_quo[14]));  // al_ip/div_signed_gate.v(4421)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4802A0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [7]),
    .sr(i_rstn),
    .q(div_signed_rem[7]));  // al_ip/div_signed_gate.v(4916)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4803B0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [10]),
    .sr(i_rstn),
    .q(div_signed_rem[10]));  // al_ip/div_signed_gate.v(4673)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4804C0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [23]),
    .sr(i_rstn),
    .q(div_signed_rem[23]));  // al_ip/div_signed_gate.v(4799)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4805D0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [26]),
    .sr(i_rstn),
    .q(div_signed_quo[26]));  // al_ip/div_signed_gate.v(4538)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4806E0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [3]),
    .sr(i_rstn),
    .q(div_signed_quo[3]));  // al_ip/div_signed_gate.v(4574)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4807F0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [29]),
    .sr(i_rstn),
    .q(div_signed_quo[29]));  // al_ip/div_signed_gate.v(4565)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA480900  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [28]),
    .sr(i_rstn),
    .q(div_signed_quo[28]));  // al_ip/div_signed_gate.v(4556)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA480A10  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D38B0 [2]),
    .sr(i_rstn),
    .q(\u_DIV_SIGNED/al_00000256AA0CE7C0 [2]));  // al_ip/div_signed_gate.v(4961)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA480B20  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [14]),
    .sr(i_rstn),
    .q(div_signed_rem[14]));  // al_ip/div_signed_gate.v(4709)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA480C30  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [13]),
    .sr(i_rstn),
    .q(div_signed_rem[13]));  // al_ip/div_signed_gate.v(4700)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA480D40  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [16]),
    .sr(i_rstn),
    .q(div_signed_rem[16]));  // al_ip/div_signed_gate.v(4727)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA480E50  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [8]),
    .sr(i_rstn),
    .q(div_signed_rem[8]));  // al_ip/div_signed_gate.v(4925)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA480F60  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [21]),
    .sr(i_rstn),
    .q(div_signed_rem[21]));  // al_ip/div_signed_gate.v(4781)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA481070  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [24]),
    .sr(i_rstn),
    .q(div_signed_quo[24]));  // al_ip/div_signed_gate.v(4520)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA481180  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [11]),
    .sr(i_rstn),
    .q(div_signed_quo[11]));  // al_ip/div_signed_gate.v(4394)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA481290  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D38B0 [3]),
    .sr(i_rstn),
    .q(\u_DIV_SIGNED/al_00000256AA0CE7C0 [3]));  // al_ip/div_signed_gate.v(4970)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4813A0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [5]),
    .sr(i_rstn),
    .q(div_signed_rem[5]));  // al_ip/div_signed_gate.v(4898)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4814B0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [9]),
    .sr(i_rstn),
    .q(div_signed_rem[9]));  // al_ip/div_signed_gate.v(4934)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4815C0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [18]),
    .sr(i_rstn),
    .q(div_signed_rem[18]));  // al_ip/div_signed_gate.v(4745)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4816D0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [7]),
    .sr(i_rstn),
    .q(div_signed_quo[7]));  // al_ip/div_signed_gate.v(4628)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4817E0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D38B0 [4]),
    .sr(i_rstn),
    .q(\u_DIV_SIGNED/al_00000256AA0CE7C0 [4]));  // al_ip/div_signed_gate.v(4979)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4818F0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [22]),
    .sr(i_rstn),
    .q(div_signed_rem[22]));  // al_ip/div_signed_gate.v(4790)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA481A00  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D38B0 [5]),
    .sr(i_rstn),
    .q(\u_DIV_SIGNED/al_00000256AA0CE7C0 [5]));  // al_ip/div_signed_gate.v(4988)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA481B10  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [4]),
    .sr(i_rstn),
    .q(div_signed_quo[4]));  // al_ip/div_signed_gate.v(4601)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA481C20  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [15]),
    .sr(i_rstn),
    .q(div_signed_rem[15]));  // al_ip/div_signed_gate.v(4718)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA481D30  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [8]),
    .sr(i_rstn),
    .q(div_signed_quo[8]));  // al_ip/div_signed_gate.v(4637)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA481E40  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [17]),
    .sr(i_rstn),
    .q(div_signed_quo[17]));  // al_ip/div_signed_gate.v(4448)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA481F50  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [20]),
    .sr(i_rstn),
    .q(div_signed_quo[20]));  // al_ip/div_signed_gate.v(4484)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA482060  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [16]),
    .sr(i_rstn),
    .q(div_signed_quo[16]));  // al_ip/div_signed_gate.v(4439)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA482170  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [23]),
    .sr(i_rstn),
    .q(div_signed_quo[23]));  // al_ip/div_signed_gate.v(4511)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA482390  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [12]),
    .sr(i_rstn),
    .q(div_signed_quo[12]));  // al_ip/div_signed_gate.v(4403)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4824A0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [15]),
    .sr(i_rstn),
    .q(div_signed_quo[15]));  // al_ip/div_signed_gate.v(4430)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4825B0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [4]),
    .sr(i_rstn),
    .q(div_signed_rem[4]));  // al_ip/div_signed_gate.v(4889)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4826C0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [24]),
    .sr(i_rstn),
    .q(div_signed_rem[24]));  // al_ip/div_signed_gate.v(4808)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4827D0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [31]),
    .sr(i_rstn),
    .q(div_signed_quo[31]));  // al_ip/div_signed_gate.v(4592)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4828E0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [25]),
    .sr(i_rstn),
    .q(div_signed_rem[25]));  // al_ip/div_signed_gate.v(4817)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA4829F0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [27]),
    .sr(i_rstn),
    .q(div_signed_rem[27]));  // al_ip/div_signed_gate.v(4835)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA482B00  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [18]),
    .sr(i_rstn),
    .q(div_signed_quo[18]));  // al_ip/div_signed_gate.v(4457)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA482C10  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [21]),
    .sr(i_rstn),
    .q(div_signed_quo[21]));  // al_ip/div_signed_gate.v(4493)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA482D20  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [22]),
    .sr(i_rstn),
    .q(div_signed_quo[22]));  // al_ip/div_signed_gate.v(4502)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA482E30  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [25]),
    .sr(i_rstn),
    .q(div_signed_quo[25]));  // al_ip/div_signed_gate.v(4529)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA482F40  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA0D38B0 [0]),
    .sr(i_rstn),
    .q(\u_DIV_SIGNED/al_00000256AA0CE7C0 [0]));  // al_ip/div_signed_gate.v(4943)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA483050  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [19]),
    .sr(i_rstn),
    .q(div_signed_quo[19]));  // al_ip/div_signed_gate.v(4466)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA483160  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [1]),
    .sr(i_rstn),
    .q(div_signed_rem[1]));  // al_ip/div_signed_gate.v(4664)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA483270  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [2]),
    .sr(i_rstn),
    .q(div_signed_rem[2]));  // al_ip/div_signed_gate.v(4763)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA483380  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4073C0 [10]),
    .sr(i_rstn),
    .q(div_signed_quo[10]));  // al_ip/div_signed_gate.v(4385)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA483AF0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [30]),
    .sr(i_rstn),
    .q(div_signed_rem[30]));  // al_ip/div_signed_gate.v(4871)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA484150  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [28]),
    .sr(i_rstn),
    .q(div_signed_rem[28]));  // al_ip/div_signed_gate.v(4844)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA485BE0  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [29]),
    .sr(i_rstn),
    .q(div_signed_rem[29]));  // al_ip/div_signed_gate.v(4853)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA486570  (
    .ce(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA4098F0 [31]),
    .sr(i_rstn),
    .q(div_signed_rem[31]));  // al_ip/div_signed_gate.v(4880)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_SIGNED/al_00000256AA4D31A0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .b(\u_DIV_SIGNED/al_00000256AA8940C0 ),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D29D0 [2]),
    .o(\u_DIV_SIGNED/al_00000256AA0D38B0 [2]));  // al_ip/div_signed_gate.v(975)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_SIGNED/al_00000256AA4D4A10  (
    .a(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .b(\u_DIV_SIGNED/al_00000256AA8940C0 ),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D29D0 [5]),
    .o(\u_DIV_SIGNED/al_00000256AA0D38B0 [5]));  // al_ip/div_signed_gate.v(948)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_SIGNED/al_00000256AA4D4B20  (
    .a(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .b(\u_DIV_SIGNED/al_00000256AA8940C0 ),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D29D0 [1]),
    .o(\u_DIV_SIGNED/al_00000256AA0D38B0 [1]));  // al_ip/div_signed_gate.v(984)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_SIGNED/al_00000256AA4D4E50  (
    .a(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .b(\u_DIV_SIGNED/al_00000256AA8940C0 ),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D29D0 [3]),
    .o(\u_DIV_SIGNED/al_00000256AA0D38B0 [3]));  // al_ip/div_signed_gate.v(966)
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'b0001))
    \u_DIV_SIGNED/al_00000256AA4D58F0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CE7C0 [1]),
    .b(\u_DIV_SIGNED/al_00000256AA0CE7C0 [2]),
    .o(\u_DIV_SIGNED/al_00000256AA895350 ));  // al_ip/div_signed_gate.v(921)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_SIGNED/al_00000256AA4D5E40  (
    .a(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .b(\u_DIV_SIGNED/al_00000256AA8940C0 ),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D29D0 [4]),
    .o(\u_DIV_SIGNED/al_00000256AA0D38B0 [4]));  // al_ip/div_signed_gate.v(957)
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~B*~A))"),
    .INIT(16'b1111000111110000))
    \u_DIV_SIGNED/al_00000256AA4D5F50  (
    .a(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .b(\u_DIV_SIGNED/al_00000256AA8940C0 ),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D29D0 [0]),
    .o(\u_DIV_SIGNED/al_00000256AA0D38B0 [0]));  // al_ip/div_signed_gate.v(1001)
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'b00000000000000000000000000000010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4D6280  (
    .a(\u_DIV_SIGNED/al_00000256AA895350 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CE7C0 [0]),
    .c(\u_DIV_SIGNED/al_00000256AA0CE7C0 [3]),
    .d(\u_DIV_SIGNED/al_00000256AA0CE7C0 [4]),
    .e(\u_DIV_SIGNED/al_00000256AA0CE7C0 [5]),
    .o(\u_DIV_SIGNED/al_00000256AA8940C0 ));  // al_ip/div_signed_gate.v(938)
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'b00000000000010000000000000000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4D6390  (
    .a(\u_DIV_SIGNED/al_00000256AA895350 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CE7C0 [0]),
    .c(\u_DIV_SIGNED/al_00000256AA0CE7C0 [3]),
    .d(\u_DIV_SIGNED/al_00000256AA0CE7C0 [4]),
    .e(\u_DIV_SIGNED/al_00000256AA0CE7C0 [5]),
    .o(\u_DIV_SIGNED/al_00000256AA3DD9A0 ));  // al_ip/div_signed_gate.v(928)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4D6D20  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [9]),
    .b(n35[31]),
    .c(n35[9]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [9]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [9]));  // al_ip/div_signed_gate.v(911)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D7490  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [17]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [17]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [17]));  // al_ip/div_signed_gate.v(1353)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D75A0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [28]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [28]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [28]));  // al_ip/div_signed_gate.v(1065)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D76B0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [5]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [5]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [5]));  // al_ip/div_signed_gate.v(1121)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D77C0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [14]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [14]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [14]));  // al_ip/div_signed_gate.v(1385)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D78D0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [7]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [7]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [7]));  // al_ip/div_signed_gate.v(1177)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D79E0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [10]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [10]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [10]));  // al_ip/div_signed_gate.v(1417)
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'b0110))
    \u_DIV_SIGNED/al_00000256AA4D7AF0  (
    .a(n34[31]),
    .b(n35[31]),
    .o(\u_DIV_SIGNED/al_00000256AA422680 ));  // al_ip/div_signed_gate.v(301)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D7C00  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [31]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [31]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [31]));  // al_ip/div_signed_gate.v(1097)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D7D10  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [0]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [0]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [0]));  // al_ip/div_signed_gate.v(1113)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D7E20  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [9]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [9]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [9]));  // al_ip/div_signed_gate.v(1153)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D7F30  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [21]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [21]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [21]));  // al_ip/div_signed_gate.v(1313)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D8040  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [20]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [20]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [20]));  // al_ip/div_signed_gate.v(1321)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D8150  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [13]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [13]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [13]));  // al_ip/div_signed_gate.v(1393)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D8260  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [13]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [13]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [13]));  // al_ip/div_signed_gate.v(1579)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D8370  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [30]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [30]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [30]));  // al_ip/div_signed_gate.v(1225)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D8480  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [25]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [25]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [25]));  // al_ip/div_signed_gate.v(1273)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D8590  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [26]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [26]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [26]));  // al_ip/div_signed_gate.v(1049)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D86A0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [24]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [24]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [24]));  // al_ip/div_signed_gate.v(1281)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D87B0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [2]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [2]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [2]));  // al_ip/div_signed_gate.v(1329)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D88C0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [12]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [12]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [12]));  // al_ip/div_signed_gate.v(1401)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D89D0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [23]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [23]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [23]));  // al_ip/div_signed_gate.v(1018)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D8AE0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [4]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [4]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [4]));  // al_ip/div_signed_gate.v(1105)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D8BF0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [8]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [8]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [8]));  // al_ip/div_signed_gate.v(1169)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D8D00  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [9]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [9]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [9]));  // al_ip/div_signed_gate.v(1161)
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'b1000))
    \u_DIV_SIGNED/al_00000256AA4D8E10  (
    .a(n34[31]),
    .b(\u_DIV_SIGNED/al_00000256AA0D5590 [31]),
    .o(\u_DIV_SIGNED/al_00000256AA0D7970 [62]));  // al_ip/div_signed_gate.v(1026)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D8F20  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [16]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [16]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [16]));  // al_ip/div_signed_gate.v(406)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9030  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [18]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [18]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [18]));  // al_ip/div_signed_gate.v(602)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9140  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [19]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [19]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [19]));  // al_ip/div_signed_gate.v(700)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9250  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [25]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [25]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [25]));  // al_ip/div_signed_gate.v(1041)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9360  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [27]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [27]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [27]));  // al_ip/div_signed_gate.v(1057)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9470  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [1]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [1]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [1]));  // al_ip/div_signed_gate.v(1201)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9580  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [17]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [17]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [17]));  // al_ip/div_signed_gate.v(504)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9690  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [2]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [2]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [2]));  // al_ip/div_signed_gate.v(797)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D97A0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [24]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [24]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [24]));  // al_ip/div_signed_gate.v(1033)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D98B0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [6]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [6]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [6]));  // al_ip/div_signed_gate.v(1185)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D99C0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [31]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [31]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [31]));  // al_ip/div_signed_gate.v(1217)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4D9AD0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [14]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [14]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [14]));  // al_ip/div_signed_gate.v(1687)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D9BE0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [3]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [3]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [3]));  // al_ip/div_signed_gate.v(1233)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D9CF0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [28]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [28]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [28]));  // al_ip/div_signed_gate.v(1249)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D9E00  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [27]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [27]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [27]));  // al_ip/div_signed_gate.v(1257)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4D9F10  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [23]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [23]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [23]));  // al_ip/div_signed_gate.v(1297)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DA020  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [26]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [26]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [26]));  // al_ip/div_signed_gate.v(1265)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DA130  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [22]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [22]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [22]));  // al_ip/div_signed_gate.v(1305)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DA240  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [7]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [7]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [7]));  // al_ip/div_signed_gate.v(1137)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DA350  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [19]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [19]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [19]));  // al_ip/div_signed_gate.v(1337)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DA460  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [3]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [3]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [3]));  // al_ip/div_signed_gate.v(1081)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DA570  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [30]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [30]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [30]));  // al_ip/div_signed_gate.v(1089)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DA680  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [5]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [5]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [5]));  // al_ip/div_signed_gate.v(1193)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DA790  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [22]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [22]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [22]));  // al_ip/div_signed_gate.v(1010)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DA8A0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [18]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [18]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [18]));  // al_ip/div_signed_gate.v(1345)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DA9B0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [15]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [15]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [15]));  // al_ip/div_signed_gate.v(308)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DAAC0  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [16]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [16]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [16]));  // al_ip/div_signed_gate.v(1361)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DABD0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [29]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [29]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [29]));  // al_ip/div_signed_gate.v(1073)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DACE0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [12]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [12]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [12]));  // al_ip/div_signed_gate.v(1471)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DADF0  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [11]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [11]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [11]));  // al_ip/div_signed_gate.v(1377)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DAF00  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [8]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [8]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [8]));  // al_ip/div_signed_gate.v(1145)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DB010  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [20]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [20]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [20]));  // al_ip/div_signed_gate.v(895)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DB120  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [4]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [4]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [4]));  // al_ip/div_signed_gate.v(1209)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DB230  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [21]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [21]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [21]));  // al_ip/div_signed_gate.v(993)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DB340  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [29]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [29]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [29]));  // al_ip/div_signed_gate.v(1241)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DB450  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [15]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [15]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [15]));  // al_ip/div_signed_gate.v(1369)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DB560  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [11]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [11]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [11]));  // al_ip/div_signed_gate.v(1409)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DB670  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [10]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [10]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [10]));  // al_ip/div_signed_gate.v(1289)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_SIGNED/al_00000256AA4DB780  (
    .a(\u_DIV_SIGNED/al_00000256AA4072E0 [6]),
    .b(\u_DIV_SIGNED/al_00000256AA3DC030 ),
    .c(\u_DIV_SIGNED/al_00000256AA0CEB40 [6]),
    .o(\u_DIV_SIGNED/al_00000256AA4073C0 [6]));  // al_ip/div_signed_gate.v(1129)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DB890  (
    .a(n34[31]),
    .b(n34[5]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [5]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [37]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [36]));  // al_ip/div_signed_gate.v(1725)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DB9A0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [10]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [10]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [10]));  // al_ip/div_signed_gate.v(334)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DBAB0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [14]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [14]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [14]));  // al_ip/div_signed_gate.v(414)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DBBC0  (
    .a(n34[31]),
    .b(n34[15]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [15]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [47]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [46]));  // al_ip/div_signed_gate.v(1519)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DBCD0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [20]),
    .b(n35[31]),
    .c(n35[20]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [20]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [20]));  // al_ip/div_signed_gate.v(556)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DBDE0  (
    .a(n34[31]),
    .b(n34[29]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [29]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [61]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [60]));  // al_ip/div_signed_gate.v(1677)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DBEF0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [16]),
    .b(n35[31]),
    .c(n35[16]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [16]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [16]));  // al_ip/div_signed_gate.v(458)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DC000  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [17]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [17]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [17]));  // al_ip/div_signed_gate.v(468)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DC110  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [19]),
    .b(n35[31]),
    .c(n35[19]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [19]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [19]));  // al_ip/div_signed_gate.v(520)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DC220  (
    .a(n34[31]),
    .b(n34[30]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [30]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [62]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [61]));  // al_ip/div_signed_gate.v(1705)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DC330  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [2]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [2]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [2]));  // al_ip/div_signed_gate.v(530)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DC440  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [20]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [20]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [20]));  // al_ip/div_signed_gate.v(548)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DC550  (
    .a(n34[31]),
    .b(n34[11]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [11]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [43]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [42]));  // al_ip/div_signed_gate.v(1479)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DC660  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [0]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [0]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [0]));  // al_ip/div_signed_gate.v(1775)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DC770  (
    .a(n34[31]),
    .b(n34[1]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [1]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [33]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [32]));  // al_ip/div_signed_gate.v(1451)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DC880  (
    .a(n34[31]),
    .b(n34[8]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [8]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [40]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [39]));  // al_ip/div_signed_gate.v(1755)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DC990  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [15]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [15]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [15]));  // al_ip/div_signed_gate.v(432)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DCAA0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [21]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [21]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [21]));  // al_ip/div_signed_gate.v(566)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DCBB0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [21]),
    .b(n35[31]),
    .c(n35[21]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [21]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [21]));  // al_ip/div_signed_gate.v(574)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DCCC0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [22]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [22]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [22]));  // al_ip/div_signed_gate.v(584)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DCDD0  (
    .a(n34[31]),
    .b(n34[12]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [12]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [44]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [43]));  // al_ip/div_signed_gate.v(1489)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DCEE0  (
    .a(n34[31]),
    .b(n34[10]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [10]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [42]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [41]));  // al_ip/div_signed_gate.v(1461)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DCFF0  (
    .a(n34[31]),
    .b(n34[16]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [16]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [48]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [47]));  // al_ip/div_signed_gate.v(1529)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DD100  (
    .a(n34[31]),
    .b(n34[18]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [18]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [50]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [49]));  // al_ip/div_signed_gate.v(1549)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DD210  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [12]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [12]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [12]));  // al_ip/div_signed_gate.v(370)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DD320  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [1]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [1]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [1]));  // al_ip/div_signed_gate.v(1425)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DD430  (
    .a(n34[31]),
    .b(n34[27]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [27]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [59]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [58]));  // al_ip/div_signed_gate.v(1657)
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'b10101100))
    \u_DIV_SIGNED/al_00000256AA4DD540  (
    .a(\u_DIV_SIGNED/al_00000256AA40B170 [0]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [0]),
    .c(\u_DIV_SIGNED/al_00000256AA3DC5B0 ),
    .o(\u_DIV_SIGNED/al_00000256AA4098F0 [0]));  // al_ip/div_signed_gate.v(1433)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DD650  (
    .a(n34[31]),
    .b(n34[3]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [3]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [35]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [34]));  // al_ip/div_signed_gate.v(1695)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DD760  (
    .a(n34[31]),
    .b(n34[7]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [7]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [39]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [38]));  // al_ip/div_signed_gate.v(1745)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DD870  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [0]),
    .b(n35[31]),
    .c(n35[0]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [0]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [0]));  // al_ip/div_signed_gate.v(1783)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DD980  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [10]),
    .b(n35[31]),
    .c(n35[10]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [10]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [10]));  // al_ip/div_signed_gate.v(342)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DDA90  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [1]),
    .b(n35[31]),
    .c(n35[1]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [1]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [1]));  // al_ip/div_signed_gate.v(324)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DDBA0  (
    .a(n34[31]),
    .b(n34[13]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [13]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [45]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [44]));  // al_ip/div_signed_gate.v(1499)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DDCB0  (
    .a(n34[31]),
    .b(n34[6]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [6]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [38]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [37]));  // al_ip/div_signed_gate.v(1735)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DDDC0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [11]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [11]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [11]));  // al_ip/div_signed_gate.v(352)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DDED0  (
    .a(n34[31]),
    .b(n34[14]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [14]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [46]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [45]));  // al_ip/div_signed_gate.v(1509)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DDFE0  (
    .a(n34[31]),
    .b(n34[17]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [17]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [49]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [48]));  // al_ip/div_signed_gate.v(1539)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE0F0  (
    .a(n34[31]),
    .b(n34[25]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [25]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [57]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [56]));  // al_ip/div_signed_gate.v(1637)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE200  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [12]),
    .b(n35[31]),
    .c(n35[12]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [12]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [12]));  // al_ip/div_signed_gate.v(378)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DE310  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [13]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [13]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [13]));  // al_ip/div_signed_gate.v(388)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE420  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [14]),
    .b(n35[31]),
    .c(n35[14]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [14]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [14]));  // al_ip/div_signed_gate.v(422)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DE530  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [18]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [18]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [18]));  // al_ip/div_signed_gate.v(486)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE640  (
    .a(n34[31]),
    .b(n34[0]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [0]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [32]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [31]));  // al_ip/div_signed_gate.v(1441)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE750  (
    .a(n34[31]),
    .b(n34[19]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [19]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [51]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [50]));  // al_ip/div_signed_gate.v(1559)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE860  (
    .a(n34[31]),
    .b(n34[2]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [2]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [34]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [33]));  // al_ip/div_signed_gate.v(1569)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DE970  (
    .a(n34[31]),
    .b(n34[21]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [21]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [53]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [52]));  // al_ip/div_signed_gate.v(1597)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DEA80  (
    .a(n34[31]),
    .b(n34[23]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [23]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [55]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [54]));  // al_ip/div_signed_gate.v(1617)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DEB90  (
    .a(n34[31]),
    .b(n34[22]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [22]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [54]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [53]));  // al_ip/div_signed_gate.v(1607)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DECA0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [1]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [1]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [1]));  // al_ip/div_signed_gate.v(316)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DEDB0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [11]),
    .b(n35[31]),
    .c(n35[11]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [11]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [11]));  // al_ip/div_signed_gate.v(360)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DEEC0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [15]),
    .b(n35[31]),
    .c(n35[15]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [15]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [15]));  // al_ip/div_signed_gate.v(440)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DEFD0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [16]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [16]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [16]));  // al_ip/div_signed_gate.v(450)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF0E0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [17]),
    .b(n35[31]),
    .c(n35[17]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [17]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [17]));  // al_ip/div_signed_gate.v(476)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF1F0  (
    .a(n34[31]),
    .b(n34[24]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [24]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [56]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [55]));  // al_ip/div_signed_gate.v(1627)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF300  (
    .a(n34[31]),
    .b(n34[4]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [4]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [36]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [35]));  // al_ip/div_signed_gate.v(1715)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF410  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [18]),
    .b(n35[31]),
    .c(n35[18]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [18]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [18]));  // al_ip/div_signed_gate.v(494)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF520  (
    .a(n34[31]),
    .b(n34[28]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [28]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [60]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [59]));  // al_ip/div_signed_gate.v(1667)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF630  (
    .a(n34[31]),
    .b(n34[9]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [9]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [41]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [40]));  // al_ip/div_signed_gate.v(1765)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF740  (
    .a(n34[31]),
    .b(n34[20]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [20]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [52]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [51]));  // al_ip/div_signed_gate.v(1587)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DF850  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [13]),
    .b(n35[31]),
    .c(n35[13]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [13]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [13]));  // al_ip/div_signed_gate.v(396)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DF960  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [19]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [19]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [19]));  // al_ip/div_signed_gate.v(512)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DFA70  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [2]),
    .b(n35[31]),
    .c(n35[2]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [2]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [2]));  // al_ip/div_signed_gate.v(538)
  AL_MAP_LUT5 #(
    .EQN("(E*~((B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A))*~(C)+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*~(C)+~(E)*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C+E*(B*~(D)*~(A)+B*D*~(A)+~(B)*D*A+B*D*A)*C)"),
    .INIT(32'b11101111010011111110000001000000),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DFB80  (
    .a(n34[31]),
    .b(n34[26]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA0D5590 [26]),
    .e(\u_DIV_SIGNED/al_00000256AA0D0BA0 [58]),
    .o(\u_DIV_SIGNED/al_00000256AA0D80E0 [57]));  // al_ip/div_signed_gate.v(1647)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4DFC90  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [24]),
    .b(n35[31]),
    .c(n35[24]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [24]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [24]));  // al_ip/div_signed_gate.v(636)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DFDA0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [26]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [26]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [26]));  // al_ip/div_signed_gate.v(664)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DFEB0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [27]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [27]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [27]));  // al_ip/div_signed_gate.v(682)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4DFFC0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [30]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [30]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [30]));  // al_ip/div_signed_gate.v(762)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E00D0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [29]),
    .b(n35[31]),
    .c(n35[29]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [29]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [29]));  // al_ip/div_signed_gate.v(734)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E02F0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [28]),
    .b(n35[31]),
    .c(n35[28]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [28]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [28]));  // al_ip/div_signed_gate.v(716)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0400  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [25]),
    .b(n35[31]),
    .c(n35[25]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [25]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [25]));  // al_ip/div_signed_gate.v(654)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E0620  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [28]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [28]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [28]));  // al_ip/div_signed_gate.v(708)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E0730  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [3]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [3]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [3]));  // al_ip/div_signed_gate.v(744)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0840  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [30]),
    .b(n35[31]),
    .c(n35[30]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [30]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [30]));  // al_ip/div_signed_gate.v(770)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0950  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [3]),
    .b(n35[31]),
    .c(n35[3]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [3]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [3]));  // al_ip/div_signed_gate.v(752)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E0A60  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [4]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [4]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [4]));  // al_ip/div_signed_gate.v(805)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0B70  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [4]),
    .b(n35[31]),
    .c(n35[4]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [4]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [4]));  // al_ip/div_signed_gate.v(813)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0C80  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [5]),
    .b(n35[31]),
    .c(n35[5]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [5]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [5]));  // al_ip/div_signed_gate.v(831)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0D90  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [6]),
    .b(n35[31]),
    .c(n35[6]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [6]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [6]));  // al_ip/div_signed_gate.v(849)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E0EA0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [7]),
    .b(n35[31]),
    .c(n35[7]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [7]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [7]));  // al_ip/div_signed_gate.v(867)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E0FB0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [8]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [8]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [8]));  // al_ip/div_signed_gate.v(877)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E10C0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [9]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [9]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [9]));  // al_ip/div_signed_gate.v(903)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E11D0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [8]),
    .b(n35[31]),
    .c(n35[8]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [8]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [8]));  // al_ip/div_signed_gate.v(885)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E12E0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [29]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [29]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [29]));  // al_ip/div_signed_gate.v(726)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E13F0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [23]),
    .b(n35[31]),
    .c(n35[23]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [23]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [23]));  // al_ip/div_signed_gate.v(618)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E1500  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [26]),
    .b(n35[31]),
    .c(n35[26]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [26]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [26]));  // al_ip/div_signed_gate.v(672)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E1610  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [5]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [5]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [5]));  // al_ip/div_signed_gate.v(823)
  AL_MAP_LUT4 #(
    .EQN("(~A*~((D*B))*~(C)+~A*(D*B)*~(C)+~(~A)*(D*B)*C+~A*(D*B)*C)"),
    .INIT(16'b1100010100000101))
    \u_DIV_SIGNED/al_00000256AA4E1720  (
    .a(\u_DIV_SIGNED/al_00000256AA893670 ),
    .b(n35[31]),
    .c(div_signed_start),
    .d(\u_DIV_SIGNED/al_00000256AA3FF0F0 [31]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [31]));  // al_ip/div_signed_gate.v(788)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E1830  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [6]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [6]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [6]));  // al_ip/div_signed_gate.v(841)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E1B60  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [7]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [7]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [7]));  // al_ip/div_signed_gate.v(859)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E1D80  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [23]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [23]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [23]));  // al_ip/div_signed_gate.v(610)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E20B0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [25]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [25]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [25]));  // al_ip/div_signed_gate.v(646)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E21C0  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [27]),
    .b(n35[31]),
    .c(n35[27]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [27]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [27]));  // al_ip/div_signed_gate.v(690)
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b11100100))
    \u_DIV_SIGNED/al_00000256AA4E22D0  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [24]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [24]),
    .o(\u_DIV_SIGNED/al_00000256AA403450 [24]));  // al_ip/div_signed_gate.v(628)
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'b00011011))
    \u_DIV_SIGNED/al_00000256AA4E2710  (
    .a(\u_DIV_SIGNED/al_00000256AA3DB7F0 ),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [31]),
    .c(\u_DIV_SIGNED/al_00000256AA400D60 [31]),
    .o(\u_DIV_SIGNED/al_00000256AA893670 ));  // al_ip/div_signed_gate.v(780)
  AL_MAP_LUT5 #(
    .EQN("(A*~((C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B))*~(D)+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*~(D)+~(A)*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D+A*(C*~(E)*~(B)+C*E*~(B)+~(C)*E*B+C*E*B)*D)"),
    .INIT(32'b11111100101010100011000010101010),
    .LOC("UNPLACED"))
    \u_DIV_SIGNED/al_00000256AA4E2B50  (
    .a(\u_DIV_SIGNED/al_00000256AA403450 [22]),
    .b(n35[31]),
    .c(n35[22]),
    .d(div_signed_start),
    .e(\u_DIV_SIGNED/al_00000256AA3FF0F0 [22]),
    .o(\u_DIV_SIGNED/al_00000256AA402C70 [22]));  // al_ip/div_signed_gate.v(592)
  EG_PHY_LSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256A66FB850_al_u414"),
    //.R_POSITION("X0Y3Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6691B0_al_u420  (
    .a({\u_DIV_SIGNED/al_00000256AA0CF470 [25],\u_DIV_SIGNED/al_00000256AA0CF470 [23]}),
    .b({\u_DIV_SIGNED/al_00000256AA0CF470 [26],\u_DIV_SIGNED/al_00000256AA0CF470 [24]}),
    .c(2'b11),
    .d({\u_DIV_SIGNED/al_00000256AA0D0BA0 [25],\u_DIV_SIGNED/al_00000256AA0D0BA0 [23]}),
    .e({\u_DIV_SIGNED/al_00000256AA0D0BA0 [26],\u_DIV_SIGNED/al_00000256AA0D0BA0 [24]}),
    .fci(\u_DIV_SIGNED/al_00000256AA898E70 ),
    .f({\u_DIV_SIGNED/al_00000256AA400D60 [25],\u_DIV_SIGNED/al_00000256AA400D60 [23]}),
    .fco(\u_DIV_SIGNED/al_00000256AA898630 ),
    .fx({\u_DIV_SIGNED/al_00000256AA400D60 [26],\u_DIV_SIGNED/al_00000256AA400D60 [24]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256A66FB850_al_u414"),
    //.R_POSITION("X0Y3Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6695F0_al_u421  (
    .a({\u_DIV_SIGNED/al_00000256AA0CF470 [29],\u_DIV_SIGNED/al_00000256AA0CF470 [27]}),
    .b({\u_DIV_SIGNED/al_00000256AA0CF470 [30],\u_DIV_SIGNED/al_00000256AA0CF470 [28]}),
    .c(2'b11),
    .d({\u_DIV_SIGNED/al_00000256AA0D0BA0 [29],\u_DIV_SIGNED/al_00000256AA0D0BA0 [27]}),
    .e({\u_DIV_SIGNED/al_00000256AA0D0BA0 [30],\u_DIV_SIGNED/al_00000256AA0D0BA0 [28]}),
    .fci(\u_DIV_SIGNED/al_00000256AA898630 ),
    .f({\u_DIV_SIGNED/al_00000256AA400D60 [29],\u_DIV_SIGNED/al_00000256AA400D60 [27]}),
    .fco(\u_DIV_SIGNED/al_00000256AA899810 ),
    .fx({\u_DIV_SIGNED/al_00000256AA400D60 [30],\u_DIV_SIGNED/al_00000256AA400D60 [28]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256A66FB850_al_u414"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA66A090_al_u415  (
    .a({\u_DIV_SIGNED/al_00000256AA0CF470 [5],\u_DIV_SIGNED/al_00000256AA0CF470 [3]}),
    .b({\u_DIV_SIGNED/al_00000256AA0CF470 [6],\u_DIV_SIGNED/al_00000256AA0CF470 [4]}),
    .c(2'b11),
    .d({\u_DIV_SIGNED/al_00000256AA0D0BA0 [5],\u_DIV_SIGNED/al_00000256AA0D0BA0 [3]}),
    .e({\u_DIV_SIGNED/al_00000256AA0D0BA0 [6],\u_DIV_SIGNED/al_00000256AA0D0BA0 [4]}),
    .fci(\u_DIV_SIGNED/al_00000256AA898FD0 ),
    .f({\u_DIV_SIGNED/al_00000256AA400D60 [5],\u_DIV_SIGNED/al_00000256AA400D60 [3]}),
    .fco(\u_DIV_SIGNED/al_00000256AA89AEC0 ),
    .fx({\u_DIV_SIGNED/al_00000256AA400D60 [6],\u_DIV_SIGNED/al_00000256AA400D60 [4]}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA66A1A0  (
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA3DD9A0 ),
    .sr(i_rstn),
    .q(div_signed_finish));  // al_ip/div_signed_gate.v(2753)
  EG_PHY_LSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256A66FB850_al_u414"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA66A800_al_u418  (
    .a({\u_DIV_SIGNED/al_00000256AA0CF470 [17],\u_DIV_SIGNED/al_00000256AA0CF470 [15]}),
    .b({\u_DIV_SIGNED/al_00000256AA0CF470 [18],\u_DIV_SIGNED/al_00000256AA0CF470 [16]}),
    .c(2'b11),
    .d({\u_DIV_SIGNED/al_00000256AA0D0BA0 [17],\u_DIV_SIGNED/al_00000256AA0D0BA0 [15]}),
    .e({\u_DIV_SIGNED/al_00000256AA0D0BA0 [18],\u_DIV_SIGNED/al_00000256AA0D0BA0 [16]}),
    .fci(\u_DIV_SIGNED/al_00000256AA899130 ),
    .f({\u_DIV_SIGNED/al_00000256AA400D60 [17],\u_DIV_SIGNED/al_00000256AA400D60 [15]}),
    .fco(\u_DIV_SIGNED/al_00000256AA898DC0 ),
    .fx({\u_DIV_SIGNED/al_00000256AA400D60 [18],\u_DIV_SIGNED/al_00000256AA400D60 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256A66FB850_al_u414"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA66AD50_al_u419  (
    .a({\u_DIV_SIGNED/al_00000256AA0CF470 [21],\u_DIV_SIGNED/al_00000256AA0CF470 [19]}),
    .b({\u_DIV_SIGNED/al_00000256AA0CF470 [22],\u_DIV_SIGNED/al_00000256AA0CF470 [20]}),
    .c(2'b11),
    .d({\u_DIV_SIGNED/al_00000256AA0D0BA0 [21],\u_DIV_SIGNED/al_00000256AA0D0BA0 [19]}),
    .e({\u_DIV_SIGNED/al_00000256AA0D0BA0 [22],\u_DIV_SIGNED/al_00000256AA0D0BA0 [20]}),
    .fci(\u_DIV_SIGNED/al_00000256AA898DC0 ),
    .f({\u_DIV_SIGNED/al_00000256AA400D60 [21],\u_DIV_SIGNED/al_00000256AA400D60 [19]}),
    .fco(\u_DIV_SIGNED/al_00000256AA898E70 ),
    .fx({\u_DIV_SIGNED/al_00000256AA400D60 [22],\u_DIV_SIGNED/al_00000256AA400D60 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256A66FB850_al_u414"),
    //.R_POSITION("X0Y4Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA66B080_al_u422  (
    .a({open_n2719,\u_DIV_SIGNED/al_00000256AA0CF470 [31]}),
    .c(2'b11),
    .d({open_n2724,\u_DIV_SIGNED/al_00000256AA0D0BA0 [31]}),
    .fci(\u_DIV_SIGNED/al_00000256AA899810 ),
    .f({open_n2741,\u_DIV_SIGNED/al_00000256AA400D60 [31]}));
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_SIGNED/al_00000256AA66B190  (
    .ce(div_signed_start),
    .clk(i_clk),
    .d(\u_DIV_SIGNED/al_00000256AA422680 ),
    .q(\u_DIV_SIGNED/al_00000256AA3DC030 ));  // al_ip/div_signed_gate.v(3215)
  EG_PHY_LSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256A66FB850_al_u414"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA66C6D0_al_u417  (
    .a({\u_DIV_SIGNED/al_00000256AA0CF470 [13],\u_DIV_SIGNED/al_00000256AA0CF470 [11]}),
    .b({\u_DIV_SIGNED/al_00000256AA0CF470 [14],\u_DIV_SIGNED/al_00000256AA0CF470 [12]}),
    .c(2'b11),
    .d({\u_DIV_SIGNED/al_00000256AA0D0BA0 [13],\u_DIV_SIGNED/al_00000256AA0D0BA0 [11]}),
    .e({\u_DIV_SIGNED/al_00000256AA0D0BA0 [14],\u_DIV_SIGNED/al_00000256AA0D0BA0 [12]}),
    .fci(\u_DIV_SIGNED/al_00000256AA899290 ),
    .f({\u_DIV_SIGNED/al_00000256AA400D60 [13],\u_DIV_SIGNED/al_00000256AA400D60 [11]}),
    .fco(\u_DIV_SIGNED/al_00000256AA899130 ),
    .fx({\u_DIV_SIGNED/al_00000256AA400D60 [14],\u_DIV_SIGNED/al_00000256AA400D60 [12]}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \u_DIV_SIGNED/al_00000256AA66ED10  (
    .clk(i_clk),
    .d(i_mdu_op1[31]),
    .sr(mdu_vld),
    .q(\u_DIV_SIGNED/al_00000256AA3DC5B0 ));  // al_ip/div_signed_gate.v(4997)
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA672780|u_DIV_SIGNED/al_00000256AA672670"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA672780|u_DIV_SIGNED/al_00000256AA672670  (
    .a({\u_DIV_SIGNED/al_00000256AA0CE7C0 [0],1'b0}),
    .b(2'b10),
    .f({\u_DIV_SIGNED/al_00000256AA0D29D0 [0],open_n2786}),
    .fco(\u_DIV_SIGNED/al_00000256AA6547B0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA672780|u_DIV_SIGNED/al_00000256AA672670"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA672DE0_al_u425  (
    .a({open_n2791,\u_DIV_SIGNED/al_00000256AA0CE7C0 [5]}),
    .b({open_n2792,1'b0}),
    .fci(\u_DIV_SIGNED/al_00000256AA653E10 ),
    .f({open_n2811,\u_DIV_SIGNED/al_00000256AA0D29D0 [5]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA672780|u_DIV_SIGNED/al_00000256AA672670"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA673880|u_DIV_SIGNED/al_00000256AA675200  (
    .a(\u_DIV_SIGNED/al_00000256AA0CE7C0 [4:3]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA653890 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D29D0 [4:3]),
    .fco(\u_DIV_SIGNED/al_00000256AA653E10 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA672780|u_DIV_SIGNED/al_00000256AA672670"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA675750|u_DIV_SIGNED/al_00000256AA672BC0  (
    .a(\u_DIV_SIGNED/al_00000256AA0CE7C0 [2:1]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA6547B0 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D29D0 [2:1]),
    .fco(\u_DIV_SIGNED/al_00000256AA653890 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA675FD0|u_DIV_SIGNED/al_00000256AA678610  (
    .a(2'b00),
    .b(n34[12:11]),
    .fci(\u_DIV_SIGNED/al_00000256AA423390 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [12:11]),
    .fco(\u_DIV_SIGNED/al_00000256AA422E10 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6760E0|u_DIV_SIGNED/al_00000256AA677D90  (
    .a(2'b00),
    .b(n34[28:27]),
    .fci(\u_DIV_SIGNED/al_00000256AA421CE0 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [28:27]),
    .fco(\u_DIV_SIGNED/al_00000256AA4216B0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA676A70|u_DIV_SIGNED/al_00000256AA679600  (
    .a(2'b00),
    .b(n34[10:9]),
    .fci(\u_DIV_SIGNED/al_00000256AA4232E0 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [10:9]),
    .fco(\u_DIV_SIGNED/al_00000256AA423390 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA676B80|u_DIV_SIGNED/al_00000256AA6772F0  (
    .a(2'b00),
    .b(n34[20:19]),
    .fci(\u_DIV_SIGNED/al_00000256AA421130 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [20:19]),
    .fco(\u_DIV_SIGNED/al_00000256AA421550 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA676C90|u_DIV_SIGNED/al_00000256AA678720  (
    .a(2'b00),
    .b(n34[22:21]),
    .fci(\u_DIV_SIGNED/al_00000256AA421550 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [22:21]),
    .fco(\u_DIV_SIGNED/al_00000256AA423700 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA676DA0|u_DIV_SIGNED/al_00000256AA676520  (
    .a(2'b00),
    .b(n34[8:7]),
    .fci(\u_DIV_SIGNED/al_00000256AA422470 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [8:7]),
    .fco(\u_DIV_SIGNED/al_00000256AA4232E0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6771E0|u_DIV_SIGNED/al_00000256AA6790B0  (
    .a(2'b00),
    .b(n34[26:25]),
    .fci(\u_DIV_SIGNED/al_00000256AA422310 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [26:25]),
    .fco(\u_DIV_SIGNED/al_00000256AA421CE0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA677400|u_DIV_SIGNED/al_00000256AA678FA0  (
    .a(2'b00),
    .b(n34[16:15]),
    .fci(\u_DIV_SIGNED/al_00000256AA422940 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [16:15]),
    .fco(\u_DIV_SIGNED/al_00000256AA421080 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6782E0|u_DIV_SIGNED/al_00000256AA677620  (
    .a(2'b00),
    .b(n34[18:17]),
    .fci(\u_DIV_SIGNED/al_00000256AA421080 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [18:17]),
    .fco(\u_DIV_SIGNED/al_00000256AA421130 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA678A50|u_DIV_SIGNED/al_00000256AA677510  (
    .a(2'b00),
    .b(n34[14:13]),
    .fci(\u_DIV_SIGNED/al_00000256AA422E10 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [14:13]),
    .fco(\u_DIV_SIGNED/al_00000256AA422940 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA678C70|u_DIV_SIGNED/al_00000256AA678B60  (
    .a(2'b00),
    .b(n34[2:1]),
    .fci(\u_DIV_SIGNED/al_00000256AA423B20 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [2:1]),
    .fco(\u_DIV_SIGNED/al_00000256AA4218C0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730  (
    .a(2'b00),
    .b({n34[0],1'b0}),
    .f({\u_DIV_SIGNED/al_00000256AA0D5590 [0],open_n3122}),
    .fco(\u_DIV_SIGNED/al_00000256AA423B20 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6791C0|u_DIV_SIGNED/al_00000256AA679710  (
    .a(2'b00),
    .b(n34[30:29]),
    .fci(\u_DIV_SIGNED/al_00000256AA4216B0 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [30:29]),
    .fco(\u_DIV_SIGNED/al_00000256AA421600 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6792D0_al_u426  (
    .a({open_n3149,1'b0}),
    .b({open_n3150,n34[31]}),
    .fci(\u_DIV_SIGNED/al_00000256AA421600 ),
    .f({open_n3169,\u_DIV_SIGNED/al_00000256AA0D5590 [31]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6793E0|u_DIV_SIGNED/al_00000256AA678D80  (
    .a(2'b00),
    .b(n34[24:23]),
    .fci(\u_DIV_SIGNED/al_00000256AA423700 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [24:23]),
    .fco(\u_DIV_SIGNED/al_00000256AA422310 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6794F0|u_DIV_SIGNED/al_00000256AA678500  (
    .a(2'b00),
    .b(n34[4:3]),
    .fci(\u_DIV_SIGNED/al_00000256AA4218C0 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [4:3]),
    .fco(\u_DIV_SIGNED/al_00000256AA421C30 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA678E90|u_DIV_SIGNED/al_00000256AA677730"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA679C60|u_DIV_SIGNED/al_00000256AA6783F0  (
    .a(2'b00),
    .b(n34[6:5]),
    .fci(\u_DIV_SIGNED/al_00000256AA421C30 ),
    .f(\u_DIV_SIGNED/al_00000256AA0D5590 [6:5]),
    .fco(\u_DIV_SIGNED/al_00000256AA422470 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67A1B0|u_DIV_SIGNED/al_00000256AA67D4B0  (
    .a(2'b00),
    .b(n35[2:1]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DD2C0 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [2:1]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DD840 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67B090|u_DIV_SIGNED/al_00000256AA67B910  (
    .a(2'b00),
    .b(n35[18:17]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DDA50 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [18:17]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DD420 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67B5E0|u_DIV_SIGNED/al_00000256AA67D5C0  (
    .a(2'b00),
    .b(n35[16:15]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DC450 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [16:15]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DDA50 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67BA20|u_DIV_SIGNED/al_00000256AA67B6F0  (
    .a(2'b00),
    .b(n35[6:5]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DB3D0 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [6:5]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DB480 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67C6E0|u_DIV_SIGNED/al_00000256AA67C7F0  (
    .a(2'b00),
    .b(n35[28:27]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DB320 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [28:27]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DC9D0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67CA10|u_DIV_SIGNED/al_00000256AA67C2A0  (
    .a(2'b00),
    .b(n35[24:23]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DB5E0 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [24:23]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DD580 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67CC30|u_DIV_SIGNED/al_00000256AA67B800  (
    .a(2'b00),
    .b(n35[22:21]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DCC90 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [22:21]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DB5E0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40  (
    .a(2'b00),
    .b({n35[0],1'b0}),
    .f({\u_DIV_SIGNED/al_00000256AA3FF0F0 [0],open_n3414}),
    .fco(\u_DIV_SIGNED/al_00000256AA3DD2C0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67D070|u_DIV_SIGNED/al_00000256AA67C900  (
    .a(2'b00),
    .b(n35[12:11]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DB110 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [12:11]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DC870 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67D290|u_DIV_SIGNED/al_00000256AA67BE60  (
    .a(2'b00),
    .b(n35[20:19]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DD420 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [20:19]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DCC90 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67D6D0|u_DIV_SIGNED/al_00000256AA67BB30  (
    .a(2'b00),
    .b(n35[26:25]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DD580 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [26:25]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DB320 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67D7E0|u_DIV_SIGNED/al_00000256AA67D180  (
    .a(2'b00),
    .b(n35[14:13]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DC870 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [14:13]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DC450 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67D8F0|u_DIV_SIGNED/al_00000256AA67DD30  (
    .a(2'b00),
    .b(n35[30:29]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DC9D0 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [30:29]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DDB00 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67DA00_al_u427  (
    .a({open_n3529,1'b0}),
    .b({open_n3530,n35[31]}),
    .fci(\u_DIV_SIGNED/al_00000256AA3DDB00 ),
    .f({open_n3549,\u_DIV_SIGNED/al_00000256AA3FF0F0 [31]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67DB10|u_DIV_SIGNED/al_00000256AA67DF50  (
    .a(2'b00),
    .b(n35[10:9]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DEA20 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [10:9]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DB110 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67DC20|u_DIV_SIGNED/al_00000256AA67E170  (
    .a(2'b00),
    .b(n35[4:3]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DD840 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [4:3]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DB3D0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA67CE50|u_DIV_SIGNED/al_00000256AA67CD40"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67DE40|u_DIV_SIGNED/al_00000256AA67CB20  (
    .a(2'b00),
    .b(n35[8:7]),
    .fci(\u_DIV_SIGNED/al_00000256AA3DB480 ),
    .f(\u_DIV_SIGNED/al_00000256AA3FF0F0 [8:7]),
    .fco(\u_DIV_SIGNED/al_00000256AA3DEA20 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67E5B0|u_DIV_SIGNED/al_00000256AA680260  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [8:7]),
    .fci(\u_DIV_SIGNED/al_00000256AA444E10 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [8:7]),
    .fco(\u_DIV_SIGNED/al_00000256AA3E0300 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67ED20|u_DIV_SIGNED/al_00000256AA67FD10  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [14:13]),
    .fci(\u_DIV_SIGNED/al_00000256AA443CE0 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [14:13]),
    .fco(\u_DIV_SIGNED/al_00000256AA443E40 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67F270|u_DIV_SIGNED/al_00000256AA67FC00  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [16:15]),
    .fci(\u_DIV_SIGNED/al_00000256AA443E40 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [16:15]),
    .fco(\u_DIV_SIGNED/al_00000256AA443760 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67F5A0|u_DIV_SIGNED/al_00000256AA67EC10  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [2:1]),
    .fci(\u_DIV_SIGNED/al_00000256AA445230 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [2:1]),
    .fco(\u_DIV_SIGNED/al_00000256AA444CB0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67F6B0|u_DIV_SIGNED/al_00000256AA67F050  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [20:19]),
    .fci(\u_DIV_SIGNED/al_00000256AA443810 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [20:19]),
    .fco(\u_DIV_SIGNED/al_00000256AA444680 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67F8D0|u_DIV_SIGNED/al_00000256AA67F160  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [24:23]),
    .fci(\u_DIV_SIGNED/al_00000256AA444100 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [24:23]),
    .fco(\u_DIV_SIGNED/al_00000256AA443130 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67F9E0|u_DIV_SIGNED/al_00000256AA67EF40  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [22:21]),
    .fci(\u_DIV_SIGNED/al_00000256AA444680 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [22:21]),
    .fco(\u_DIV_SIGNED/al_00000256AA444100 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA67FAF0|u_DIV_SIGNED/al_00000256AA681CF0  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [10:9]),
    .fci(\u_DIV_SIGNED/al_00000256AA3E0300 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [10:9]),
    .fco(\u_DIV_SIGNED/al_00000256AA4436B0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA680150|u_DIV_SIGNED/al_00000256AA680040  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [30:29]),
    .fci(\u_DIV_SIGNED/al_00000256AA444260 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [30:29]),
    .fco(\u_DIV_SIGNED/al_00000256AA4445D0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240  (
    .a(2'b00),
    .b({\u_DIV_SIGNED/al_00000256AA0CEB40 [0],1'b0}),
    .f({\u_DIV_SIGNED/al_00000256AA4072E0 [0],open_n3838}),
    .fco(\u_DIV_SIGNED/al_00000256AA445230 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA680AE0|u_DIV_SIGNED/al_00000256AA682130  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [6:5]),
    .fci(\u_DIV_SIGNED/al_00000256AA444940 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [6:5]),
    .fco(\u_DIV_SIGNED/al_00000256AA444E10 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA680E10|u_DIV_SIGNED/al_00000256AA67FF30  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [28:27]),
    .fci(\u_DIV_SIGNED/al_00000256AA444B50 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [28:27]),
    .fco(\u_DIV_SIGNED/al_00000256AA444260 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA680F20|u_DIV_SIGNED/al_00000256AA67FE20  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [12:11]),
    .fci(\u_DIV_SIGNED/al_00000256AA4436B0 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [12:11]),
    .fco(\u_DIV_SIGNED/al_00000256AA443CE0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA681030_al_u428  (
    .a({open_n3909,1'b0}),
    .b({open_n3910,\u_DIV_SIGNED/al_00000256AA0CEB40 [31]}),
    .fci(\u_DIV_SIGNED/al_00000256AA4445D0 ),
    .f({open_n3929,\u_DIV_SIGNED/al_00000256AA4072E0 [31]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6817A0|u_DIV_SIGNED/al_00000256AA682460  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [26:25]),
    .fci(\u_DIV_SIGNED/al_00000256AA443130 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [26:25]),
    .fco(\u_DIV_SIGNED/al_00000256AA444B50 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6819C0|u_DIV_SIGNED/al_00000256AA682350  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [4:3]),
    .fci(\u_DIV_SIGNED/al_00000256AA444CB0 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [4:3]),
    .fco(\u_DIV_SIGNED/al_00000256AA444940 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA6807B0|u_DIV_SIGNED/al_00000256AA682240"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA682020|u_DIV_SIGNED/al_00000256AA6818B0  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CEB40 [18:17]),
    .fci(\u_DIV_SIGNED/al_00000256AA443760 ),
    .f(\u_DIV_SIGNED/al_00000256AA4072E0 [18:17]),
    .fco(\u_DIV_SIGNED/al_00000256AA443810 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6828A0|u_DIV_SIGNED/al_00000256AA686530  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [4:3]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [4:3]),
    .fci(\u_DIV_SIGNED/al_00000256AA88C450 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88ADA0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA682CE0|u_DIV_SIGNED/al_00000256AA684880  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [12:11]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [12:11]),
    .fci(\u_DIV_SIGNED/al_00000256AA88BCC0 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88A8D0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA683010|u_DIV_SIGNED/al_00000256AA684CC0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [16:15]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [16:15]),
    .fci(\u_DIV_SIGNED/al_00000256AA88C3A0 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88B110 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA683340|u_DIV_SIGNED/al_00000256AA683120  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [18:17]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [18:17]),
    .fci(\u_DIV_SIGNED/al_00000256AA88B110 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88B480 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA683450|u_DIV_SIGNED/al_00000256AA684BB0  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [6:5]),
    .fci(\u_DIV_SIGNED/al_00000256AA88B270 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [6:5]),
    .fco(\u_DIV_SIGNED/al_00000256AA88B530 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA683890|u_DIV_SIGNED/al_00000256AA686310  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [2:1]),
    .fci(\u_DIV_SIGNED/al_00000256AA88C190 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [2:1]),
    .fco(\u_DIV_SIGNED/al_00000256AA88AC40 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6839A0|u_DIV_SIGNED/al_00000256AA683670  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [8:7]),
    .fci(\u_DIV_SIGNED/al_00000256AA88B530 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [8:7]),
    .fco(\u_DIV_SIGNED/al_00000256AA88AF00 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA683AB0|u_DIV_SIGNED/al_00000256AA682F00  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [18:17]),
    .fci(\u_DIV_SIGNED/al_00000256AA88BED0 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [18:17]),
    .fco(\u_DIV_SIGNED/al_00000256AA88CEA0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA683BC0|u_DIV_SIGNED/al_00000256AA685870  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [6:5]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [6:5]),
    .fci(\u_DIV_SIGNED/al_00000256AA88ADA0 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88D0B0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA684000|u_DIV_SIGNED/al_00000256AA683230  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [10:9]),
    .fci(\u_DIV_SIGNED/al_00000256AA88AF00 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [10:9]),
    .fco(\u_DIV_SIGNED/al_00000256AA88D420 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA684110|u_DIV_SIGNED/al_00000256AA684DD0  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [26:25]),
    .fci(\u_DIV_SIGNED/al_00000256AA88CA80 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [26:25]),
    .fco(\u_DIV_SIGNED/al_00000256AA88B950 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA684440|u_DIV_SIGNED/al_00000256AA683EF0  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [22:21]),
    .fci(\u_DIV_SIGNED/al_00000256AA88CBE0 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [22:21]),
    .fco(\u_DIV_SIGNED/al_00000256AA88C5B0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA684550|u_DIV_SIGNED/al_00000256AA685CB0  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [4:3]),
    .fci(\u_DIV_SIGNED/al_00000256AA88AC40 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [4:3]),
    .fco(\u_DIV_SIGNED/al_00000256AA88B270 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA684990|u_DIV_SIGNED/al_00000256AA682DF0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [14:13]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [14:13]),
    .fci(\u_DIV_SIGNED/al_00000256AA88A8D0 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88C3A0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA684AA0|u_DIV_SIGNED/al_00000256AA683780  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [14:13]),
    .fci(\u_DIV_SIGNED/al_00000256AA88C240 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [14:13]),
    .fco(\u_DIV_SIGNED/al_00000256AA88C660 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA685100|u_DIV_SIGNED/al_00000256AA684EE0  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [20:19]),
    .fci(\u_DIV_SIGNED/al_00000256AA88CEA0 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [20:19]),
    .fco(\u_DIV_SIGNED/al_00000256AA88CBE0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660  (
    .a(2'b00),
    .b({\u_DIV_SIGNED/al_00000256AA0CF470 [0],1'b0}),
    .f({\u_DIV_SIGNED/al_00000256AA40B170 [0],open_n4384}),
    .fco(\u_DIV_SIGNED/al_00000256AA88C190 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA685760|u_DIV_SIGNED/al_00000256AA686420  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [2:1]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [2:1]),
    .fci(\u_DIV_SIGNED/al_00000256AA88C500 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88C450 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA685980|u_DIV_SIGNED/al_00000256AA682BD0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [10:9]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [10:9]),
    .fci(\u_DIV_SIGNED/al_00000256AA88A980 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88BCC0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA685A90|u_DIV_SIGNED/al_00000256AA685540  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [24:23]),
    .fci(\u_DIV_SIGNED/al_00000256AA88C5B0 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [24:23]),
    .fco(\u_DIV_SIGNED/al_00000256AA88CA80 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA685BA0|u_DIV_SIGNED/al_00000256AA683CD0  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [16:15]),
    .fci(\u_DIV_SIGNED/al_00000256AA88C660 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [16:15]),
    .fco(\u_DIV_SIGNED/al_00000256AA88BED0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA685ED0|u_DIV_SIGNED/al_00000256AA685210  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [30:29]),
    .fci(\u_DIV_SIGNED/al_00000256AA88B060 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [30:29]),
    .fco(\u_DIV_SIGNED/al_00000256AA88C710 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA686200_al_u429  (
    .a({open_n4503,1'b0}),
    .b({open_n4504,\u_DIV_SIGNED/al_00000256AA0CF470 [31]}),
    .fci(\u_DIV_SIGNED/al_00000256AA88C710 ),
    .f({open_n4523,\u_DIV_SIGNED/al_00000256AA40B170 [31]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA686640|u_DIV_SIGNED/al_00000256AA682AC0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [8:7]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [8:7]),
    .fci(\u_DIV_SIGNED/al_00000256AA88D0B0 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88A980 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA686860|u_DIV_SIGNED/al_00000256AA686970  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [12:11]),
    .fci(\u_DIV_SIGNED/al_00000256AA88D420 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [12:11]),
    .fco(\u_DIV_SIGNED/al_00000256AA88C240 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA685430|u_DIV_SIGNED/al_00000256AA684660"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA686A80|u_DIV_SIGNED/al_00000256AA685650  (
    .a(2'b00),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [28:27]),
    .fci(\u_DIV_SIGNED/al_00000256AA88B950 ),
    .f(\u_DIV_SIGNED/al_00000256AA40B170 [28:27]),
    .fco(\u_DIV_SIGNED/al_00000256AA88B060 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530  (
    .a({\u_DIV_SIGNED/al_00000256AA0D0BA0 [0],1'b1}),
    .b({\u_DIV_SIGNED/al_00000256AA0CF470 [0],1'b0}),
    .fco(\u_DIV_SIGNED/al_00000256AA88C500 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y14Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA686CA0|u_DIV_SIGNED/al_00000256AA689B60  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [56:55]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88DFD0 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88F680 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA686DB0|u_DIV_SIGNED/al_00000256AA6890C0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [26:25]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [26:25]),
    .fci(\u_DIV_SIGNED/al_00000256AA88BC10 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88BE20 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y14Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA686EC0|u_DIV_SIGNED/al_00000256AA687850  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [58:57]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88F680 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88E340 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y10Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6870E0|u_DIV_SIGNED/al_00000256AA688730  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [42:41]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88F890 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88E130 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y15Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6871F0|u_DIV_SIGNED/al_00000256AA686FD0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [62:61]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88F730 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88D630 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y9Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA687300|u_DIV_SIGNED/al_00000256AA688B70  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [38:37]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88F470 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88F3C0 ));
  EG_PHY_LSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256A66FB850_al_u414"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA687740_al_u416  (
    .a({\u_DIV_SIGNED/al_00000256AA0CF470 [9],\u_DIV_SIGNED/al_00000256AA0CF470 [7]}),
    .b({\u_DIV_SIGNED/al_00000256AA0CF470 [10],\u_DIV_SIGNED/al_00000256AA0CF470 [8]}),
    .c(2'b11),
    .d({\u_DIV_SIGNED/al_00000256AA0D0BA0 [9],\u_DIV_SIGNED/al_00000256AA0D0BA0 [7]}),
    .e({\u_DIV_SIGNED/al_00000256AA0D0BA0 [10],\u_DIV_SIGNED/al_00000256AA0D0BA0 [8]}),
    .fci(\u_DIV_SIGNED/al_00000256AA89AEC0 ),
    .f({\u_DIV_SIGNED/al_00000256AA400D60 [9],\u_DIV_SIGNED/al_00000256AA400D60 [7]}),
    .fco(\u_DIV_SIGNED/al_00000256AA899290 ),
    .fx({\u_DIV_SIGNED/al_00000256AA400D60 [10],\u_DIV_SIGNED/al_00000256AA400D60 [8]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA687C90|u_DIV_SIGNED/al_00000256AA683560  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [20:19]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [20:19]),
    .fci(\u_DIV_SIGNED/al_00000256AA88B480 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88BA00 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA687DA0|u_DIV_SIGNED/al_00000256AA6892E0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [22:21]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [22:21]),
    .fci(\u_DIV_SIGNED/al_00000256AA88BA00 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88BAB0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6880D0|u_DIV_SIGNED/al_00000256AA687EB0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [24:23]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [24:23]),
    .fci(\u_DIV_SIGNED/al_00000256AA88BAB0 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88BC10 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y8Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6881E0|u_DIV_SIGNED/al_00000256AA687520  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [34:33]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88DB00 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88EE40 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6882F0|u_DIV_SIGNED/al_00000256AA687FC0  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [28:27]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [28:27]),
    .fci(\u_DIV_SIGNED/al_00000256AA88BE20 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88C030 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y10Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA688400|u_DIV_SIGNED/al_00000256AA689C70  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [40:39]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88F3C0 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88F890 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y11Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA688840|u_DIV_SIGNED/al_00000256AA688C80  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [46:45]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88DE70 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88E1E0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA688A60|u_DIV_SIGNED/al_00000256AA688620  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [32:31]),
    .b({1'b0,\u_DIV_SIGNED/al_00000256AA0CF470 [31]}),
    .fci(\u_DIV_SIGNED/al_00000256AA88FC00 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88DB00 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y12Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA688EA0|u_DIV_SIGNED/al_00000256AA688D90  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [50:49]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88DF20 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88F520 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y11Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA688FB0|u_DIV_SIGNED/al_00000256AA688510  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [44:43]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88E130 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88DE70 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y12Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6891D0|u_DIV_SIGNED/al_00000256AA688950  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [48:47]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88E1E0 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88DF20 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y13Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA6893F0|u_DIV_SIGNED/al_00000256AA689D80  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [52:51]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88F520 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88F9F0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y13Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA689610|u_DIV_SIGNED/al_00000256AA689500  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [54:53]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88F9F0 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88DFD0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y9Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA689720|u_DIV_SIGNED/al_00000256AA689E90  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [36:35]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88EE40 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88F470 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA689940|u_DIV_SIGNED/al_00000256AA687B80  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [30:29]),
    .b(\u_DIV_SIGNED/al_00000256AA0CF470 [30:29]),
    .fci(\u_DIV_SIGNED/al_00000256AA88C030 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88FC00 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_SIGNED/al_00000256AA686B90|u_DIV_SIGNED/al_00000256AA675530"),
    //.R_POSITION("X0Y15Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_SIGNED/al_00000256AA689A50|u_DIV_SIGNED/al_00000256AA689830  (
    .a(\u_DIV_SIGNED/al_00000256AA0D0BA0 [60:59]),
    .b(2'b00),
    .fci(\u_DIV_SIGNED/al_00000256AA88E340 ),
    .fco(\u_DIV_SIGNED/al_00000256AA88F730 ));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE91F6C0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [30]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [30]));  // al_ip/div_unsigned_gate.v(2099)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE91F7D0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [6]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [7]));  // al_ip/div_unsigned_gate.v(2432)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE91F8E0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [5]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [6]));  // al_ip/div_unsigned_gate.v(2423)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE91F9F0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [7]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [8]));  // al_ip/div_unsigned_gate.v(2441)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE91FB00  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [8]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [9]));  // al_ip/div_unsigned_gate.v(2450)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE91FC10  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [20]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [21]));  // al_ip/div_unsigned_gate.v(2297)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE91FD20  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [22]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [23]));  // al_ip/div_unsigned_gate.v(2315)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE91FF40  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [13]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [14]));  // al_ip/div_unsigned_gate.v(2225)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE920050  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [16]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [16]));  // al_ip/div_unsigned_gate.v(1955)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE920160  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [19]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [19]));  // al_ip/div_unsigned_gate.v(1982)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE920270  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [27]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [27]));  // al_ip/div_unsigned_gate.v(2063)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE920490  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [21]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [22]));  // al_ip/div_unsigned_gate.v(2306)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE9205A0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [23]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [24]));  // al_ip/div_unsigned_gate.v(2324)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE9206B0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [24]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [25]));  // al_ip/div_unsigned_gate.v(2333)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE9207C0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [27]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [28]));  // al_ip/div_unsigned_gate.v(2360)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE9208D0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [28]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [29]));  // al_ip/div_unsigned_gate.v(2369)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE9209E0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [28]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [28]));  // al_ip/div_unsigned_gate.v(2072)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE920D10  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [1]),
    .sr(i_rstn),
    .q(div_unsigned_quo[1]));  // al_ip/div_unsigned_gate.v(2468)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE920E20  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [3]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [4]));  // al_ip/div_unsigned_gate.v(2405)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE920F30  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [26]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [26]));  // al_ip/div_unsigned_gate.v(2054)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE921040  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [14]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [15]));  // al_ip/div_unsigned_gate.v(2234)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE921150  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [29]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [30]));  // al_ip/div_unsigned_gate.v(2387)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE921260  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [0]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [1]));  // al_ip/div_unsigned_gate.v(2180)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE921370  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [26]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [27]));  // al_ip/div_unsigned_gate.v(2351)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE921480  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [30]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [31]));  // al_ip/div_unsigned_gate.v(2396)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE921590  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [15]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [15]));  // al_ip/div_unsigned_gate.v(1946)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE9216A0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [12]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [13]));  // al_ip/div_unsigned_gate.v(2216)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE9217B0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [15]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [16]));  // al_ip/div_unsigned_gate.v(2243)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE9218C0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [19]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [20]));  // al_ip/div_unsigned_gate.v(2288)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE921AE0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [4]),
    .sr(i_rstn),
    .q(div_unsigned_quo[4]));  // al_ip/div_unsigned_gate.v(2693)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE921BF0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [5]),
    .sr(i_rstn),
    .q(div_unsigned_quo[5]));  // al_ip/div_unsigned_gate.v(2702)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE921D00  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [20]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [20]));  // al_ip/div_unsigned_gate.v(2000)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE921E10  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [24]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [24]));  // al_ip/div_unsigned_gate.v(2036)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE921F20  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [10]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [11]));  // al_ip/div_unsigned_gate.v(2198)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE922030  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [17]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [17]));  // al_ip/div_unsigned_gate.v(1964)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE922140  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [2]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [3]));  // al_ip/div_unsigned_gate.v(2378)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE922250  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [4]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [5]));  // al_ip/div_unsigned_gate.v(2414)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE922360  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [1]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [2]));  // al_ip/div_unsigned_gate.v(2279)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE922470  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [11]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [12]));  // al_ip/div_unsigned_gate.v(2207)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE9227A0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [0]),
    .sr(i_rstn),
    .q(div_unsigned_quo[0]));  // al_ip/div_unsigned_gate.v(2459)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE9228B0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [25]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [25]));  // al_ip/div_unsigned_gate.v(2045)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE9229C0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [6]),
    .sr(i_rstn),
    .q(div_unsigned_quo[6]));  // al_ip/div_unsigned_gate.v(2711)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE922AD0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [23]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [23]));  // al_ip/div_unsigned_gate.v(2027)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE922BE0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [3]),
    .sr(i_rstn),
    .q(div_unsigned_quo[3]));  // al_ip/div_unsigned_gate.v(2666)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE922CF0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [7]),
    .sr(i_rstn),
    .q(div_unsigned_quo[7]));  // al_ip/div_unsigned_gate.v(2720)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE922E00  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [21]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [21]));  // al_ip/div_unsigned_gate.v(2009)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE922F10  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [16]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [17]));  // al_ip/div_unsigned_gate.v(2252)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE923020  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [17]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [18]));  // al_ip/div_unsigned_gate.v(2261)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE923130  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [31]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [31]));  // al_ip/div_unsigned_gate.v(2108)
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y16Z0"),
    .ALUTYPE("A_LE_B"),
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"),
    .REG0_REGSET("RESET"),
    .REG0_SD("F"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE923240_al_u430  (
    .a({open_n5224,1'b0}),
    .b({open_n5225,1'b1}),
    .clk(i_clk),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A26D40 ),
    .sr(div_unsigned_start),
    .f({open_n5242,\u_DIV_UNSIGNED/al_00000286E5A5D8C0 }),
    .q({open_n5246,\u_DIV_UNSIGNED/al_00000286E57DBF10 [0]}));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE923350  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [25]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [26]));  // al_ip/div_unsigned_gate.v(2342)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE923460  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [29]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [29]));  // al_ip/div_unsigned_gate.v(2081)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE923570  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [2]),
    .sr(i_rstn),
    .q(div_unsigned_quo[2]));  // al_ip/div_unsigned_gate.v(2567)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE923680  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [22]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [22]));  // al_ip/div_unsigned_gate.v(2018)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE923790  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [9]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [10]));  // al_ip/div_unsigned_gate.v(2189)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286DE9238A0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [18]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DBF10 [19]));  // al_ip/div_unsigned_gate.v(2270)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286DE9239B0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [18]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [18]));  // al_ip/div_unsigned_gate.v(1973)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE923AC0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [2]),
    .sr(i_rstn),
    .q(div_unsigned_rem[2]));  // al_ip/div_unsigned_gate.v(2855)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE923CE0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [12]),
    .sr(i_rstn),
    .q(div_unsigned_quo[12]));  // al_ip/div_unsigned_gate.v(2495)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE923DF0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [14]),
    .sr(i_rstn),
    .q(div_unsigned_quo[14]));  // al_ip/div_unsigned_gate.v(2513)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE923F00  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [16]),
    .sr(i_rstn),
    .q(div_unsigned_quo[16]));  // al_ip/div_unsigned_gate.v(2531)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE924230  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [28]),
    .sr(i_rstn),
    .q(div_unsigned_quo[28]));  // al_ip/div_unsigned_gate.v(2648)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE924450  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [0]),
    .sr(i_rstn),
    .q(div_unsigned_rem[0]));  // al_ip/div_unsigned_gate.v(2747)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE924560  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [7]),
    .sr(i_rstn),
    .q(div_unsigned_rem[7]));  // al_ip/div_unsigned_gate.v(3008)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE924890  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [13]),
    .sr(i_rstn),
    .q(div_unsigned_quo[13]));  // al_ip/div_unsigned_gate.v(2504)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE924DE0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [15]),
    .sr(i_rstn),
    .q(div_unsigned_quo[15]));  // al_ip/div_unsigned_gate.v(2522)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE925000  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [19]),
    .sr(i_rstn),
    .q(div_unsigned_quo[19]));  // al_ip/div_unsigned_gate.v(2558)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE925110  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [23]),
    .sr(i_rstn),
    .q(div_unsigned_quo[23]));  // al_ip/div_unsigned_gate.v(2603)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE925220  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [24]),
    .sr(i_rstn),
    .q(div_unsigned_quo[24]));  // al_ip/div_unsigned_gate.v(2612)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE925330  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [27]),
    .sr(i_rstn),
    .q(div_unsigned_quo[27]));  // al_ip/div_unsigned_gate.v(2639)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE925550  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [8]),
    .sr(i_rstn),
    .q(div_unsigned_quo[8]));  // al_ip/div_unsigned_gate.v(2729)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE925660  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [9]),
    .sr(i_rstn),
    .q(div_unsigned_quo[9]));  // al_ip/div_unsigned_gate.v(2738)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE925770  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [17]),
    .sr(i_rstn),
    .q(div_unsigned_quo[17]));  // al_ip/div_unsigned_gate.v(2540)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE925880  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [30]),
    .sr(i_rstn),
    .q(div_unsigned_quo[30]));  // al_ip/div_unsigned_gate.v(2675)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE925AA0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [31]),
    .sr(i_rstn),
    .q(div_unsigned_quo[31]));  // al_ip/div_unsigned_gate.v(2684)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE925BB0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [25]),
    .sr(i_rstn),
    .q(div_unsigned_quo[25]));  // al_ip/div_unsigned_gate.v(2621)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE925CC0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [22]),
    .sr(i_rstn),
    .q(div_unsigned_quo[22]));  // al_ip/div_unsigned_gate.v(2594)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE926430  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [26]),
    .sr(i_rstn),
    .q(div_unsigned_quo[26]));  // al_ip/div_unsigned_gate.v(2630)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE926540  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [18]),
    .sr(i_rstn),
    .q(div_unsigned_quo[18]));  // al_ip/div_unsigned_gate.v(2549)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE926650  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [20]),
    .sr(i_rstn),
    .q(div_unsigned_quo[20]));  // al_ip/div_unsigned_gate.v(2576)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE926870  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [3]),
    .sr(i_rstn),
    .q(div_unsigned_rem[3]));  // al_ip/div_unsigned_gate.v(2954)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE926980  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [4]),
    .sr(i_rstn),
    .q(div_unsigned_rem[4]));  // al_ip/div_unsigned_gate.v(2981)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE926A90  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [5]),
    .sr(i_rstn),
    .q(div_unsigned_rem[5]));  // al_ip/div_unsigned_gate.v(2990)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE926CB0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [6]),
    .sr(i_rstn),
    .q(div_unsigned_rem[6]));  // al_ip/div_unsigned_gate.v(2999)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE926ED0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [11]),
    .sr(i_rstn),
    .q(div_unsigned_quo[11]));  // al_ip/div_unsigned_gate.v(2486)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE926FE0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [21]),
    .sr(i_rstn),
    .q(div_unsigned_quo[21]));  // al_ip/div_unsigned_gate.v(2585)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE9270F0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [29]),
    .sr(i_rstn),
    .q(div_unsigned_quo[29]));  // al_ip/div_unsigned_gate.v(2657)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE927200  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DBF10 [10]),
    .sr(i_rstn),
    .q(div_unsigned_quo[10]));  // al_ip/div_unsigned_gate.v(2477)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DE927420  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [1]),
    .sr(i_rstn),
    .q(div_unsigned_rem[1]));  // al_ip/div_unsigned_gate.v(2756)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA92230  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [11]),
    .sr(i_rstn),
    .q(div_unsigned_rem[11]));  // al_ip/div_unsigned_gate.v(2774)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA92340  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [25]),
    .sr(i_rstn),
    .q(div_unsigned_rem[25]));  // al_ip/div_unsigned_gate.v(2909)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA92450  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E04A0 [4]),
    .sr(i_rstn),
    .q(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [4]));  // al_ip/div_unsigned_gate.v(3071)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA92AB0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [9]),
    .sr(i_rstn),
    .q(div_unsigned_rem[9]));  // al_ip/div_unsigned_gate.v(3026)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA92BC0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [20]),
    .sr(i_rstn),
    .q(div_unsigned_rem[20]));  // al_ip/div_unsigned_gate.v(2864)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA93220  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [18]),
    .sr(i_rstn),
    .q(div_unsigned_rem[18]));  // al_ip/div_unsigned_gate.v(2837)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA93330  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [23]),
    .sr(i_rstn),
    .q(div_unsigned_rem[23]));  // al_ip/div_unsigned_gate.v(2891)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA93550  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [17]),
    .sr(i_rstn),
    .q(div_unsigned_rem[17]));  // al_ip/div_unsigned_gate.v(2828)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA93660  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [29]),
    .sr(i_rstn),
    .q(div_unsigned_rem[29]));  // al_ip/div_unsigned_gate.v(2945)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA93880  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [8]),
    .sr(i_rstn),
    .q(div_unsigned_rem[8]));  // al_ip/div_unsigned_gate.v(3017)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA93AA0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E04A0 [2]),
    .sr(i_rstn),
    .q(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [2]));  // al_ip/div_unsigned_gate.v(3053)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA93DD0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [16]),
    .sr(i_rstn),
    .q(div_unsigned_rem[16]));  // al_ip/div_unsigned_gate.v(2819)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA94320  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [19]),
    .sr(i_rstn),
    .q(div_unsigned_rem[19]));  // al_ip/div_unsigned_gate.v(2846)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA94540  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [13]),
    .sr(i_rstn),
    .q(div_unsigned_rem[13]));  // al_ip/div_unsigned_gate.v(2792)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA94870  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [10]),
    .sr(i_rstn),
    .q(div_unsigned_rem[10]));  // al_ip/div_unsigned_gate.v(2765)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA94980  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [12]),
    .sr(i_rstn),
    .q(div_unsigned_rem[12]));  // al_ip/div_unsigned_gate.v(2783)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA94A90  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [15]),
    .sr(i_rstn),
    .q(div_unsigned_rem[15]));  // al_ip/div_unsigned_gate.v(2810)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA94CB0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [14]),
    .sr(i_rstn),
    .q(div_unsigned_rem[14]));  // al_ip/div_unsigned_gate.v(2801)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA94DC0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [21]),
    .sr(i_rstn),
    .q(div_unsigned_rem[21]));  // al_ip/div_unsigned_gate.v(2873)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA94ED0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [22]),
    .sr(i_rstn),
    .q(div_unsigned_rem[22]));  // al_ip/div_unsigned_gate.v(2882)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA94FE0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [26]),
    .sr(i_rstn),
    .q(div_unsigned_rem[26]));  // al_ip/div_unsigned_gate.v(2918)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA950F0  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [28]),
    .sr(i_rstn),
    .q(div_unsigned_rem[28]));  // al_ip/div_unsigned_gate.v(2936)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA95200  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [30]),
    .sr(i_rstn),
    .q(div_unsigned_rem[30]));  // al_ip/div_unsigned_gate.v(2963)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA95310  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E04A0 [0]),
    .sr(i_rstn),
    .q(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [0]));  // al_ip/div_unsigned_gate.v(3035)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA95420  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E04A0 [1]),
    .sr(i_rstn),
    .q(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [1]));  // al_ip/div_unsigned_gate.v(3044)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA95530  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E04A0 [3]),
    .sr(i_rstn),
    .q(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [3]));  // al_ip/div_unsigned_gate.v(3062)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA95640  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E04A0 [5]),
    .sr(i_rstn),
    .q(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [5]));  // al_ip/div_unsigned_gate.v(3080)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA95750  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [24]),
    .sr(i_rstn),
    .q(div_unsigned_rem[24]));  // al_ip/div_unsigned_gate.v(2900)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA95860  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [31]),
    .sr(i_rstn),
    .q(div_unsigned_rem[31]));  // al_ip/div_unsigned_gate.v(2972)
  AL_MAP_SEQ #(
    .CEMUX("CE"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286DEA95970  (
    .ce(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [27]),
    .sr(i_rstn),
    .q(div_unsigned_rem[27]));  // al_ip/div_unsigned_gate.v(2927)
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443B780|u_DIV_UNSIGNED/al_00000286E4444F70  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [10:9]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [10:9]),
    .fci(\u_DIV_UNSIGNED/al_00000286E44833F0 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [10:9]),
    .fco(\u_DIV_UNSIGNED/al_00000286E4481B30 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443B9A0|u_DIV_UNSIGNED/al_00000286E443C990  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [12:11]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [12:11]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4481B30 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [12:11]),
    .fco(\u_DIV_UNSIGNED/al_00000286E44810E0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443BAB0|u_DIV_UNSIGNED/al_00000286E443E970  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [14:13]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [14:13]),
    .fci(\u_DIV_UNSIGNED/al_00000286E44810E0 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [14:13]),
    .fco(\u_DIV_UNSIGNED/al_00000286E44808A0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443BCD0|u_DIV_UNSIGNED/al_00000286E443CFF0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [18:17]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [18:17]),
    .fci(\u_DIV_UNSIGNED/al_00000286E44819D0 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [18:17]),
    .fco(\u_DIV_UNSIGNED/al_00000286E4480480 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443C110|u_DIV_UNSIGNED/al_00000286E443C000  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [2:1]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [2:1]),
    .fci(\u_DIV_UNSIGNED/al_00000286E447F350 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [2:1]),
    .fco(\u_DIV_UNSIGNED/al_00000286E44805E0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("SUB_CARRY"),
    .INIT_LUT0(16'b0000000000000101),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0  (
    .a({\u_DIV_UNSIGNED/al_00000286E57DC290 [0],1'b0}),
    .b({\u_DIV_UNSIGNED/al_00000286E57DE2F0 [0],1'b0}),
    .f({\u_DIV_UNSIGNED/al_00000286E57E1690 [0],open_n5391}),
    .fco(\u_DIV_UNSIGNED/al_00000286E447F350 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443C440|u_DIV_UNSIGNED/al_00000286E443C330  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [26:25]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [26:25]),
    .fci(\u_DIV_UNSIGNED/al_00000286E447FF00 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [26:25]),
    .fco(\u_DIV_UNSIGNED/al_00000286E4480530 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443CAA0|u_DIV_UNSIGNED/al_00000286E443BBC0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [16:15]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [16:15]),
    .fci(\u_DIV_UNSIGNED/al_00000286E44808A0 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [16:15]),
    .fco(\u_DIV_UNSIGNED/al_00000286E44819D0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443D210|u_DIV_UNSIGNED/al_00000286E443C550  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [28:27]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [28:27]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4480530 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [28:27]),
    .fco(\u_DIV_UNSIGNED/al_00000286E44812F0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443DCB0|u_DIV_UNSIGNED/al_00000286E443D320  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [20:19]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [20:19]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4480480 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [20:19]),
    .fco(\u_DIV_UNSIGNED/al_00000286E447FE50 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443DED0|u_DIV_UNSIGNED/al_00000286E443D100  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [24:23]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [24:23]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4480CC0 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [24:23]),
    .fco(\u_DIV_UNSIGNED/al_00000286E447FF00 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443DFE0|u_DIV_UNSIGNED/al_00000286E443D430  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [30:29]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [30:29]),
    .fci(\u_DIV_UNSIGNED/al_00000286E44812F0 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [30:29]),
    .fco(\u_DIV_UNSIGNED/al_00000286E4480B60 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443E0F0_al_u431  (
    .a({open_n5528,\u_DIV_UNSIGNED/al_00000286E57DC290 [31]}),
    .b({open_n5529,\u_DIV_UNSIGNED/al_00000286E57DE2F0 [31]}),
    .fci(\u_DIV_UNSIGNED/al_00000286E4480B60 ),
    .f({open_n5548,\u_DIV_UNSIGNED/al_00000286E57E1690 [31]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443E200|u_DIV_UNSIGNED/al_00000286E443D540  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [4:3]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [4:3]),
    .fci(\u_DIV_UNSIGNED/al_00000286E44805E0 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [4:3]),
    .fco(\u_DIV_UNSIGNED/al_00000286E44815B0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443E530|u_DIV_UNSIGNED/al_00000286E443E310  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [6:5]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [6:5]),
    .fci(\u_DIV_UNSIGNED/al_00000286E44815B0 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [6:5]),
    .fco(\u_DIV_UNSIGNED/al_00000286E4481710 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443EA80|u_DIV_UNSIGNED/al_00000286E443DDC0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [22:21]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [22:21]),
    .fci(\u_DIV_UNSIGNED/al_00000286E447FE50 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [22:21]),
    .fco(\u_DIV_UNSIGNED/al_00000286E4480CC0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443ECA0|u_DIV_UNSIGNED/al_00000286E44424F0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [8:7]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [8:7]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A24FB0 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A24820 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y3Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443EEC0|u_DIV_UNSIGNED/al_00000286E44412E0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [12:11]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [12:11]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A25740 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A23F30 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443F300|u_DIV_UNSIGNED/al_00000286E44411D0"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("ADD_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443F300|u_DIV_UNSIGNED/al_00000286E44411D0  (
    .a({\u_DIV_UNSIGNED/al_00000286E57DB3B0 [0],1'b0}),
    .b(2'b10),
    .f({\u_DIV_UNSIGNED/al_00000286E57E03C0 [0],open_n5687}),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A24560 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y3Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443F630|u_DIV_UNSIGNED/al_00000286E443EFD0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [14:13]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [14:13]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A23F30 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A23FE0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y4Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443FA70|u_DIV_UNSIGNED/al_00000286E443F960  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [18:17]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [18:17]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A25060 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A258A0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443F300|u_DIV_UNSIGNED/al_00000286E44411D0"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443FC90|u_DIV_UNSIGNED/al_00000286E4442D70  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [4:3]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A24E50 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E03C0 [4:3]),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A24A30 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y5Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E443FFC0|u_DIV_UNSIGNED/al_00000286E443FEB0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [22:21]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [22:21]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A25950 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A25ED0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y6Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44401E0|u_DIV_UNSIGNED/al_00000286E44400D0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [24:23]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [24:23]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A25ED0 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A25A00 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y6Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44402F0|u_DIV_UNSIGNED/al_00000286E4441500  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [26:25]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [26:25]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A25A00 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A25C10 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y7Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4440620|u_DIV_UNSIGNED/al_00000286E4440510  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [30:29]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [30:29]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A25F80 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A260E0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4440840|u_DIV_UNSIGNED/al_00000286E443FDA0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [2:1]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [2:1]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A25530 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A23D20 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y8Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4440A60|u_DIV_UNSIGNED/al_00000286E4440950  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [34:33]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A27BB0 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A28810 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y7Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4440D90|u_DIV_UNSIGNED/al_00000286E4440400  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [28:27]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [28:27]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A25C10 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A25F80 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y8Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4440FB0|u_DIV_UNSIGNED/al_00000286E4440730  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [32:31]),
    .b({1'b0,\u_DIV_UNSIGNED/al_00000286E57DC290 [31]}),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A260E0 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A27BB0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y9Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44410C0|u_DIV_UNSIGNED/al_00000286E4440EA0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [36:35]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A28810 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A26A80 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y0Z0"),
    .ALUTYPE("A_LE_B_CARRY"),
    .INIT_LUT0(16'b0000000000001010),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600  (
    .a({\u_DIV_UNSIGNED/al_00000286E57DE2F0 [0],1'b1}),
    .b({\u_DIV_UNSIGNED/al_00000286E57DC290 [0],1'b0}),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A25530 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4441830|u_DIV_UNSIGNED/al_00000286E4442930  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [6:5]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [6:5]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A25690 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A24FB0 ));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286E4441A50  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .sr(i_rstn),
    .q(div_unsigned_finish));  // al_ip/div_unsigned_gate.v(854)
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443F300|u_DIV_UNSIGNED/al_00000286E44411D0"),
    //.R_POSITION("X0Y0Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4441E90|u_DIV_UNSIGNED/al_00000286E4441D80  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [2:1]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A24560 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E03C0 [2:1]),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A24E50 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443F300|u_DIV_UNSIGNED/al_00000286E44411D0"),
    //.R_POSITION("X0Y1Z1"),
    .ALUTYPE("ADD"),
    .INIT_LUT0(16'b0110011001101010),
    .INIT_LUT1(16'b0110011001101010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4441FA0_al_u432  (
    .a({open_n6050,\u_DIV_UNSIGNED/al_00000286E57DB3B0 [5]}),
    .b({open_n6051,1'b0}),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A24A30 ),
    .f({open_n6070,\u_DIV_UNSIGNED/al_00000286E57E03C0 [5]}));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y2Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44420B0|u_DIV_UNSIGNED/al_00000286E443EDB0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [10:9]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [10:9]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A24820 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A25740 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y4Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44422D0|u_DIV_UNSIGNED/al_00000286E443F850  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [16:15]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [16:15]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A23FE0 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A25060 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y5Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44423E0|u_DIV_UNSIGNED/al_00000286E443FB80  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [20:19]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [20:19]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A258A0 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A25950 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y1Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4442F90|u_DIV_UNSIGNED/al_00000286E4442820  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [4:3]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DC290 [4:3]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A23D20 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A25690 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y14Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44432C0|u_DIV_UNSIGNED/al_00000286E4446180  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [58:57]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A272C0 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A28E40 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y11Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44433D0|u_DIV_UNSIGNED/al_00000286E4443700  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [46:45]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A27C60 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A27370 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y13Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44435F0|u_DIV_UNSIGNED/al_00000286E4446070  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [52:51]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A28B80 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A26BE0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y9Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4443A30|u_DIV_UNSIGNED/al_00000286E4441720  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [38:37]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A26A80 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A26F50 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y10Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4443C50|u_DIV_UNSIGNED/al_00000286E44457F0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [40:39]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A26F50 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A276E0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y11Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44443C0|u_DIV_UNSIGNED/al_00000286E4445F60  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [44:43]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A270B0 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A27C60 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y15Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44445E0|u_DIV_UNSIGNED/al_00000286E44455D0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [60:59]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A28E40 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A27160 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y10Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44454C0|u_DIV_UNSIGNED/al_00000286E4444800  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [42:41]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A276E0 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A270B0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y12Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E44464B0|u_DIV_UNSIGNED/al_00000286E44453B0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [48:47]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A27370 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A27210 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y12Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4446C20|u_DIV_UNSIGNED/al_00000286E44434E0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [50:49]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A27210 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A28B80 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y15Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4446E40|u_DIV_UNSIGNED/al_00000286E4443810  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [62:61]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A27160 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A26D40 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y13Z1"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4447060|u_DIV_UNSIGNED/al_00000286E44444D0  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [54:53]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A26BE0 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A27B00 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E443C220|u_DIV_UNSIGNED/al_00000286E44446F0"),
    //.R_POSITION("X0Y2Z0"),
    .ALUTYPE("SUB"),
    .INIT_LUT0(16'b1001100110011010),
    .INIT_LUT1(16'b1001100110011010),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4447280|u_DIV_UNSIGNED/al_00000286E4447170  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DC290 [8:7]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [8:7]),
    .fci(\u_DIV_UNSIGNED/al_00000286E4481710 ),
    .f(\u_DIV_UNSIGNED/al_00000286E57E1690 [8:7]),
    .fco(\u_DIV_UNSIGNED/al_00000286E44833F0 ));
  EG_PHY_MSLICE #(
    //.MACRO("u_DIV_UNSIGNED/al_00000286E44413F0|u_DIV_UNSIGNED/al_00000286E4442600"),
    //.R_POSITION("X0Y14Z0"),
    .ALUTYPE("A_LE_B"),
    .INIT_LUT0(16'b1001100110011100),
    .INIT_LUT1(16'b1001100110011100),
    .MODE("RIPPLE"))
    \u_DIV_UNSIGNED/al_00000286E4447390|u_DIV_UNSIGNED/al_00000286E4443B40  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [56:55]),
    .b(2'b00),
    .fci(\u_DIV_UNSIGNED/al_00000286E4A27B00 ),
    .fco(\u_DIV_UNSIGNED/al_00000286E4A272C0 ));
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC86D0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [55]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [55]));  // al_ip/div_unsigned_gate.v(1775)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC87E0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [5]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [5]));  // al_ip/div_unsigned_gate.v(2126)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC8B10  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [57]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [57]));  // al_ip/div_unsigned_gate.v(1793)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC8D30  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [3]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [3]));  // al_ip/div_unsigned_gate.v(2090)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC8E40  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [7]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [7]));  // al_ip/div_unsigned_gate.v(2144)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC8F50  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [8]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [8]));  // al_ip/div_unsigned_gate.v(2153)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC94A0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [4]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [4]));  // al_ip/div_unsigned_gate.v(2117)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC95B0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [2]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [2]));  // al_ip/div_unsigned_gate.v(1991)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC96C0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [6]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [6]));  // al_ip/div_unsigned_gate.v(2135)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC97D0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [9]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [9]));  // al_ip/div_unsigned_gate.v(2162)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC99F0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [56]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [56]));  // al_ip/div_unsigned_gate.v(1784)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC9B00  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [10]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [10]));  // al_ip/div_unsigned_gate.v(1901)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC9E30  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [11]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [11]));  // al_ip/div_unsigned_gate.v(1910)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BC9F40  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [12]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [12]));  // al_ip/div_unsigned_gate.v(1919)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BCA050  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [13]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [13]));  // al_ip/div_unsigned_gate.v(1928)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BCA270  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [14]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [14]));  // al_ip/div_unsigned_gate.v(1937)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BCB7B0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [58]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [58]));  // al_ip/div_unsigned_gate.v(1802)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BCB8C0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [59]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [59]));  // al_ip/div_unsigned_gate.v(1811)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BCB9D0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [60]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [60]));  // al_ip/div_unsigned_gate.v(1829)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BCBAE0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [61]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [61]));  // al_ip/div_unsigned_gate.v(1838)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("INV"))
    \u_DIV_UNSIGNED/al_00000286E4BCBBF0  (
    .clk(i_clk),
    .d(n34[31]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [62]));  // al_ip/div_unsigned_gate.v(1847)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BCBD00  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [0]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [0]));  // al_ip/div_unsigned_gate.v(1883)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BCC580  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57E4870 [1]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DC290 [1]));  // al_ip/div_unsigned_gate.v(1892)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDD8B0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [47]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [47]));  // al_ip/div_unsigned_gate.v(1694)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDD9C0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [20]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [19]));  // al_ip/div_unsigned_gate.v(1415)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDDAD0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [52]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [52]));  // al_ip/div_unsigned_gate.v(1748)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDDBE0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [53]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [53]));  // al_ip/div_unsigned_gate.v(1757)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDDE00  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [54]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [54]));  // al_ip/div_unsigned_gate.v(1766)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDDF10  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [28]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [27]));  // al_ip/div_unsigned_gate.v(1496)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDE020  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [38]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [38]));  // al_ip/div_unsigned_gate.v(1604)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDE130  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [9]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [8]));  // al_ip/div_unsigned_gate.v(1865)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDE460  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [12]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [11]));  // al_ip/div_unsigned_gate.v(1343)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDE570  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [21]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [20]));  // al_ip/div_unsigned_gate.v(1433)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDE790  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [48]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [48]));  // al_ip/div_unsigned_gate.v(1703)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDE8A0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [2]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [1]));  // al_ip/div_unsigned_gate.v(1325)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDE9B0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [4]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [3]));  // al_ip/div_unsigned_gate.v(1523)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDEAC0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [7]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [6]));  // al_ip/div_unsigned_gate.v(1820)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDEBD0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [8]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [7]));  // al_ip/div_unsigned_gate.v(1856)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDECE0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [11]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [10]));  // al_ip/div_unsigned_gate.v(1334)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDEDF0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [35]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [35]));  // al_ip/div_unsigned_gate.v(1577)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDEF00  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [27]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [26]));  // al_ip/div_unsigned_gate.v(1487)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDF010  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [34]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [34]));  // al_ip/div_unsigned_gate.v(1568)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDF120  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [32]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [32]));  // al_ip/div_unsigned_gate.v(1550)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDF230  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [39]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [39]));  // al_ip/div_unsigned_gate.v(1613)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDF340  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [24]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [23]));  // al_ip/div_unsigned_gate.v(1460)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDF450  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [45]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [45]));  // al_ip/div_unsigned_gate.v(1676)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDF560  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [49]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [49]));  // al_ip/div_unsigned_gate.v(1712)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDF670  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [36]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [36]));  // al_ip/div_unsigned_gate.v(1586)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDF780  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [50]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [50]));  // al_ip/div_unsigned_gate.v(1730)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BDF890  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [51]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [51]));  // al_ip/div_unsigned_gate.v(1739)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDF9A0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [22]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [21]));  // al_ip/div_unsigned_gate.v(1442)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDFAB0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [17]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [16]));  // al_ip/div_unsigned_gate.v(1388)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDFCD0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [1]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [0]));  // al_ip/div_unsigned_gate.v(1316)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDFDE0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [6]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [5]));  // al_ip/div_unsigned_gate.v(1721)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BDFEF0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [5]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [4]));  // al_ip/div_unsigned_gate.v(1622)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE0110  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [30]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [29]));  // al_ip/div_unsigned_gate.v(1514)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE0220  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [25]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [24]));  // al_ip/div_unsigned_gate.v(1469)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE0330  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [15]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [14]));  // al_ip/div_unsigned_gate.v(1370)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE0440  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [26]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [25]));  // al_ip/div_unsigned_gate.v(1478)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE0550  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [31]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [30]));  // al_ip/div_unsigned_gate.v(1532)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BE0660  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [37]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [37]));  // al_ip/div_unsigned_gate.v(1595)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE0770  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [3]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [2]));  // al_ip/div_unsigned_gate.v(1424)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE0990  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [14]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [13]));  // al_ip/div_unsigned_gate.v(1361)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE0AA0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [29]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [28]));  // al_ip/div_unsigned_gate.v(1505)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE0BB0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [10]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [9]));  // al_ip/div_unsigned_gate.v(1874)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BE0CC0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [33]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [33]));  // al_ip/div_unsigned_gate.v(1559)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BE0DD0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [40]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [40]));  // al_ip/div_unsigned_gate.v(1631)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BE0EE0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [42]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [42]));  // al_ip/div_unsigned_gate.v(1649)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE0FF0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [19]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [18]));  // al_ip/div_unsigned_gate.v(1406)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BE1100  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [43]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [43]));  // al_ip/div_unsigned_gate.v(1658)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE1210  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [23]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [22]));  // al_ip/div_unsigned_gate.v(1451)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BE1320  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [44]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [44]));  // al_ip/div_unsigned_gate.v(1667)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BE1430  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [46]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [46]));  // al_ip/div_unsigned_gate.v(1685)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE1540  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [16]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [15]));  // al_ip/div_unsigned_gate.v(1379)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BE1650  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [41]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [41]));  // al_ip/div_unsigned_gate.v(1640)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE1760  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [13]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [12]));  // al_ip/div_unsigned_gate.v(1352)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("SYNC"),
    .SRMUX("SR"))
    \u_DIV_UNSIGNED/al_00000286E4BE1A90  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [18]),
    .sr(div_unsigned_start),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [17]));  // al_ip/div_unsigned_gate.v(1397)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("0"))
    \u_DIV_UNSIGNED/al_00000286E4BE1BA0  (
    .clk(i_clk),
    .d(\u_DIV_UNSIGNED/al_00000286E57DEE50 [31]),
    .q(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [31]));  // al_ip/div_unsigned_gate.v(1541)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E578F490  (
    .a(n35[16]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [16]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [16]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [16]));  // al_ip/div_unsigned_gate.v(441)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E578F5A0  (
    .a(n35[19]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [19]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [19]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [19]));  // al_ip/div_unsigned_gate.v(479)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E578F6B0  (
    .a(n35[2]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [2]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [2]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [2]));  // al_ip/div_unsigned_gate.v(489)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E578F7C0  (
    .a(n34[6]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [38]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [37]));  // al_ip/div_unsigned_gate.v(667)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E578F8D0  (
    .a(n34[18]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [50]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [49]));  // al_ip/div_unsigned_gate.v(241)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E578F9E0  (
    .a(n35[21]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [21]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [21]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [21]));  // al_ip/div_unsigned_gate.v(509)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E578FAF0  (
    .a(n34[9]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [41]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [40]));  // al_ip/div_unsigned_gate.v(802)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E578FC00  (
    .a(n34[10]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [42]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [41]));  // al_ip/div_unsigned_gate.v(177)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E578FD10  (
    .a(n34[22]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [54]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [53]));  // al_ip/div_unsigned_gate.v(281)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E578FE20  (
    .a(n35[3]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [3]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [3]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [3]));  // al_ip/div_unsigned_gate.v(607)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E578FF30  (
    .a(n35[4]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [4]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [4]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [4]));  // al_ip/div_unsigned_gate.v(637)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5790040  (
    .a(n34[14]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [46]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [45]));  // al_ip/div_unsigned_gate.v(209)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5790150  (
    .a(n35[5]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [5]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [5]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [5]));  // al_ip/div_unsigned_gate.v(647)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5790260  (
    .a(n35[20]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [20]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [20]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [20]));  // al_ip/div_unsigned_gate.v(499)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5790370  (
    .a(n34[16]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [48]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [47]));  // al_ip/div_unsigned_gate.v(225)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5790480  (
    .a(n34[20]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [52]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [51]));  // al_ip/div_unsigned_gate.v(265)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5790590  (
    .a(n34[24]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [56]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [55]));  // al_ip/div_unsigned_gate.v(297)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E57906A0  (
    .a(n34[29]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [61]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [60]));  // al_ip/div_unsigned_gate.v(337)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E57907B0  (
    .a(n34[30]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [62]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [61]));  // al_ip/div_unsigned_gate.v(353)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E57908C0  (
    .a(n34[7]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [39]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [38]));  // al_ip/div_unsigned_gate.v(768)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E57909D0  (
    .a(n35[11]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [11]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [11]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [11]));  // al_ip/div_unsigned_gate.v(391)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5790AE0  (
    .a(n34[21]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [53]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [52]));  // al_ip/div_unsigned_gate.v(273)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5790BF0  (
    .a(n35[17]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [17]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [17]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [17]));  // al_ip/div_unsigned_gate.v(459)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5790D00  (
    .a(n35[26]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [26]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [26]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [26]));  // al_ip/div_unsigned_gate.v(567)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5790E10  (
    .a(n34[15]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [47]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [46]));  // al_ip/div_unsigned_gate.v(217)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5790F20  (
    .a(n35[28]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [28]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [28]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [28]));  // al_ip/div_unsigned_gate.v(587)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791030  (
    .a(n35[7]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [7]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [7]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [7]));  // al_ip/div_unsigned_gate.v(675)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5791140  (
    .a(n34[3]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [35]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [34]));  // al_ip/div_unsigned_gate.v(345)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5791250  (
    .a(n34[2]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [34]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [33]));  // al_ip/div_unsigned_gate.v(257)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791360  (
    .a(n35[1]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [1]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [1]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [1]));  // al_ip/div_unsigned_gate.v(371)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5791470  (
    .a(n34[4]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [36]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [35]));  // al_ip/div_unsigned_gate.v(451)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5791580  (
    .a(n34[17]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [49]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [48]));  // al_ip/div_unsigned_gate.v(233)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791690  (
    .a(n35[22]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [22]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [22]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [22]));  // al_ip/div_unsigned_gate.v(519)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E57917A0  (
    .a(n35[23]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [23]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [23]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [23]));  // al_ip/div_unsigned_gate.v(529)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E57918B0  (
    .a(n34[5]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [37]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [36]));  // al_ip/div_unsigned_gate.v(559)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E57919C0  (
    .a(n35[24]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [24]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [24]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [24]));  // al_ip/div_unsigned_gate.v(539)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791AD0  (
    .a(n35[30]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [30]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [30]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [30]));  // al_ip/div_unsigned_gate.v(617)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791BE0  (
    .a(n35[10]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [10]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [10]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [10]));  // al_ip/div_unsigned_gate.v(381)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791CF0  (
    .a(n35[31]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [31]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [31]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [31]));  // al_ip/div_unsigned_gate.v(627)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791E00  (
    .a(n35[8]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [8]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [8]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [8]));  // al_ip/div_unsigned_gate.v(685)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5791F10  (
    .a(n35[18]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [18]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [18]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [18]));  // al_ip/div_unsigned_gate.v(469)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792020  (
    .a(n34[26]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [58]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [57]));  // al_ip/div_unsigned_gate.v(313)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792130  (
    .a(n34[27]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [59]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [58]));  // al_ip/div_unsigned_gate.v(321)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792240  (
    .a(n34[12]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [44]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [43]));  // al_ip/div_unsigned_gate.v(193)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792350  (
    .a(n34[25]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [57]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [56]));  // al_ip/div_unsigned_gate.v(305)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5792460  (
    .a(n35[14]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [14]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [14]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [14]));  // al_ip/div_unsigned_gate.v(421)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5792570  (
    .a(n35[25]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [25]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [25]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [25]));  // al_ip/div_unsigned_gate.v(549)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5792680  (
    .a(n35[27]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [27]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [27]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [27]));  // al_ip/div_unsigned_gate.v(577)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5792790  (
    .a(n35[9]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [9]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [9]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [9]));  // al_ip/div_unsigned_gate.v(695)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E57928A0  (
    .a(n35[6]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [6]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [6]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [6]));  // al_ip/div_unsigned_gate.v(657)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E57929B0  (
    .a(n34[0]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [32]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [31]));  // al_ip/div_unsigned_gate.v(161)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5792AC0  (
    .a(n35[0]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [0]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [0]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [0]));  // al_ip/div_unsigned_gate.v(361)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5792BD0  (
    .a(n35[13]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [13]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [13]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [13]));  // al_ip/div_unsigned_gate.v(411)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792CE0  (
    .a(n34[13]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [45]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [44]));  // al_ip/div_unsigned_gate.v(201)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792DF0  (
    .a(n34[28]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [60]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [59]));  // al_ip/div_unsigned_gate.v(329)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5792F00  (
    .a(n34[19]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [51]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [50]));  // al_ip/div_unsigned_gate.v(249)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5793010  (
    .a(n34[23]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [55]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [54]));  // al_ip/div_unsigned_gate.v(289)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5793120  (
    .a(n35[15]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [15]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [15]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [15]));  // al_ip/div_unsigned_gate.v(431)
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'b0001))
    \u_DIV_UNSIGNED/al_00000286E5793230  (
    .a(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [1]),
    .b(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [2]),
    .o(\u_DIV_UNSIGNED/al_00000286E4688A90 ));  // al_ip/div_unsigned_gate.v(705)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5793340  (
    .a(n35[29]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [29]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [29]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [29]));  // al_ip/div_unsigned_gate.v(597)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5793450  (
    .a(n34[1]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [33]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [32]));  // al_ip/div_unsigned_gate.v(169)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5793560  (
    .a(n34[11]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [43]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [42]));  // al_ip/div_unsigned_gate.v(185)
  AL_MAP_LUT3 #(
    .EQN("(C*~(A)*~(B)+C*A*~(B)+~(C)*A*B+C*A*B)"),
    .INIT(8'b10111000))
    \u_DIV_UNSIGNED/al_00000286E5793670  (
    .a(n34[8]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E57DE2F0 [40]),
    .o(\u_DIV_UNSIGNED/al_00000286E57DEE50 [39]));  // al_ip/div_unsigned_gate.v(794)
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*~(A)*~(B)+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*~(B)+~((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C))*A*B+(D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)*A*B)"),
    .INIT(32'b10111011101110001000101110001000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5793780  (
    .a(n35[12]),
    .b(div_unsigned_start),
    .c(\u_DIV_UNSIGNED/al_00000286E5A5D8C0 ),
    .d(\u_DIV_UNSIGNED/al_00000286E57DC290 [12]),
    .e(\u_DIV_UNSIGNED/al_00000286E57E1690 [12]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E4870 [12]));  // al_ip/div_unsigned_gate.v(401)
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'b00000000000000000000000000000010),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5794000  (
    .a(\u_DIV_UNSIGNED/al_00000286E4688A90 ),
    .b(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [0]),
    .c(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [3]),
    .d(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [4]),
    .e(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [5]),
    .o(\u_DIV_UNSIGNED/al_00000286E468A980 ));  // al_ip/div_unsigned_gate.v(722)
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'b00000000000010000000000000000000),
    .LOC("UNPLACED"))
    \u_DIV_UNSIGNED/al_00000286E5794220  (
    .a(\u_DIV_UNSIGNED/al_00000286E4688A90 ),
    .b(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [0]),
    .c(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [3]),
    .d(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [4]),
    .e(\u_DIV_UNSIGNED/al_00000286E57DB3B0 [5]),
    .o(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ));  // al_ip/div_unsigned_gate.v(712)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_UNSIGNED/al_00000286E5794770  (
    .a(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .b(\u_DIV_UNSIGNED/al_00000286E468A980 ),
    .c(div_unsigned_start),
    .d(\u_DIV_UNSIGNED/al_00000286E57E03C0 [5]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E04A0 [5]));  // al_ip/div_unsigned_gate.v(732)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_UNSIGNED/al_00000286E5795540  (
    .a(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .b(\u_DIV_UNSIGNED/al_00000286E468A980 ),
    .c(div_unsigned_start),
    .d(\u_DIV_UNSIGNED/al_00000286E57E03C0 [3]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E04A0 [3]));  // al_ip/div_unsigned_gate.v(750)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_UNSIGNED/al_00000286E5796530  (
    .a(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .b(\u_DIV_UNSIGNED/al_00000286E468A980 ),
    .c(div_unsigned_start),
    .d(\u_DIV_UNSIGNED/al_00000286E57E03C0 [1]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E04A0 [1]));  // al_ip/div_unsigned_gate.v(776)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_UNSIGNED/al_00000286E5796A80  (
    .a(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .b(\u_DIV_UNSIGNED/al_00000286E468A980 ),
    .c(div_unsigned_start),
    .d(\u_DIV_UNSIGNED/al_00000286E57E03C0 [4]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E04A0 [4]));  // al_ip/div_unsigned_gate.v(741)
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'b0000000100000000))
    \u_DIV_UNSIGNED/al_00000286E5797740  (
    .a(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .b(\u_DIV_UNSIGNED/al_00000286E468A980 ),
    .c(div_unsigned_start),
    .d(\u_DIV_UNSIGNED/al_00000286E57E03C0 [2]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E04A0 [2]));  // al_ip/div_unsigned_gate.v(759)
  AL_MAP_LUT4 #(
    .EQN("~(~C*~(D*~B*~A))"),
    .INIT(16'b1111000111110000))
    \u_DIV_UNSIGNED/al_00000286E5797B80  (
    .a(\u_DIV_UNSIGNED/al_00000286E5A5E1B0 ),
    .b(\u_DIV_UNSIGNED/al_00000286E468A980 ),
    .c(div_unsigned_start),
    .d(\u_DIV_UNSIGNED/al_00000286E57E03C0 [0]),
    .o(\u_DIV_UNSIGNED/al_00000286E57E04A0 [0]));  // al_ip/div_unsigned_gate.v(785)
  AL_MAP_SEQ #(
    .CEMUX("1"),
    .CLKMUX("CLK"),
    .DFFMODE("FF"),
    .REGSET("RESET"),
    .SRMODE("ASYNC"),
    .SRMUX("INV"))
    working_reg (
    .clk(i_clk),
    .d(n8),
    .sr(i_rstn),
    .q(working));  // ../RTL/core/exu_mdu.v(52)

endmodule 

module add_sub_1  // ../RTL/core/fpu.v(83)
  (
  n1,
  n2,
  sub,
  Exception,
  Overflow,
  Underflow,
  result
  );

  input [31:0] n1;  // ../RTL/core/fpu.v(84)
  input [31:0] n2;  // ../RTL/core/fpu.v(85)
  input sub;  // ../RTL/core/fpu.v(87)
  output Exception;  // ../RTL/core/fpu.v(90)
  output Overflow;  // ../RTL/core/fpu.v(88)
  output Underflow;  // ../RTL/core/fpu.v(89)
  output [31:0] result;  // ../RTL/core/fpu.v(86)

  wire [7:0] \C023/outtemp ;  // ../RTL/core/fpu_utils.v(93)
  wire [23:0] \C03/outtemp ;  // ../RTL/core/fpu_utils.v(99)
  wire [7:0] E;  // ../RTL/core/fpu.v(95)
  wire [23:0] M_result;  // ../RTL/core/fpu.v(97)
  wire [23:0] M_result2;  // ../RTL/core/fpu.v(97)
  wire [22:0] \NM/n4 ;
  wire [7:0] exp_diff;  // ../RTL/core/fpu.v(95)
  wire \ADD01/ADD01/c1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/n10 ;
  wire \ADD01/ADD01/n20 ;
  wire \ADD01/ADD01/n3 ;
  wire \ADD01/ADD01/p2_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/p3_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/n17 ;
  wire \ADD01/ADD02/n21 ;
  wire \ADD01/ADD02/n7 ;
  wire \ADD01/ADD02/p0_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/p1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/p2_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/p3_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ctemp_lutinv ;  // ../RTL/core/fpu_utils.v(76)
  wire \ADD02/ADD01/ADD01/c0_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/p2_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/p3_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/n14 ;
  wire \ADD02/ADD01/ADD02/n7 ;
  wire \ADD02/ADD01/ADD02/p1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/n17 ;
  wire \ADD02/ADD02/ADD01/n20 ;
  wire \ADD02/ADD02/ADD01/n3 ;
  wire \ADD02/ADD02/ADD01/p0_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/p1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/p2_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/p3_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/n3 ;
  wire \ADD02/ADD02/ADD02/p0_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/p1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/p2_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/p3_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/n14 ;
  wire \ADD02/ADD03/ADD01/n3 ;
  wire \ADD02/ADD03/ADD01/p0_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/p1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/p2_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/p3_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/n1 ;
  wire \ADD02/ADD03/ADD02/n16_lutinv ;
  wire \ADD02/ADD03/ADD02/n3 ;
  wire \ADD02/ADD03/ADD02/p0_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/p1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/p2_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/p3_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD0212/ADD01/n1 ;
  wire \ADD0212/ADD01/n8 ;
  wire \ADD03/ADD01/p0_neg ;
  wire \C023/ADD01/ADD02/n0 ;
  wire \NM/add0/c11 ;  // ../RTL/core/fpu_utils.v(158)
  wire \NM/add0/c15 ;  // ../RTL/core/fpu_utils.v(158)
  wire \NM/add0/c19 ;  // ../RTL/core/fpu_utils.v(158)
  wire \NM/add0/c3 ;  // ../RTL/core/fpu_utils.v(158)
  wire \NM/add0/c7 ;  // ../RTL/core/fpu_utils.v(158)
  wire _al_u101_o;
  wire _al_u102_o;
  wire _al_u103_o;
  wire _al_u105_o;
  wire _al_u107_o;
  wire _al_u108_o;
  wire _al_u109_o;
  wire _al_u110_o;
  wire _al_u111_o;
  wire _al_u112_o;
  wire _al_u113_o;
  wire _al_u115_o;
  wire _al_u116_o;
  wire _al_u118_o;
  wire _al_u119_o;
  wire _al_u120_o;
  wire _al_u121_o;
  wire _al_u124_o;
  wire _al_u127_o;
  wire _al_u128_o;
  wire _al_u131_o;
  wire _al_u132_o;
  wire _al_u133_o;
  wire _al_u134_o;
  wire _al_u136_o;
  wire _al_u139_o;
  wire _al_u142_o;
  wire _al_u145_o;
  wire _al_u146_o;
  wire _al_u147_o;
  wire _al_u148_o;
  wire _al_u149_o;
  wire _al_u150_o;
  wire _al_u151_o;
  wire _al_u153_o;
  wire _al_u154_o;
  wire _al_u155_o;
  wire _al_u156_o;
  wire _al_u157_o;
  wire _al_u158_o;
  wire _al_u159_o;
  wire _al_u160_o;
  wire _al_u162_o;
  wire _al_u163_o;
  wire _al_u164_o;
  wire _al_u165_o;
  wire _al_u166_o;
  wire _al_u167_o;
  wire _al_u168_o;
  wire _al_u169_o;
  wire _al_u170_o;
  wire _al_u171_o;
  wire _al_u172_o;
  wire _al_u173_o;
  wire _al_u174_o;
  wire _al_u175_o;
  wire _al_u176_o;
  wire _al_u177_o;
  wire _al_u179_o;
  wire _al_u180_o;
  wire _al_u183_o;
  wire _al_u184_o;
  wire _al_u187_o;
  wire _al_u190_o;
  wire _al_u191_o;
  wire _al_u193_o;
  wire _al_u194_o;
  wire _al_u195_o;
  wire _al_u196_o;
  wire _al_u198_o;
  wire _al_u201_o;
  wire _al_u202_o;
  wire _al_u205_o;
  wire _al_u208_o;
  wire _al_u209_o;
  wire _al_u210_o;
  wire _al_u211_o;
  wire _al_u212_o;
  wire _al_u213_o;
  wire _al_u214_o;
  wire _al_u215_o;
  wire _al_u216_o;
  wire _al_u217_o;
  wire _al_u218_o;
  wire _al_u219_o;
  wire _al_u221_o;
  wire _al_u222_o;
  wire _al_u223_o;
  wire _al_u224_o;
  wire _al_u225_o;
  wire _al_u226_o;
  wire _al_u227_o;
  wire _al_u228_o;
  wire _al_u229_o;
  wire _al_u230_o;
  wire _al_u232_o;
  wire _al_u233_o;
  wire _al_u234_o;
  wire _al_u235_o;
  wire _al_u236_o;
  wire _al_u237_o;
  wire _al_u238_o;
  wire _al_u240_o;
  wire _al_u241_o;
  wire _al_u242_o;
  wire _al_u243_o;
  wire _al_u244_o;
  wire _al_u245_o;
  wire _al_u246_o;
  wire _al_u247_o;
  wire _al_u248_o;
  wire _al_u249_o;
  wire _al_u250_o;
  wire _al_u251_o;
  wire _al_u253_o;
  wire _al_u254_o;
  wire _al_u255_o;
  wire _al_u256_o;
  wire _al_u257_o;
  wire _al_u259_o;
  wire _al_u260_o;
  wire _al_u261_o;
  wire _al_u262_o;
  wire _al_u263_o;
  wire _al_u264_o;
  wire _al_u265_o;
  wire _al_u266_o;
  wire _al_u268_o;
  wire _al_u269_o;
  wire _al_u271_o;
  wire _al_u272_o;
  wire _al_u273_o;
  wire _al_u274_o;
  wire _al_u275_o;
  wire _al_u277_o;
  wire _al_u278_o;
  wire _al_u279_o;
  wire _al_u280_o;
  wire _al_u281_o;
  wire _al_u282_o;
  wire _al_u283_o;
  wire _al_u284_o;
  wire _al_u285_o;
  wire _al_u286_o;
  wire _al_u287_o;
  wire _al_u288_o;
  wire _al_u289_o;
  wire _al_u290_o;
  wire _al_u291_o;
  wire _al_u292_o;
  wire _al_u294_o;
  wire _al_u295_o;
  wire _al_u296_o;
  wire _al_u297_o;
  wire _al_u298_o;
  wire _al_u299_o;
  wire _al_u300_o;
  wire _al_u301_o;
  wire _al_u302_o;
  wire _al_u303_o;
  wire _al_u304_o;
  wire _al_u305_o;
  wire _al_u306_o;
  wire _al_u307_o;
  wire _al_u308_o;
  wire _al_u309_o;
  wire _al_u310_o;
  wire _al_u311_o;
  wire _al_u312_o;
  wire _al_u313_o;
  wire _al_u314_o;
  wire _al_u315_o;
  wire _al_u316_o;
  wire _al_u317_o;
  wire _al_u318_o;
  wire _al_u320_o;
  wire _al_u321_o;
  wire _al_u323_o;
  wire _al_u324_o;
  wire _al_u325_o;
  wire _al_u326_o;
  wire _al_u327_o;
  wire _al_u328_o;
  wire _al_u329_o;
  wire _al_u330_o;
  wire _al_u331_o;
  wire _al_u332_o;
  wire _al_u334_o;
  wire _al_u335_o;
  wire _al_u336_o;
  wire _al_u337_o;
  wire _al_u338_o;
  wire _al_u339_o;
  wire _al_u341_o;
  wire _al_u344_o;
  wire _al_u345_o;
  wire _al_u346_o;
  wire _al_u347_o;
  wire _al_u348_o;
  wire _al_u349_o;
  wire _al_u350_o;
  wire _al_u351_o;
  wire _al_u352_o;
  wire _al_u353_o;
  wire _al_u354_o;
  wire _al_u355_o;
  wire _al_u356_o;
  wire _al_u357_o;
  wire _al_u358_o;
  wire _al_u359_o;
  wire _al_u360_o;
  wire _al_u361_o;
  wire _al_u362_o;
  wire _al_u363_o;
  wire _al_u364_o;
  wire _al_u365_o;
  wire _al_u366_o;
  wire _al_u368_o;
  wire _al_u369_o;
  wire _al_u370_o;
  wire _al_u371_o;
  wire _al_u372_o;
  wire _al_u373_o;
  wire _al_u374_o;
  wire _al_u375_o;
  wire _al_u377_o;
  wire _al_u380_o;
  wire _al_u381_o;
  wire _al_u382_o;
  wire _al_u384_o;
  wire _al_u385_o;
  wire _al_u386_o;
  wire _al_u389_o;
  wire _al_u390_o;
  wire _al_u394_o;
  wire _al_u395_o;
  wire _al_u396_o;
  wire _al_u400_o;
  wire _al_u401_o;
  wire _al_u402_o;
  wire _al_u403_o;
  wire _al_u404_o;
  wire _al_u405_o;
  wire _al_u406_o;
  wire _al_u407_o;
  wire _al_u409_o;
  wire _al_u410_o;
  wire _al_u411_o;
  wire _al_u412_o;
  wire _al_u413_o;
  wire _al_u414_o;
  wire _al_u415_o;
  wire _al_u416_o;
  wire _al_u417_o;
  wire _al_u420_o;
  wire _al_u425_o;
  wire _al_u426_o;
  wire _al_u427_o;
  wire _al_u428_o;
  wire _al_u431_o;
  wire _al_u432_o;
  wire _al_u433_o;
  wire _al_u434_o;
  wire _al_u435_o;
  wire _al_u436_o;
  wire _al_u438_o;
  wire _al_u439_o;
  wire _al_u440_o;
  wire _al_u441_o;
  wire _al_u442_o;
  wire _al_u443_o;
  wire _al_u445_o;
  wire _al_u447_o;
  wire _al_u448_o;
  wire _al_u449_o;
  wire _al_u450_o;
  wire _al_u453_o;
  wire _al_u454_o;
  wire _al_u455_o;
  wire _al_u456_o;
  wire _al_u459_o;
  wire _al_u461_o;
  wire _al_u462_o;
  wire _al_u463_o;
  wire _al_u465_o;
  wire _al_u468_o;
  wire _al_u469_o;
  wire _al_u470_o;
  wire _al_u473_o;
  wire _al_u474_o;
  wire _al_u475_o;
  wire _al_u477_o;
  wire _al_u481_o;
  wire _al_u482_o;
  wire _al_u483_o;
  wire _al_u485_o;
  wire _al_u486_o;
  wire _al_u487_o;
  wire _al_u489_o;
  wire _al_u494_o;
  wire _al_u495_o;
  wire _al_u496_o;
  wire _al_u498_o;
  wire _al_u500_o;
  wire _al_u501_o;
  wire _al_u503_o;
  wire _al_u504_o;
  wire _al_u506_o;
  wire _al_u507_o;
  wire _al_u509_o;
  wire _al_u510_o;
  wire _al_u512_o;
  wire _al_u513_o;
  wire _al_u515_o;
  wire _al_u517_o;
  wire _al_u518_o;
  wire _al_u519_o;
  wire _al_u520_o;
  wire _al_u522_o;
  wire _al_u524_o;
  wire _al_u525_o;
  wire _al_u527_o;
  wire _al_u528_o;
  wire _al_u529_o;
  wire _al_u531_o;
  wire _al_u532_o;
  wire _al_u533_o;
  wire _al_u535_o;
  wire _al_u536_o;
  wire _al_u537_o;
  wire _al_u539_o;
  wire _al_u540_o;
  wire _al_u541_o;
  wire _al_u542_o;
  wire _al_u543_o;
  wire _al_u545_o;
  wire _al_u546_o;
  wire _al_u547_o;
  wire _al_u548_o;
  wire _al_u549_o;
  wire _al_u550_o;
  wire _al_u552_o;
  wire _al_u553_o;
  wire _al_u554_o;
  wire _al_u555_o;
  wire _al_u556_o;
  wire _al_u557_o;
  wire _al_u558_o;
  wire _al_u559_o;
  wire _al_u560_o;
  wire _al_u561_o;
  wire _al_u563_o;
  wire _al_u564_o;
  wire _al_u565_o;
  wire _al_u566_o;
  wire _al_u567_o;
  wire _al_u568_o;
  wire _al_u569_o;
  wire _al_u570_o;
  wire _al_u571_o;
  wire _al_u572_o;
  wire _al_u573_o;
  wire _al_u575_o;
  wire _al_u576_o;
  wire _al_u577_o;
  wire _al_u578_o;
  wire _al_u579_o;
  wire _al_u581_o;
  wire _al_u582_o;
  wire _al_u583_o;
  wire _al_u584_o;
  wire _al_u585_o;
  wire _al_u586_o;
  wire _al_u587_o;
  wire _al_u588_o;
  wire _al_u589_o;
  wire _al_u590_o;
  wire _al_u592_o;
  wire _al_u593_o;
  wire _al_u594_o;
  wire _al_u595_o;
  wire _al_u596_o;
  wire _al_u597_o;
  wire _al_u598_o;
  wire _al_u599_o;
  wire _al_u600_o;
  wire _al_u601_o;
  wire _al_u602_o;
  wire _al_u603_o;
  wire _al_u605_o;
  wire _al_u606_o;
  wire _al_u607_o;
  wire _al_u608_o;
  wire _al_u609_o;
  wire _al_u610_o;
  wire _al_u611_o;
  wire _al_u613_o;
  wire _al_u614_o;
  wire _al_u615_o;
  wire _al_u616_o;
  wire _al_u617_o;
  wire _al_u618_o;
  wire _al_u619_o;
  wire _al_u620_o;
  wire _al_u621_o;
  wire _al_u622_o;
  wire _al_u623_o;
  wire _al_u624_o;
  wire _al_u625_o;
  wire _al_u627_o;
  wire _al_u628_o;
  wire _al_u629_o;
  wire _al_u630_o;
  wire _al_u631_o;
  wire _al_u632_o;
  wire _al_u633_o;
  wire _al_u634_o;
  wire _al_u635_o;
  wire _al_u636_o;
  wire _al_u637_o;
  wire _al_u638_o;
  wire _al_u639_o;
  wire _al_u640_o;
  wire _al_u641_o;
  wire _al_u642_o;
  wire _al_u643_o;
  wire _al_u644_o;
  wire _al_u645_o;
  wire _al_u646_o;
  wire _al_u648_o;
  wire _al_u649_o;
  wire _al_u64_o;
  wire _al_u650_o;
  wire _al_u651_o;
  wire _al_u652_o;
  wire _al_u653_o;
  wire _al_u654_o;
  wire _al_u655_o;
  wire _al_u657_o;
  wire _al_u658_o;
  wire _al_u659_o;
  wire _al_u660_o;
  wire _al_u661_o;
  wire _al_u662_o;
  wire _al_u663_o;
  wire _al_u664_o;
  wire _al_u665_o;
  wire _al_u666_o;
  wire _al_u667_o;
  wire _al_u668_o;
  wire _al_u669_o;
  wire _al_u670_o;
  wire _al_u671_o;
  wire _al_u673_o;
  wire _al_u674_o;
  wire _al_u675_o;
  wire _al_u676_o;
  wire _al_u677_o;
  wire _al_u678_o;
  wire _al_u679_o;
  wire _al_u67_o;
  wire _al_u680_o;
  wire _al_u681_o;
  wire _al_u682_o;
  wire _al_u683_o;
  wire _al_u684_o;
  wire _al_u685_o;
  wire _al_u686_o;
  wire _al_u688_o;
  wire _al_u689_o;
  wire _al_u68_o;
  wire _al_u690_o;
  wire _al_u691_o;
  wire _al_u692_o;
  wire _al_u693_o;
  wire _al_u694_o;
  wire _al_u695_o;
  wire _al_u696_o;
  wire _al_u697_o;
  wire _al_u698_o;
  wire _al_u699_o;
  wire _al_u700_o;
  wire _al_u701_o;
  wire _al_u702_o;
  wire _al_u703_o;
  wire _al_u704_o;
  wire _al_u705_o;
  wire _al_u707_o;
  wire _al_u708_o;
  wire _al_u709_o;
  wire _al_u710_o;
  wire _al_u711_o;
  wire _al_u712_o;
  wire _al_u713_o;
  wire _al_u714_o;
  wire _al_u715_o;
  wire _al_u716_o;
  wire _al_u717_o;
  wire _al_u718_o;
  wire _al_u719_o;
  wire _al_u71_o;
  wire _al_u720_o;
  wire _al_u721_o;
  wire _al_u722_o;
  wire _al_u723_o;
  wire _al_u724_o;
  wire _al_u725_o;
  wire _al_u727_o;
  wire _al_u728_o;
  wire _al_u729_o;
  wire _al_u730_o;
  wire _al_u731_o;
  wire _al_u732_o;
  wire _al_u733_o;
  wire _al_u734_o;
  wire _al_u735_o;
  wire _al_u736_o;
  wire _al_u737_o;
  wire _al_u738_o;
  wire _al_u739_o;
  wire _al_u741_o;
  wire _al_u742_o;
  wire _al_u743_o;
  wire _al_u744_o;
  wire _al_u745_o;
  wire _al_u746_o;
  wire _al_u747_o;
  wire _al_u748_o;
  wire _al_u749_o;
  wire _al_u74_o;
  wire _al_u750_o;
  wire _al_u751_o;
  wire _al_u752_o;
  wire _al_u753_o;
  wire _al_u754_o;
  wire _al_u755_o;
  wire _al_u756_o;
  wire _al_u757_o;
  wire _al_u758_o;
  wire _al_u759_o;
  wire _al_u760_o;
  wire _al_u762_o;
  wire _al_u763_o;
  wire _al_u764_o;
  wire _al_u765_o;
  wire _al_u766_o;
  wire _al_u767_o;
  wire _al_u768_o;
  wire _al_u769_o;
  wire _al_u770_o;
  wire _al_u771_o;
  wire _al_u772_o;
  wire _al_u773_o;
  wire _al_u774_o;
  wire _al_u775_o;
  wire _al_u776_o;
  wire _al_u778_o;
  wire _al_u779_o;
  wire _al_u77_o;
  wire _al_u780_o;
  wire _al_u781_o;
  wire _al_u782_o;
  wire _al_u783_o;
  wire _al_u784_o;
  wire _al_u785_o;
  wire _al_u786_o;
  wire _al_u787_o;
  wire _al_u788_o;
  wire _al_u789_o;
  wire _al_u78_o;
  wire _al_u790_o;
  wire _al_u791_o;
  wire _al_u793_o;
  wire _al_u794_o;
  wire _al_u795_o;
  wire _al_u796_o;
  wire _al_u797_o;
  wire _al_u798_o;
  wire _al_u801_o;
  wire _al_u802_o;
  wire _al_u803_o;
  wire _al_u804_o;
  wire _al_u805_o;
  wire _al_u806_o;
  wire _al_u807_o;
  wire _al_u808_o;
  wire _al_u809_o;
  wire _al_u811_o;
  wire _al_u812_o;
  wire _al_u813_o;
  wire _al_u814_o;
  wire _al_u817_o;
  wire _al_u818_o;
  wire _al_u820_o;
  wire _al_u821_o;
  wire _al_u822_o;
  wire _al_u823_o;
  wire _al_u824_o;
  wire _al_u827_o;
  wire _al_u828_o;
  wire _al_u829_o;
  wire _al_u82_o;
  wire _al_u830_o;
  wire _al_u832_o;
  wire _al_u833_o;
  wire _al_u834_o;
  wire _al_u835_o;
  wire _al_u837_o;
  wire _al_u838_o;
  wire _al_u840_o;
  wire _al_u841_o;
  wire _al_u842_o;
  wire _al_u844_o;
  wire _al_u846_o;
  wire _al_u847_o;
  wire _al_u848_o;
  wire _al_u849_o;
  wire _al_u92_o;
  wire _al_u93_o;
  wire _al_u95_o;
  wire _al_u96_o;
  wire _al_u98_o;
  wire n100_lutinv;
  wire n101_lutinv;
  wire n102_lutinv;
  wire n103_lutinv;
  wire n104_lutinv;
  wire n105_lutinv;
  wire n106_lutinv;
  wire n107_lutinv;
  wire n198_lutinv;
  wire n221_lutinv;
  wire n222_lutinv;
  wire n223_lutinv;
  wire n224_lutinv;
  wire n225_lutinv;
  wire n226_lutinv;
  wire n227_lutinv;
  wire n228_lutinv;
  wire n229_lutinv;
  wire n230_lutinv;
  wire n231_lutinv;
  wire n232_lutinv;
  wire n233_lutinv;
  wire n234_lutinv;
  wire n235_lutinv;
  wire n236_lutinv;
  wire n237_lutinv;
  wire n238_lutinv;
  wire n239_lutinv;
  wire n86_lutinv;
  wire n87_lutinv;
  wire n89_lutinv;
  wire n90_lutinv;
  wire n91_lutinv;
  wire n92_lutinv;
  wire n93_lutinv;
  wire n94_lutinv;
  wire n95_lutinv;
  wire n96_lutinv;
  wire n97_lutinv;
  wire n98_lutinv;
  wire n99_lutinv;
  wire u194_sel_is_0_o;

  assign result[23] = \ADD03/ADD01/p0_neg ;
  EG_PHY_LSLICE #(
    //.MACRO("NM/add0/ucin_al_u852"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \NM/add0/u11_al_u855  (
    .a({M_result2[14],M_result2[12]}),
    .b({M_result2[15],M_result2[13]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\NM/add0/c11 ),
    .f({\NM/n4 [13],\NM/n4 [11]}),
    .fco(\NM/add0/c15 ),
    .fx({\NM/n4 [14],\NM/n4 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("NM/add0/ucin_al_u852"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \NM/add0/u15_al_u856  (
    .a({M_result2[18],M_result2[16]}),
    .b({M_result2[19],M_result2[17]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\NM/add0/c15 ),
    .f({\NM/n4 [17],\NM/n4 [15]}),
    .fco(\NM/add0/c19 ),
    .fx({\NM/n4 [18],\NM/n4 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("NM/add0/ucin_al_u852"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \NM/add0/u19_al_u857  (
    .a({M_result2[22],M_result2[20]}),
    .b({M_result2[23],M_result2[21]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\NM/add0/c19 ),
    .f({\NM/n4 [21],\NM/n4 [19]}),
    .fx({\NM/n4 [22],\NM/n4 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("NM/add0/ucin_al_u852"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \NM/add0/u3_al_u853  (
    .a({M_result2[6],M_result2[4]}),
    .b({M_result2[7],M_result2[5]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\NM/add0/c3 ),
    .f({\NM/n4 [5],\NM/n4 [3]}),
    .fco(\NM/add0/c7 ),
    .fx({\NM/n4 [6],\NM/n4 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("NM/add0/ucin_al_u852"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \NM/add0/u7_al_u854  (
    .a({M_result2[10],M_result2[8]}),
    .b({M_result2[11],M_result2[9]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\NM/add0/c7 ),
    .f({\NM/n4 [9],\NM/n4 [7]}),
    .fco(\NM/add0/c11 ),
    .fx({\NM/n4 [10],\NM/n4 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("NM/add0/ucin_al_u852"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \NM/add0/ucin_al_u852  (
    .a({M_result2[2],1'b0}),
    .b({M_result2[3],M_result2[1]}),
    .c(2'b00),
    .d(2'b01),
    .e({1'b0,M_result[0]}),
    .f({\NM/n4 [1],open_n108}),
    .fco(\NM/add0/c3 ),
    .fx({\NM/n4 [2],\NM/n4 [0]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u100 (
    .a(_al_u64_o),
    .b(n2[17]),
    .c(n2[16]),
    .o(n225_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u101 (
    .a(n223_lutinv),
    .b(n225_lutinv),
    .c(_al_u67_o),
    .o(_al_u101_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(16'h0a03))
    _al_u102 (
    .a(_al_u98_o),
    .b(_al_u101_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u102_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(B*(A*~(D)*~(E)+~(A)*D*~(E)+A*D*~(E)+A*D*E)))"),
    .INIT(32'h70f03070))
    _al_u103 (
    .a(\ADD01/ctemp_lutinv ),
    .b(\ADD01/ADD02/n17 ),
    .c(_al_u78_o),
    .d(n1[27]),
    .e(n2[27]),
    .o(_al_u103_o));
  AL_MAP_LUT3 #(
    .EQN("(B@(~C*A))"),
    .INIT(8'hc6))
    _al_u104 (
    .a(_al_u103_o),
    .b(_al_u67_o),
    .c(_al_u64_o),
    .o(exp_diff[1]));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u105 (
    .a(_al_u64_o),
    .b(n2[1]),
    .c(n2[0]),
    .o(_al_u105_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u106 (
    .a(_al_u64_o),
    .b(n2[3]),
    .c(n2[2]),
    .o(n239_lutinv));
  AL_MAP_LUT5 #(
    .EQN("(~C*~B*(~D*~(E)*~(A)+~D*E*~(A)+~(~D)*E*A+~D*E*A))"),
    .INIT(32'h02030001))
    _al_u107 (
    .a(exp_diff[1]),
    .b(exp_diff[3]),
    .c(exp_diff[2]),
    .d(_al_u105_o),
    .e(n239_lutinv),
    .o(_al_u107_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u108 (
    .a(\ADD01/ADD02/g0 ),
    .b(\ADD01/ctemp_lutinv ),
    .o(_al_u108_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u109 (
    .a(n1[27]),
    .b(n2[27]),
    .o(_al_u109_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C)*~((~D*~A))+~(B)*C*~((~D*~A))+B*C*~((~D*~A))+~(B)*~(C)*(~D*~A)+B*~(C)*(~D*~A)+~(B)*C*(~D*~A))"),
    .INIT(16'hfcbd))
    _al_u110 (
    .a(_al_u108_o),
    .b(_al_u78_o),
    .c(\ADD01/ADD02/p1_lutinv ),
    .d(_al_u109_o),
    .o(_al_u110_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h7f133701))
    _al_u111 (
    .a(\ADD01/ADD02/g0 ),
    .b(n1[29]),
    .c(n1[28]),
    .d(n2[29]),
    .e(n2[28]),
    .o(_al_u111_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@(B*~(E*C*A)))"),
    .INIT(32'h4cb3cc33))
    _al_u112 (
    .a(\ADD01/ctemp_lutinv ),
    .b(_al_u111_o),
    .c(\ADD01/ADD02/n7 ),
    .d(\ADD01/ADD02/p3_lutinv ),
    .e(\ADD01/ADD02/p0_lutinv ),
    .o(_al_u112_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+~(A)*B*C)"),
    .INIT(8'h71))
    _al_u113 (
    .a(\ADD01/ADD02/g0 ),
    .b(n1[28]),
    .c(n2[28]),
    .o(_al_u113_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u114 (
    .a(n1[29]),
    .b(n2[29]),
    .o(\ADD01/ADD02/p2_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("~(C@(B*~(E*D*A)))"),
    .INIT(32'h4bc3c3c3))
    _al_u115 (
    .a(\ADD01/ctemp_lutinv ),
    .b(_al_u113_o),
    .c(\ADD01/ADD02/p2_lutinv ),
    .d(\ADD01/ADD02/p1_lutinv ),
    .e(\ADD01/ADD02/p0_lutinv ),
    .o(_al_u115_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u116 (
    .a(_al_u110_o),
    .b(_al_u112_o),
    .c(_al_u115_o),
    .o(_al_u116_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E@D))"),
    .INIT(32'h80000080))
    _al_u117 (
    .a(\ADD01/ADD01/p3_lutinv ),
    .b(\ADD01/ADD01/p2_lutinv ),
    .c(_al_u64_o),
    .d(n1[24]),
    .e(n2[24]),
    .o(\ADD01/ADD01/n20 ));
  AL_MAP_LUT4 #(
    .EQN("(C@(A*~(B)*~(D)+A*B*~(D)+~(A)*~(B)*D+~(A)*B*D+A*B*D))"),
    .INIT(16'h2d5a))
    _al_u118 (
    .a(\ADD01/ctemp_lutinv ),
    .b(\ADD01/ADD01/n20 ),
    .c(\ADD01/ADD02/p0_lutinv ),
    .d(_al_u103_o),
    .o(_al_u118_o));
  AL_MAP_LUT5 #(
    .EQN("(D*(~(~C*A)*~(B)*~(E)+~(~C*A)*B*~(E)+~(~(~C*A))*B*E+~(~C*A)*B*E))"),
    .INIT(32'hcc00f500))
    _al_u119 (
    .a(_al_u95_o),
    .b(_al_u102_o),
    .c(_al_u107_o),
    .d(_al_u116_o),
    .e(_al_u118_o),
    .o(_al_u119_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u120 (
    .a(n1[26]),
    .b(n1[25]),
    .c(n1[24]),
    .d(n1[23]),
    .o(_al_u120_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u121 (
    .a(_al_u120_o),
    .b(n1[30]),
    .c(n1[29]),
    .d(n1[28]),
    .e(n1[27]),
    .o(_al_u121_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u122 (
    .a(_al_u121_o),
    .b(_al_u64_o),
    .c(n1[22]),
    .o(n87_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u123 (
    .a(_al_u64_o),
    .b(n1[21]),
    .c(n1[20]),
    .o(n89_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'hacca))
    _al_u124 (
    .a(n87_lutinv),
    .b(n89_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u124_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u125 (
    .a(_al_u64_o),
    .b(n1[19]),
    .c(n1[18]),
    .o(n91_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u126 (
    .a(_al_u64_o),
    .b(n1[17]),
    .c(n1[16]),
    .o(n93_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u127 (
    .a(n91_lutinv),
    .b(n93_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u127_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u128 (
    .a(_al_u124_o),
    .b(_al_u127_o),
    .c(exp_diff[2]),
    .o(_al_u128_o));
  AL_MAP_LUT3 #(
    .EQN("~(B@(~C*~A))"),
    .INIT(8'h36))
    _al_u129 (
    .a(_al_u108_o),
    .b(\ADD01/ADD02/p1_lutinv ),
    .c(_al_u109_o),
    .o(\C023/outtemp [5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u130 (
    .a(\ADD01/ADD01/n20 ),
    .b(\ADD01/ADD02/p0_lutinv ),
    .o(\C023/ADD01/ADD02/n0 ));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*~A)"),
    .INIT(32'h10000000))
    _al_u131 (
    .a(\C023/outtemp [5]),
    .b(\C023/ADD01/ADD02/n0 ),
    .c(_al_u103_o),
    .d(_al_u112_o),
    .e(_al_u115_o),
    .o(_al_u131_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u132 (
    .a(exp_diff[3]),
    .b(_al_u118_o),
    .o(_al_u132_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u133 (
    .a(_al_u103_o),
    .b(n1[0]),
    .o(_al_u133_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*B*~A))"),
    .INIT(16'h00bf))
    _al_u134 (
    .a(_al_u128_o),
    .b(_al_u131_o),
    .c(_al_u132_o),
    .d(_al_u133_o),
    .o(_al_u134_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u135 (
    .a(_al_u64_o),
    .b(n1[3]),
    .c(n1[2]),
    .o(n107_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h717d))
    _al_u136 (
    .a(n107_lutinv),
    .b(_al_u67_o),
    .c(_al_u64_o),
    .d(n1[1]),
    .o(_al_u136_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u137 (
    .a(_al_u64_o),
    .b(n1[7]),
    .c(n1[6]),
    .o(n103_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u138 (
    .a(_al_u64_o),
    .b(n1[5]),
    .c(n1[4]),
    .o(n105_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u139 (
    .a(n103_lutinv),
    .b(n105_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u139_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u140 (
    .a(_al_u64_o),
    .b(n1[15]),
    .c(n1[14]),
    .o(n95_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u141 (
    .a(_al_u64_o),
    .b(n1[13]),
    .c(n1[12]),
    .o(n97_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u142 (
    .a(n95_lutinv),
    .b(n97_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u142_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u143 (
    .a(_al_u64_o),
    .b(n1[11]),
    .c(n1[10]),
    .o(n99_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u144 (
    .a(_al_u64_o),
    .b(n1[9]),
    .c(n1[8]),
    .o(n101_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u145 (
    .a(n99_lutinv),
    .b(n101_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u145_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u146 (
    .a(_al_u142_o),
    .b(_al_u145_o),
    .c(exp_diff[2]),
    .d(exp_diff[3]),
    .o(_al_u146_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u147 (
    .a(_al_u136_o),
    .b(_al_u139_o),
    .c(_al_u146_o),
    .d(exp_diff[3]),
    .o(_al_u147_o));
  AL_MAP_LUT3 #(
    .EQN("(A@(~C*B))"),
    .INIT(8'ha6))
    _al_u148 (
    .a(\ADD01/ADD02/p1_lutinv ),
    .b(n1[27]),
    .c(n2[27]),
    .o(_al_u148_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u149 (
    .a(\C023/ADD01/ADD02/n0 ),
    .b(_al_u112_o),
    .c(_al_u115_o),
    .o(_al_u149_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*~A)"),
    .INIT(16'h4000))
    _al_u150 (
    .a(_al_u118_o),
    .b(_al_u148_o),
    .c(_al_u103_o),
    .d(_al_u149_o),
    .o(_al_u150_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u151 (
    .a(_al_u103_o),
    .b(n2[0]),
    .o(_al_u151_o));
  AL_MAP_LUT5 #(
    .EQN("((~E*~A)@(~(D*~C)*B))"),
    .INIT(32'hc0cc9599))
    _al_u152 (
    .a(_al_u119_o),
    .b(_al_u134_o),
    .c(_al_u147_o),
    .d(_al_u150_o),
    .e(_al_u151_o),
    .o(M_result[0]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u153 (
    .a(n89_lutinv),
    .b(n91_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u153_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(A)*~((D@C))+B*A*~((D@C))+~(B)*A*(D@C)+B*A*(D@C))"),
    .INIT(16'h3553))
    _al_u154 (
    .a(n95_lutinv),
    .b(n93_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u154_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hafc0))
    _al_u155 (
    .a(_al_u153_o),
    .b(_al_u154_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u155_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u156 (
    .a(n97_lutinv),
    .b(n99_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u156_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~B*~A))"),
    .INIT(16'h00ef))
    _al_u157 (
    .a(_al_u156_o),
    .b(exp_diff[3]),
    .c(exp_diff[2]),
    .d(_al_u118_o),
    .o(_al_u157_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(A)*~((D@C))+B*A*~((D@C))+~(B)*A*(D@C)+B*A*(D@C))"),
    .INIT(16'h3553))
    _al_u158 (
    .a(n103_lutinv),
    .b(n101_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u158_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~A*~(~D*C)))"),
    .INIT(16'h88c8))
    _al_u159 (
    .a(_al_u155_o),
    .b(_al_u157_o),
    .c(_al_u158_o),
    .d(exp_diff[3]),
    .o(_al_u159_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u160 (
    .a(n87_lutinv),
    .b(_al_u67_o),
    .c(_al_u64_o),
    .o(_al_u160_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u161 (
    .a(\ADD01/ctemp_lutinv ),
    .b(\ADD01/ADD02/n17 ),
    .c(\ADD01/ADD02/p0_lutinv ),
    .o(\ADD01/ADD02/n21 ));
  AL_MAP_LUT4 #(
    .EQN("(~((B*~A))*~(C)*~(D)+(B*~A)*~(C)*~(D)+(B*~A)*C*~(D)+~((B*~A))*~(C)*D+~((B*~A))*C*D+(B*~A)*C*D)"),
    .INIT(16'hfb4f))
    _al_u162 (
    .a(\ADD01/ADD02/n21 ),
    .b(_al_u92_o),
    .c(\C023/outtemp [3]),
    .d(_al_u93_o),
    .o(_al_u162_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*B)))"),
    .INIT(16'h08aa))
    _al_u163 (
    .a(_al_u131_o),
    .b(_al_u160_o),
    .c(_al_u162_o),
    .d(_al_u118_o),
    .o(_al_u163_o));
  AL_MAP_LUT4 #(
    .EQN("~(C*~((D*~A))*~(B)+C*(D*~A)*~(B)+~(C)*(D*~A)*B+C*(D*~A)*B)"),
    .INIT(16'h8bcf))
    _al_u164 (
    .a(_al_u159_o),
    .b(_al_u103_o),
    .c(n1[6]),
    .d(_al_u163_o),
    .o(_al_u164_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u165 (
    .a(exp_diff[2]),
    .b(_al_u96_o),
    .c(_al_u67_o),
    .o(_al_u165_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u166 (
    .a(_al_u103_o),
    .b(n2[6]),
    .o(_al_u166_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(E*~D*B*A))"),
    .INIT(32'h0f070f0f))
    _al_u167 (
    .a(_al_u165_o),
    .b(_al_u116_o),
    .c(_al_u166_o),
    .d(exp_diff[3]),
    .e(_al_u118_o),
    .o(_al_u167_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u168 (
    .a(\C023/outtemp [5]),
    .b(_al_u112_o),
    .c(_al_u115_o),
    .o(_al_u168_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u169 (
    .a(\C023/outtemp [3]),
    .b(_al_u93_o),
    .o(_al_u169_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u170 (
    .a(n229_lutinv),
    .b(n231_lutinv),
    .c(_al_u67_o),
    .o(_al_u170_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*A*~(C*B))"),
    .INIT(32'h0000002a))
    _al_u171 (
    .a(_al_u168_o),
    .b(_al_u169_o),
    .c(_al_u170_o),
    .d(_al_u118_o),
    .e(_al_u103_o),
    .o(_al_u171_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u172 (
    .a(n221_lutinv),
    .b(n223_lutinv),
    .c(_al_u67_o),
    .o(_al_u172_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u173 (
    .a(n225_lutinv),
    .b(n227_lutinv),
    .c(_al_u67_o),
    .o(_al_u173_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u174 (
    .a(_al_u172_o),
    .b(_al_u173_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u174_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u175 (
    .a(n233_lutinv),
    .b(n235_lutinv),
    .c(_al_u67_o),
    .o(_al_u175_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u176 (
    .a(_al_u175_o),
    .b(exp_diff[3]),
    .c(exp_diff[2]),
    .o(_al_u176_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~C*B))"),
    .INIT(16'haaa2))
    _al_u177 (
    .a(_al_u167_o),
    .b(_al_u171_o),
    .c(_al_u174_o),
    .d(_al_u176_o),
    .o(_al_u177_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u178 (
    .a(_al_u64_o),
    .b(n2[20]),
    .c(n2[19]),
    .o(n222_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u179 (
    .a(_al_u64_o),
    .b(n2[22]),
    .c(n2[21]),
    .o(_al_u179_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(B)*~(C)+~A*B*~(C)+~(~A)*B*C+~A*B*C)"),
    .INIT(8'hc5))
    _al_u180 (
    .a(n222_lutinv),
    .b(_al_u179_o),
    .c(_al_u67_o),
    .o(_al_u180_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u181 (
    .a(_al_u64_o),
    .b(n2[18]),
    .c(n2[17]),
    .o(n224_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u182 (
    .a(_al_u64_o),
    .b(n2[16]),
    .c(n2[15]),
    .o(n226_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u183 (
    .a(n224_lutinv),
    .b(n226_lutinv),
    .c(_al_u67_o),
    .o(_al_u183_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u184 (
    .a(_al_u180_o),
    .b(_al_u183_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u184_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u185 (
    .a(_al_u64_o),
    .b(n2[14]),
    .c(n2[13]),
    .o(n228_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u186 (
    .a(_al_u64_o),
    .b(n2[12]),
    .c(n2[11]),
    .o(n230_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u187 (
    .a(n228_lutinv),
    .b(n230_lutinv),
    .c(_al_u67_o),
    .o(_al_u187_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u188 (
    .a(_al_u64_o),
    .b(n2[10]),
    .c(n2[9]),
    .o(n232_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u189 (
    .a(_al_u64_o),
    .b(n2[8]),
    .c(n2[7]),
    .o(n234_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u190 (
    .a(n232_lutinv),
    .b(n234_lutinv),
    .c(_al_u67_o),
    .o(_al_u190_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)))"),
    .INIT(32'h0000f5f3))
    _al_u191 (
    .a(_al_u187_o),
    .b(_al_u190_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .e(_al_u118_o),
    .o(_al_u191_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u192 (
    .a(_al_u93_o),
    .b(_al_u121_o),
    .c(\ADD01/ADD01/n3 ),
    .o(n198_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u193 (
    .a(exp_diff[3]),
    .b(_al_u118_o),
    .c(n198_lutinv),
    .o(_al_u193_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u194 (
    .a(_al_u103_o),
    .b(n2[7]),
    .o(_al_u194_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*~(~C*~(B*~A))))"),
    .INIT(32'h00000bff))
    _al_u195 (
    .a(_al_u184_o),
    .b(_al_u191_o),
    .c(_al_u193_o),
    .d(_al_u116_o),
    .e(_al_u194_o),
    .o(_al_u195_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u196 (
    .a(_al_u64_o),
    .b(n1[22]),
    .c(n1[21]),
    .o(_al_u196_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u197 (
    .a(_al_u64_o),
    .b(n1[20]),
    .c(n1[19]),
    .o(n90_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~(B)*~((D@C))+~A*B*~((D@C))+~(~A)*B*(D@C)+~A*B*(D@C))"),
    .INIT(16'ha33a))
    _al_u198 (
    .a(_al_u196_o),
    .b(n90_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u198_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u199 (
    .a(_al_u64_o),
    .b(n1[18]),
    .c(n1[17]),
    .o(n92_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u200 (
    .a(_al_u64_o),
    .b(n1[16]),
    .c(n1[15]),
    .o(n94_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u201 (
    .a(n92_lutinv),
    .b(n94_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u201_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u202 (
    .a(_al_u198_o),
    .b(_al_u201_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u202_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u203 (
    .a(_al_u64_o),
    .b(n1[14]),
    .c(n1[13]),
    .o(n96_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u204 (
    .a(_al_u64_o),
    .b(n1[12]),
    .c(n1[11]),
    .o(n98_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u205 (
    .a(n96_lutinv),
    .b(n98_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u205_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u206 (
    .a(_al_u64_o),
    .b(n1[10]),
    .c(n1[9]),
    .o(n100_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u207 (
    .a(_al_u64_o),
    .b(n1[8]),
    .c(n1[7]),
    .o(n102_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u208 (
    .a(n100_lutinv),
    .b(n102_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u208_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)))"),
    .INIT(32'h0000f5f3))
    _al_u209 (
    .a(_al_u205_o),
    .b(_al_u208_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .e(_al_u118_o),
    .o(_al_u209_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u210 (
    .a(_al_u103_o),
    .b(n1[7]),
    .o(_al_u210_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*~(~D*~(B*~A))))"),
    .INIT(32'h00000fbf))
    _al_u211 (
    .a(_al_u202_o),
    .b(_al_u209_o),
    .c(_al_u131_o),
    .d(_al_u193_o),
    .e(_al_u210_o),
    .o(_al_u211_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u212 (
    .a(n1[31]),
    .b(n2[31]),
    .o(_al_u212_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hbf0bfee0))
    _al_u213 (
    .a(_al_u164_o),
    .b(_al_u177_o),
    .c(_al_u195_o),
    .d(_al_u211_o),
    .e(_al_u212_o),
    .o(_al_u213_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*A))"),
    .INIT(8'h07))
    _al_u214 (
    .a(_al_u131_o),
    .b(_al_u193_o),
    .c(_al_u210_o),
    .o(_al_u214_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u215 (
    .a(_al_u205_o),
    .b(_al_u208_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u215_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(A*~(D*~C*~B)))"),
    .INIT(32'h5755a8aa))
    _al_u216 (
    .a(_al_u214_o),
    .b(_al_u202_o),
    .c(_al_u215_o),
    .d(_al_u150_o),
    .e(_al_u212_o),
    .o(_al_u216_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(C*~(~B*~(~E*D))))"),
    .INIT(32'h2a2a0a2a))
    _al_u217 (
    .a(_al_u163_o),
    .b(_al_u155_o),
    .c(_al_u157_o),
    .d(_al_u158_o),
    .e(exp_diff[3]),
    .o(_al_u217_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(A*~(~D*~C*B)))"),
    .INIT(32'h555daaa2))
    _al_u218 (
    .a(_al_u167_o),
    .b(_al_u171_o),
    .c(_al_u174_o),
    .d(_al_u176_o),
    .e(_al_u212_o),
    .o(_al_u218_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u219 (
    .a(_al_u103_o),
    .b(n1[6]),
    .o(_al_u219_o));
  AL_MAP_LUT5 #(
    .EQN("(((~E*~B)@C)*(D@A))"),
    .INIT(32'h50a04182))
    _al_u220 (
    .a(_al_u216_o),
    .b(_al_u217_o),
    .c(_al_u218_o),
    .d(_al_u195_o),
    .e(_al_u219_o),
    .o(\ADD02/ADD01/ADD02/n14 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*B)))"),
    .INIT(16'h08aa))
    _al_u221 (
    .a(_al_u131_o),
    .b(_al_u124_o),
    .c(_al_u162_o),
    .d(_al_u118_o),
    .o(_al_u221_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'hc0a0))
    _al_u222 (
    .a(_al_u142_o),
    .b(_al_u127_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u222_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(A*~(B)*~(D)+A*B*~(D)+~(A)*B*D+A*B*D))"),
    .INIT(16'h0c0a))
    _al_u223 (
    .a(_al_u139_o),
    .b(_al_u145_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u223_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u224 (
    .a(_al_u103_o),
    .b(n1[4]),
    .o(_al_u224_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(A*~(~E*~(~C*~B))))"),
    .INIT(32'h005500fd))
    _al_u225 (
    .a(_al_u221_o),
    .b(_al_u222_o),
    .c(_al_u223_o),
    .d(_al_u224_o),
    .e(_al_u118_o),
    .o(_al_u225_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h550f33ff))
    _al_u226 (
    .a(_al_u101_o),
    .b(_al_u68_o),
    .c(_al_u71_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u226_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*B)))"),
    .INIT(16'h08aa))
    _al_u227 (
    .a(_al_u116_o),
    .b(_al_u98_o),
    .c(_al_u162_o),
    .d(_al_u118_o),
    .o(_al_u227_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u228 (
    .a(_al_u162_o),
    .b(_al_u74_o),
    .o(_al_u228_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u229 (
    .a(_al_u103_o),
    .b(n2[4]),
    .o(_al_u229_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(B*~(~E*~(~C*A))))"),
    .INIT(32'h003300f7))
    _al_u230 (
    .a(_al_u226_o),
    .b(_al_u227_o),
    .c(_al_u228_o),
    .d(_al_u229_o),
    .e(_al_u118_o),
    .o(_al_u230_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D@C@B))"),
    .INIT(16'h1441))
    _al_u231 (
    .a(_al_u225_o),
    .b(_al_u230_o),
    .c(n1[31]),
    .d(n2[31]),
    .o(\ADD02/ADD01/ADD02/g0 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u232 (
    .a(_al_u67_o),
    .b(_al_u64_o),
    .o(_al_u232_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u233 (
    .a(_al_u179_o),
    .b(_al_u67_o),
    .o(_al_u233_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~(~D*~(~C*~B))))"),
    .INIT(32'h00a8aaaa))
    _al_u234 (
    .a(_al_u116_o),
    .b(_al_u232_o),
    .c(_al_u233_o),
    .d(_al_u162_o),
    .e(_al_u118_o),
    .o(_al_u234_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u235 (
    .a(n222_lutinv),
    .b(n224_lutinv),
    .c(_al_u67_o),
    .o(_al_u235_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u236 (
    .a(n226_lutinv),
    .b(n228_lutinv),
    .c(_al_u67_o),
    .o(_al_u236_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u237 (
    .a(n230_lutinv),
    .b(n232_lutinv),
    .c(_al_u67_o),
    .o(_al_u237_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h550f33ff))
    _al_u238 (
    .a(_al_u235_o),
    .b(_al_u236_o),
    .c(_al_u237_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u238_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u239 (
    .a(_al_u64_o),
    .b(n2[6]),
    .c(n2[5]),
    .o(n236_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u240 (
    .a(n234_lutinv),
    .b(n236_lutinv),
    .c(_al_u67_o),
    .o(_al_u240_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u241 (
    .a(_al_u162_o),
    .b(_al_u240_o),
    .o(_al_u241_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u242 (
    .a(_al_u103_o),
    .b(n2[5]),
    .o(_al_u242_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(A*~(~E*~(~C*B))))"),
    .INIT(32'h005500f7))
    _al_u243 (
    .a(_al_u234_o),
    .b(_al_u238_o),
    .c(_al_u241_o),
    .d(_al_u242_o),
    .e(_al_u118_o),
    .o(_al_u243_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u244 (
    .a(_al_u243_o),
    .b(_al_u212_o),
    .o(_al_u244_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(~D*~(A)*~(C)+~D*A*~(C)+~(~D)*A*C+~D*A*C))"),
    .INIT(16'h4c40))
    _al_u245 (
    .a(_al_u121_o),
    .b(_al_u67_o),
    .c(_al_u64_o),
    .d(n1[22]),
    .o(_al_u245_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u246 (
    .a(_al_u196_o),
    .b(_al_u67_o),
    .c(_al_u64_o),
    .o(_al_u246_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~(~B*~(~D*~C))))"),
    .INIT(32'h2220aaaa))
    _al_u247 (
    .a(_al_u131_o),
    .b(_al_u162_o),
    .c(_al_u245_o),
    .d(_al_u246_o),
    .e(_al_u118_o),
    .o(_al_u247_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u248 (
    .a(n90_lutinv),
    .b(n92_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u248_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u249 (
    .a(n94_lutinv),
    .b(n96_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u249_o));
  AL_MAP_LUT4 #(
    .EQN("(C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'ha0c0))
    _al_u250 (
    .a(_al_u248_o),
    .b(_al_u249_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u250_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u251 (
    .a(n98_lutinv),
    .b(n100_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u251_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u252 (
    .a(_al_u64_o),
    .b(n1[6]),
    .c(n1[5]),
    .o(n104_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u253 (
    .a(n102_lutinv),
    .b(n104_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u253_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u254 (
    .a(_al_u251_o),
    .b(_al_u253_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u254_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u255 (
    .a(_al_u103_o),
    .b(n1[5]),
    .o(_al_u255_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(A*~(~E*~(~C*~B))))"),
    .INIT(32'h005500fd))
    _al_u256 (
    .a(_al_u247_o),
    .b(_al_u250_o),
    .c(_al_u254_o),
    .d(_al_u255_o),
    .e(_al_u118_o),
    .o(_al_u256_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B*(~(C)*~(D)*~(E)+C*~(D)*~(E)+C*D*~(E)+C*~(D)*E)))"),
    .INIT(32'haa2a2a22))
    _al_u257 (
    .a(_al_u213_o),
    .b(\ADD02/ADD01/ADD02/n14 ),
    .c(\ADD02/ADD01/ADD02/g0 ),
    .d(_al_u244_o),
    .e(_al_u256_o),
    .o(_al_u257_o));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u258 (
    .a(_al_u256_o),
    .b(_al_u243_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD01/ADD02/p1_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("~(E@A@(~D*~(C*~B)))"),
    .INIT(32'haa65559a))
    _al_u259 (
    .a(_al_u177_o),
    .b(_al_u159_o),
    .c(_al_u163_o),
    .d(_al_u219_o),
    .e(_al_u212_o),
    .o(_al_u259_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~D*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)))"),
    .INIT(32'haa22aa0a))
    _al_u260 (
    .a(_al_u150_o),
    .b(_al_u205_o),
    .c(_al_u208_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u260_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@A@(C*~(~D*B)))"),
    .INIT(32'h5a9aa565))
    _al_u261 (
    .a(_al_u195_o),
    .b(_al_u260_o),
    .c(_al_u214_o),
    .d(_al_u202_o),
    .e(_al_u212_o),
    .o(_al_u261_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u262 (
    .a(_al_u71_o),
    .b(_al_u74_o),
    .c(exp_diff[2]),
    .d(exp_diff[3]),
    .o(_al_u262_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h530f))
    _al_u263 (
    .a(_al_u101_o),
    .b(_al_u68_o),
    .c(_al_u262_o),
    .d(exp_diff[3]),
    .o(_al_u263_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(~C*~(B*~(~D*~A))))"),
    .INIT(32'hfcf80307))
    _al_u264 (
    .a(_al_u263_o),
    .b(_al_u227_o),
    .c(_al_u229_o),
    .d(_al_u118_o),
    .e(_al_u212_o),
    .o(_al_u264_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~B*A*(E@D))"),
    .INIT(32'h00020200))
    _al_u265 (
    .a(\ADD02/ADD01/ADD02/p1_lutinv ),
    .b(_al_u259_o),
    .c(_al_u261_o),
    .d(_al_u264_o),
    .e(_al_u225_o),
    .o(_al_u265_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~D*~B*A))"),
    .INIT(16'hf0d0))
    _al_u266 (
    .a(_al_u131_o),
    .b(_al_u147_o),
    .c(_al_u134_o),
    .d(_al_u118_o),
    .o(_al_u266_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D)*~((~C*~B))+~A*D*~((~C*~B))+~(~A)*D*(~C*~B)+~A*D*(~C*~B))"),
    .INIT(16'h5754))
    _al_u267 (
    .a(_al_u266_o),
    .b(_al_u119_o),
    .c(_al_u151_o),
    .d(_al_u212_o),
    .o(\ADD02/ADD01/ADD01/c0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u268 (
    .a(_al_u245_o),
    .b(_al_u246_o),
    .o(_al_u268_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(A)*~(D)+C*A*~(D)+~(C)*A*D+C*A*D))"),
    .INIT(16'h440c))
    _al_u269 (
    .a(_al_u268_o),
    .b(_al_u132_o),
    .c(_al_u248_o),
    .d(exp_diff[2]),
    .o(_al_u269_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u270 (
    .a(_al_u64_o),
    .b(n1[4]),
    .c(n1[3]),
    .o(n106_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h717d))
    _al_u271 (
    .a(n106_lutinv),
    .b(_al_u67_o),
    .c(_al_u64_o),
    .d(n1[2]),
    .o(_al_u271_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u272 (
    .a(_al_u253_o),
    .b(_al_u271_o),
    .c(exp_diff[2]),
    .d(exp_diff[3]),
    .o(_al_u272_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u273 (
    .a(_al_u249_o),
    .b(_al_u251_o),
    .c(_al_u272_o),
    .d(exp_diff[3]),
    .o(_al_u273_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u274 (
    .a(_al_u103_o),
    .b(n1[1]),
    .o(_al_u274_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(C*~(~A*~(~E*~B))))"),
    .INIT(32'h005f004f))
    _al_u275 (
    .a(_al_u269_o),
    .b(_al_u273_o),
    .c(_al_u131_o),
    .d(_al_u274_o),
    .e(_al_u118_o),
    .o(_al_u275_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u276 (
    .a(_al_u64_o),
    .b(n2[4]),
    .c(n2[3]),
    .o(n238_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u277 (
    .a(_al_u64_o),
    .b(n2[2]),
    .c(n2[1]),
    .o(_al_u277_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u278 (
    .a(n238_lutinv),
    .b(_al_u277_o),
    .c(_al_u67_o),
    .o(_al_u278_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ac))
    _al_u279 (
    .a(_al_u240_o),
    .b(_al_u278_o),
    .c(exp_diff[2]),
    .d(exp_diff[3]),
    .o(_al_u279_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hacf0))
    _al_u280 (
    .a(_al_u236_o),
    .b(_al_u237_o),
    .c(_al_u279_o),
    .d(exp_diff[3]),
    .o(_al_u280_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(A*~((~C*~B))*~(E)+A*(~C*~B)*~(E)+~(A)*(~C*~B)*E+A*(~C*~B)*E))"),
    .INIT(32'h00fc0055))
    _al_u281 (
    .a(_al_u235_o),
    .b(_al_u232_o),
    .c(_al_u233_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u281_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u282 (
    .a(_al_u103_o),
    .b(n2[1]),
    .o(_al_u282_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(C*(~A*~(B)*~(E)+~A*B*~(E)+~(~A)*B*E+~A*B*E)))"),
    .INIT(32'h003f00af))
    _al_u283 (
    .a(_al_u280_o),
    .b(_al_u281_o),
    .c(_al_u116_o),
    .d(_al_u282_o),
    .e(_al_u118_o),
    .o(_al_u283_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~((D@C))+A*~(B)*~((D@C))+A*B*~((D@C))+A*~(B)*(D@C))"),
    .INIT(16'hb22b))
    _al_u284 (
    .a(\ADD02/ADD01/ADD01/c0_lutinv ),
    .b(_al_u275_o),
    .c(_al_u283_o),
    .d(_al_u212_o),
    .o(_al_u284_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h503f))
    _al_u285 (
    .a(_al_u154_o),
    .b(_al_u156_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u285_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h0123))
    _al_u286 (
    .a(exp_diff[1]),
    .b(exp_diff[3]),
    .c(n107_lutinv),
    .d(n105_lutinv),
    .o(_al_u286_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~(~D*~C)*~(B)*~(A)+~(~D*~C)*B*~(A)+~(~(~D*~C))*B*A+~(~D*~C)*B*A))"),
    .INIT(32'h00002227))
    _al_u287 (
    .a(_al_u285_o),
    .b(_al_u286_o),
    .c(_al_u158_o),
    .d(exp_diff[3]),
    .e(_al_u118_o),
    .o(_al_u287_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(~C*~(B)*~(D)+~C*B*~(D)+~(~C)*B*D+~C*B*D))"),
    .INIT(16'h880a))
    _al_u288 (
    .a(_al_u132_o),
    .b(_al_u160_o),
    .c(_al_u153_o),
    .d(exp_diff[2]),
    .o(_al_u288_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*~D)*~(C*~(~B*~A)))"),
    .INIT(32'h1f001f1f))
    _al_u289 (
    .a(_al_u287_o),
    .b(_al_u288_o),
    .c(_al_u131_o),
    .d(_al_u103_o),
    .e(n1[2]),
    .o(_al_u289_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u290 (
    .a(_al_u201_o),
    .b(_al_u205_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u290_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5135))
    _al_u291 (
    .a(n104_lutinv),
    .b(n106_lutinv),
    .c(_al_u67_o),
    .d(_al_u64_o),
    .o(_al_u291_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D)))"),
    .INIT(32'h0000fafc))
    _al_u292 (
    .a(_al_u208_o),
    .b(_al_u291_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .e(_al_u118_o),
    .o(_al_u292_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u293 (
    .a(_al_u121_o),
    .b(_al_u64_o),
    .o(n86_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u294 (
    .a(n86_lutinv),
    .b(_al_u93_o),
    .c(_al_u67_o),
    .o(_al_u294_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~C*~(~A*~(~D*~B))))"),
    .INIT(32'hf5f40000))
    _al_u295 (
    .a(_al_u294_o),
    .b(_al_u198_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .e(_al_u118_o),
    .o(_al_u295_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u296 (
    .a(_al_u103_o),
    .b(n1[3]),
    .o(_al_u296_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*~C*~(B*~A)))"),
    .INIT(32'h0000f4ff))
    _al_u297 (
    .a(_al_u290_o),
    .b(_al_u292_o),
    .c(_al_u295_o),
    .d(_al_u131_o),
    .e(_al_u296_o),
    .o(_al_u297_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u298 (
    .a(_al_u183_o),
    .b(_al_u187_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u298_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u299 (
    .a(n236_lutinv),
    .b(n238_lutinv),
    .c(_al_u67_o),
    .o(_al_u299_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)))"),
    .INIT(32'h0000faf3))
    _al_u300 (
    .a(_al_u190_o),
    .b(_al_u299_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .e(_al_u118_o),
    .o(_al_u300_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~C*~(~A*~(~D*~B))))"),
    .INIT(32'hf5f40000))
    _al_u301 (
    .a(_al_u294_o),
    .b(_al_u180_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .e(_al_u118_o),
    .o(_al_u301_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u302 (
    .a(_al_u103_o),
    .b(n2[3]),
    .o(_al_u302_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*~C*~(B*~A)))"),
    .INIT(32'h0000f4ff))
    _al_u303 (
    .a(_al_u298_o),
    .b(_al_u300_o),
    .c(_al_u301_o),
    .d(_al_u116_o),
    .e(_al_u302_o),
    .o(_al_u303_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h5030))
    _al_u304 (
    .a(_al_u173_o),
    .b(_al_u170_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u304_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u305 (
    .a(n237_lutinv),
    .b(n239_lutinv),
    .c(_al_u67_o),
    .o(_al_u305_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)))"),
    .INIT(32'h0000faf3))
    _al_u306 (
    .a(_al_u175_o),
    .b(_al_u305_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .e(_al_u118_o),
    .o(_al_u306_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u307 (
    .a(_al_u96_o),
    .b(_al_u67_o),
    .o(_al_u307_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~C*(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D)))"),
    .INIT(32'hf5fc0000))
    _al_u308 (
    .a(_al_u307_o),
    .b(_al_u172_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .e(_al_u118_o),
    .o(_al_u308_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u309 (
    .a(_al_u103_o),
    .b(n2[2]),
    .o(_al_u309_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*~C*~(B*~A)))"),
    .INIT(32'h0000f4ff))
    _al_u310 (
    .a(_al_u304_o),
    .b(_al_u306_o),
    .c(_al_u308_o),
    .d(_al_u116_o),
    .e(_al_u309_o),
    .o(_al_u310_o));
  AL_MAP_LUT5 #(
    .EQN("(A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*B*C*D*E)"),
    .INIT(32'h8ecffce8))
    _al_u311 (
    .a(_al_u289_o),
    .b(_al_u297_o),
    .c(_al_u303_o),
    .d(_al_u310_o),
    .e(_al_u212_o),
    .o(_al_u311_o));
  AL_MAP_LUT5 #(
    .EQN("(~((C@B))*~((D@A))*~(E)+(C@B)*~((D@A))*~(E)+~((C@B))*(D@A)*~(E)+(C@B)*~((D@A))*E+~((C@B))*(D@A)*E+(C@B)*(D@A)*E)"),
    .INIT(32'h7dbeebd7))
    _al_u312 (
    .a(_al_u289_o),
    .b(_al_u297_o),
    .c(_al_u303_o),
    .d(_al_u310_o),
    .e(_al_u212_o),
    .o(_al_u312_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B*~(D*~(~E*C))))"),
    .INIT(32'haa222a22))
    _al_u313 (
    .a(_al_u257_o),
    .b(_al_u265_o),
    .c(_al_u284_o),
    .d(_al_u311_o),
    .e(_al_u312_o),
    .o(_al_u313_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfff055cc))
    _al_u314 (
    .a(_al_u124_o),
    .b(_al_u142_o),
    .c(_al_u127_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u314_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u315 (
    .a(_al_u314_o),
    .b(_al_u150_o),
    .c(_al_u103_o),
    .d(n1[12]),
    .o(_al_u315_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hffcc55f0))
    _al_u316 (
    .a(_al_u98_o),
    .b(_al_u101_o),
    .c(_al_u68_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u316_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u317 (
    .a(_al_u118_o),
    .b(_al_u110_o),
    .c(_al_u112_o),
    .d(_al_u115_o),
    .o(_al_u317_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u318 (
    .a(_al_u316_o),
    .b(_al_u317_o),
    .c(_al_u103_o),
    .d(n2[12]),
    .o(_al_u318_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    _al_u319 (
    .a(_al_u315_o),
    .b(_al_u318_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD02/ADD02/g0 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hffccaaf0))
    _al_u320 (
    .a(_al_u268_o),
    .b(_al_u248_o),
    .c(_al_u249_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u320_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u321 (
    .a(_al_u148_o),
    .b(_al_u103_o),
    .o(_al_u321_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C))"),
    .INIT(16'h00ac))
    _al_u322 (
    .a(_al_u149_o),
    .b(_al_u116_o),
    .c(_al_u321_o),
    .d(_al_u118_o),
    .o(u194_sel_is_0_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((B*~A))*~(C)+D*(B*~A)*~(C)+~(D)*(B*~A)*C+D*(B*~A)*C)"),
    .INIT(16'hb0bf))
    _al_u323 (
    .a(_al_u320_o),
    .b(u194_sel_is_0_o),
    .c(_al_u103_o),
    .d(n1[13]),
    .o(_al_u323_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u324 (
    .a(_al_u232_o),
    .b(_al_u233_o),
    .o(_al_u324_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hffccaaf0))
    _al_u325 (
    .a(_al_u324_o),
    .b(_al_u235_o),
    .c(_al_u236_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u325_o));
  AL_MAP_LUT5 #(
    .EQN("(D@~((B*~A)*~(E)*~(C)+(B*~A)*E*~(C)+~((B*~A))*E*C+(B*~A)*E*C))"),
    .INIT(32'hf40b04fb))
    _al_u326 (
    .a(_al_u325_o),
    .b(u194_sel_is_0_o),
    .c(_al_u103_o),
    .d(_al_u212_o),
    .e(n2[13]),
    .o(_al_u326_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*B*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'hd4))
    _al_u327 (
    .a(\ADD02/ADD02/ADD02/g0 ),
    .b(_al_u323_o),
    .c(_al_u326_o),
    .o(_al_u327_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hffcc55f0))
    _al_u328 (
    .a(_al_u307_o),
    .b(_al_u172_o),
    .c(_al_u173_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u328_o));
  AL_MAP_LUT4 #(
    .EQN("~((~B*A)*~(D)*~(C)+(~B*A)*D*~(C)+~((~B*A))*D*C+(~B*A)*D*C)"),
    .INIT(16'h0dfd))
    _al_u329 (
    .a(u194_sel_is_0_o),
    .b(_al_u328_o),
    .c(_al_u103_o),
    .d(n2[14]),
    .o(_al_u329_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u330 (
    .a(_al_u329_o),
    .b(_al_u212_o),
    .o(_al_u330_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hffcc55f0))
    _al_u331 (
    .a(_al_u160_o),
    .b(_al_u153_o),
    .c(_al_u154_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u331_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u332 (
    .a(_al_u331_o),
    .b(_al_u150_o),
    .c(_al_u103_o),
    .d(n1[14]),
    .o(_al_u332_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u333 (
    .a(_al_u330_o),
    .b(_al_u332_o),
    .o(\ADD02/ADD02/ADD02/p2_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u334 (
    .a(_al_u198_o),
    .b(_al_u201_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u334_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u335 (
    .a(exp_diff[3]),
    .b(n198_lutinv),
    .o(_al_u335_o));
  AL_MAP_LUT5 #(
    .EQN("~(E*~((~C*~B*A))*~(D)+E*(~C*~B*A)*~(D)+~(E)*(~C*~B*A)*D+E*(~C*~B*A)*D)"),
    .INIT(32'hfd00fdff))
    _al_u336 (
    .a(u194_sel_is_0_o),
    .b(_al_u334_o),
    .c(_al_u335_o),
    .d(_al_u103_o),
    .e(n1[15]),
    .o(_al_u336_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u337 (
    .a(_al_u180_o),
    .b(_al_u183_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u337_o));
  AL_MAP_LUT5 #(
    .EQN("~((~C*~B*A)*~(E)*~(D)+(~C*~B*A)*E*~(D)+~((~C*~B*A))*E*D+(~C*~B*A)*E*D)"),
    .INIT(32'h00fdfffd))
    _al_u338 (
    .a(u194_sel_is_0_o),
    .b(_al_u337_o),
    .c(_al_u335_o),
    .d(_al_u103_o),
    .e(n2[15]),
    .o(_al_u338_o));
  AL_MAP_LUT5 #(
    .EQN("(A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hbb2beee8))
    _al_u339 (
    .a(_al_u336_o),
    .b(_al_u338_o),
    .c(_al_u329_o),
    .d(_al_u332_o),
    .e(_al_u212_o),
    .o(_al_u339_o));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u340 (
    .a(_al_u336_o),
    .b(_al_u338_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD02/ADD02/p3_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*B*~A))"),
    .INIT(16'hb0f0))
    _al_u341 (
    .a(_al_u327_o),
    .b(\ADD02/ADD02/ADD02/p2_lutinv ),
    .c(_al_u339_o),
    .d(\ADD02/ADD02/ADD02/p3_lutinv ),
    .o(_al_u341_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u342 (
    .a(_al_u323_o),
    .b(_al_u326_o),
    .o(\ADD02/ADD02/ADD02/p1_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u343 (
    .a(_al_u315_o),
    .b(_al_u318_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD02/ADD02/p0_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u344 (
    .a(\ADD02/ADD02/ADD02/p2_lutinv ),
    .b(\ADD02/ADD02/ADD02/p1_lutinv ),
    .c(\ADD02/ADD02/ADD02/p3_lutinv ),
    .d(\ADD02/ADD02/ADD02/p0_lutinv ),
    .o(_al_u344_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~((~C*~B))*~(D)*~(E)+A*~((~C*~B))*~(D)*~(E)+~(A)*(~C*~B)*~(D)*~(E)+A*(~C*~B)*~(D)*~(E)+~(A)*~((~C*~B))*D*~(E)+~(A)*(~C*~B)*D*~(E)+~(A)*~((~C*~B))*D*E+A*~((~C*~B))*D*E)"),
    .INIT(32'hfc0055ff))
    _al_u345 (
    .a(_al_u235_o),
    .b(_al_u232_o),
    .c(_al_u233_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u345_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*A*~(C*~B))"),
    .INIT(32'h0000008a))
    _al_u346 (
    .a(_al_u168_o),
    .b(_al_u162_o),
    .c(_al_u237_o),
    .d(_al_u118_o),
    .e(_al_u103_o),
    .o(_al_u346_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u347 (
    .a(_al_u236_o),
    .b(exp_diff[3]),
    .o(_al_u347_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u348 (
    .a(_al_u103_o),
    .b(n2[9]),
    .o(_al_u348_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~(B*~(~C*~A))))"),
    .INIT(32'hffc80037))
    _al_u349 (
    .a(_al_u345_o),
    .b(_al_u346_o),
    .c(_al_u347_o),
    .d(_al_u348_o),
    .e(_al_u212_o),
    .o(_al_u349_o));
  AL_MAP_LUT5 #(
    .EQN("(D*(C*~((~B*~A))*~(E)+C*(~B*~A)*~(E)+~(C)*(~B*~A)*E+C*(~B*~A)*E))"),
    .INIT(32'h1100f000))
    _al_u350 (
    .a(_al_u245_o),
    .b(_al_u246_o),
    .c(_al_u248_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u350_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u351 (
    .a(_al_u249_o),
    .b(_al_u251_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u351_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*~D)*~(C*~B*~A))"),
    .INIT(32'hef00efef))
    _al_u352 (
    .a(_al_u350_o),
    .b(_al_u351_o),
    .c(_al_u150_o),
    .d(_al_u103_o),
    .e(n1[9]),
    .o(_al_u352_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u353 (
    .a(_al_u142_o),
    .b(_al_u145_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u353_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u354 (
    .a(_al_u103_o),
    .b(n1[8]),
    .o(_al_u354_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(C*~B*~(E*A)))"),
    .INIT(32'h00ef00cf))
    _al_u355 (
    .a(_al_u128_o),
    .b(_al_u353_o),
    .c(_al_u150_o),
    .d(_al_u354_o),
    .e(exp_diff[3]),
    .o(_al_u355_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u356 (
    .a(_al_u68_o),
    .b(_al_u71_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u356_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C))"),
    .INIT(16'h005c))
    _al_u357 (
    .a(_al_u98_o),
    .b(_al_u101_o),
    .c(exp_diff[2]),
    .d(\C023/outtemp [3]),
    .o(_al_u357_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u358 (
    .a(_al_u103_o),
    .b(n2[8]),
    .o(_al_u358_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~(C*~B*~A)))"),
    .INIT(32'hff1000ef))
    _al_u359 (
    .a(_al_u356_o),
    .b(_al_u357_o),
    .c(_al_u317_o),
    .d(_al_u358_o),
    .e(_al_u212_o),
    .o(_al_u359_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~((~D*~C))+~(A)*B*~((~D*~C))+A*B*~((~D*~C))+A*B*(~D*~C))"),
    .INIT(16'heee8))
    _al_u360 (
    .a(_al_u349_o),
    .b(_al_u352_o),
    .c(_al_u355_o),
    .d(_al_u359_o),
    .o(_al_u360_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u361 (
    .a(_al_u183_o),
    .b(_al_u187_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u361_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~A*~((~E*C))*~(B)+~A*(~E*C)*~(B)+~(~A)*(~E*C)*B+~A*(~E*C)*B))"),
    .INIT(32'h00ee002e))
    _al_u362 (
    .a(_al_u180_o),
    .b(exp_diff[2]),
    .c(n86_lutinv),
    .d(\C023/outtemp [3]),
    .e(_al_u67_o),
    .o(_al_u362_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u363 (
    .a(_al_u103_o),
    .b(n2[11]),
    .o(_al_u363_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~(C*~B*~A)))"),
    .INIT(32'hff1000ef))
    _al_u364 (
    .a(_al_u361_o),
    .b(_al_u362_o),
    .c(_al_u317_o),
    .d(_al_u363_o),
    .e(_al_u212_o),
    .o(_al_u364_o));
  AL_MAP_LUT4 #(
    .EQN("~(~A*~((~D*C))*~(B)+~A*(~D*C)*~(B)+~(~A)*(~D*C)*B+~A*(~D*C)*B)"),
    .INIT(16'hee2e))
    _al_u365 (
    .a(_al_u198_o),
    .b(exp_diff[2]),
    .c(n86_lutinv),
    .d(_al_u67_o),
    .o(_al_u365_o));
  AL_MAP_LUT5 #(
    .EQN("~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*~(A)*~(D)+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*~(D)+~((C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E))*A*D+(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)*A*D)"),
    .INIT(32'h5533550f))
    _al_u366 (
    .a(_al_u365_o),
    .b(_al_u201_o),
    .c(_al_u205_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u366_o));
  AL_MAP_LUT5 #(
    .EQN("(A@(~(E*~D)*~(C*B)))"),
    .INIT(32'h95aa9595))
    _al_u367 (
    .a(_al_u364_o),
    .b(_al_u366_o),
    .c(_al_u150_o),
    .d(_al_u103_o),
    .e(n1[11]),
    .o(\ADD02/ADD02/ADD01/p3_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~D*(C*~(B)*~(E)+C*B*~(E)+~(C)*B*E+C*B*E)))"),
    .INIT(32'haa22aa0a))
    _al_u368 (
    .a(_al_u150_o),
    .b(_al_u154_o),
    .c(_al_u156_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u368_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(16'h50c0))
    _al_u369 (
    .a(_al_u160_o),
    .b(_al_u153_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u369_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(~B*A))"),
    .INIT(16'hd0dd))
    _al_u370 (
    .a(_al_u368_o),
    .b(_al_u369_o),
    .c(_al_u103_o),
    .d(n1[10]),
    .o(_al_u370_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(A)*~(D)+~B*A*~(D)+~(~B)*A*D+~B*A*D))"),
    .INIT(16'h50c0))
    _al_u371 (
    .a(_al_u307_o),
    .b(_al_u172_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u371_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*(B*~(A)*~(D)+B*A*~(D)+~(B)*A*D+B*A*D))"),
    .INIT(16'h0a0c))
    _al_u372 (
    .a(_al_u173_o),
    .b(_al_u170_o),
    .c(exp_diff[3]),
    .d(exp_diff[2]),
    .o(_al_u372_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u373 (
    .a(_al_u103_o),
    .b(n2[10]),
    .o(_al_u373_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~(C*~B*~A)))"),
    .INIT(32'hff1000ef))
    _al_u374 (
    .a(_al_u371_o),
    .b(_al_u372_o),
    .c(_al_u317_o),
    .d(_al_u373_o),
    .e(_al_u212_o),
    .o(_al_u374_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~((~(A)*~(C)*~(D)+A*~(C)*~(D)+~(A)*C*~(D)+~(A)*~(C)*D))*~(B)+~E*(~(A)*~(C)*~(D)+A*~(C)*~(D)+~(A)*C*~(D)+~(A)*~(C)*D)*~(B)+~(~E)*(~(A)*~(C)*~(D)+A*~(C)*~(D)+~(A)*C*~(D)+~(A)*~(C)*D)*B+~E*(~(A)*~(C)*~(D)+A*~(C)*~(D)+~(A)*C*~(D)+~(A)*~(C)*D)*B)"),
    .INIT(32'h044c377f))
    _al_u375 (
    .a(_al_u360_o),
    .b(\ADD02/ADD02/ADD01/p3_lutinv ),
    .c(_al_u370_o),
    .d(_al_u374_o),
    .e(_al_u364_o),
    .o(_al_u375_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u376 (
    .a(_al_u349_o),
    .b(_al_u352_o),
    .o(\ADD02/ADD02/ADD01/p1_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u377 (
    .a(_al_u128_o),
    .b(_al_u150_o),
    .c(exp_diff[3]),
    .o(_al_u377_o));
  AL_MAP_LUT5 #(
    .EQN("(A@(~(E*~D)*~(~C*B)))"),
    .INIT(32'h59aa5959))
    _al_u378 (
    .a(_al_u359_o),
    .b(_al_u377_o),
    .c(_al_u353_o),
    .d(_al_u103_o),
    .e(n1[8]),
    .o(\ADD02/ADD02/ADD01/p0_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*(E@D))"),
    .INIT(32'h00808000))
    _al_u379 (
    .a(\ADD02/ADD02/ADD01/p1_lutinv ),
    .b(\ADD02/ADD02/ADD01/p0_lutinv ),
    .c(\ADD02/ADD02/ADD01/p3_lutinv ),
    .d(_al_u370_o),
    .e(_al_u374_o),
    .o(\ADD02/ADD02/ADD01/n20 ));
  AL_MAP_LUT5 #(
    .EQN("(B*~(C*~(~D*~(E*~A))))"),
    .INIT(32'h0c8c0ccc))
    _al_u380 (
    .a(_al_u313_o),
    .b(_al_u341_o),
    .c(_al_u344_o),
    .d(_al_u375_o),
    .e(\ADD02/ADD02/ADD01/n20 ),
    .o(_al_u380_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*~(B)*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'hd3))
    _al_u381 (
    .a(_al_u103_o),
    .b(_al_u121_o),
    .c(_al_u212_o),
    .o(_al_u381_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~E*D)*~(C*~B*A))"),
    .INIT(32'hdfdf00df))
    _al_u382 (
    .a(u194_sel_is_0_o),
    .b(exp_diff[3]),
    .c(n198_lutinv),
    .d(_al_u103_o),
    .e(_al_u121_o),
    .o(_al_u382_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(D@A))"),
    .INIT(16'h0201))
    _al_u383 (
    .a(_al_u382_o),
    .b(_al_u103_o),
    .c(_al_u121_o),
    .d(_al_u212_o),
    .o(\ADD02/ADD03/ADD02/g3 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u384 (
    .a(_al_u317_o),
    .b(exp_diff[3]),
    .o(_al_u384_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u385 (
    .a(_al_u384_o),
    .b(_al_u165_o),
    .c(_al_u103_o),
    .d(n2[22]),
    .o(_al_u385_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*~D)*~(~C*B*A))"),
    .INIT(32'hf700f7f7))
    _al_u386 (
    .a(_al_u150_o),
    .b(_al_u160_o),
    .c(_al_u162_o),
    .d(_al_u103_o),
    .e(n1[22]),
    .o(_al_u386_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C@A))"),
    .INIT(8'h21))
    _al_u387 (
    .a(_al_u385_o),
    .b(_al_u386_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD03/ADD02/g2 ));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u388 (
    .a(_al_u385_o),
    .b(_al_u386_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD03/ADD02/p2_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~(E*~D)*~(~C*B*~A))"),
    .INIT(32'hfb00fbfb))
    _al_u389 (
    .a(_al_u268_o),
    .b(_al_u150_o),
    .c(_al_u162_o),
    .d(_al_u103_o),
    .e(n1[21]),
    .o(_al_u389_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D)*~(~C*B*~A))"),
    .INIT(32'h00fbfbfb))
    _al_u390 (
    .a(_al_u324_o),
    .b(_al_u317_o),
    .c(_al_u162_o),
    .d(_al_u103_o),
    .e(n2[21]),
    .o(_al_u390_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    _al_u391 (
    .a(_al_u389_o),
    .b(_al_u390_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD03/ADD02/g1 ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~C*~B*~(E*D)))"),
    .INIT(32'haaa8a8a8))
    _al_u392 (
    .a(_al_u381_o),
    .b(\ADD02/ADD03/ADD02/g3 ),
    .c(\ADD02/ADD03/ADD02/g2 ),
    .d(\ADD02/ADD03/ADD02/p2_lutinv ),
    .e(\ADD02/ADD03/ADD02/g1 ),
    .o(\ADD02/ADD03/ADD02/n16_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u393 (
    .a(_al_u381_o),
    .b(\ADD02/ADD03/ADD02/g3 ),
    .o(\ADD02/ADD03/ADD02/p3_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u394 (
    .a(_al_u317_o),
    .b(_al_u98_o),
    .c(_al_u162_o),
    .o(_al_u394_o));
  AL_MAP_LUT4 #(
    .EQN("(C@(~A*~(D*B)))"),
    .INIT(16'he1a5))
    _al_u395 (
    .a(_al_u394_o),
    .b(_al_u103_o),
    .c(_al_u212_o),
    .d(n2[20]),
    .o(_al_u395_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*~D)*~(~C*B*A))"),
    .INIT(32'hf700f7f7))
    _al_u396 (
    .a(_al_u150_o),
    .b(_al_u124_o),
    .c(_al_u162_o),
    .d(_al_u103_o),
    .e(n1[20]),
    .o(_al_u396_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u397 (
    .a(_al_u395_o),
    .b(_al_u396_o),
    .o(\ADD02/ADD03/ADD02/g0 ));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u398 (
    .a(_al_u389_o),
    .b(_al_u390_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD03/ADD02/p1_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u399 (
    .a(\ADD02/ADD03/ADD02/g0 ),
    .b(\ADD02/ADD03/ADD02/p1_lutinv ),
    .o(\ADD02/ADD03/ADD02/n1 ));
  AL_MAP_LUT5 #(
    .EQN("(E*~A*~(D*C*B))"),
    .INIT(32'h15550000))
    _al_u400 (
    .a(\ADD02/ADD03/ADD02/n16_lutinv ),
    .b(\ADD02/ADD03/ADD02/p3_lutinv ),
    .c(\ADD02/ADD03/ADD02/n1 ),
    .d(\ADD02/ADD03/ADD02/p2_lutinv ),
    .e(_al_u212_o),
    .o(_al_u400_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u401 (
    .a(_al_u149_o),
    .b(_al_u321_o),
    .c(exp_diff[3]),
    .d(_al_u118_o),
    .o(_al_u401_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(~B*A))"),
    .INIT(16'hd0dd))
    _al_u402 (
    .a(_al_u401_o),
    .b(_al_u128_o),
    .c(_al_u103_o),
    .d(n1[16]),
    .o(_al_u402_o));
  AL_MAP_LUT4 #(
    .EQN("~((B*A)*~(D)*~(C)+(B*A)*D*~(C)+~((B*A))*D*C+(B*A)*D*C)"),
    .INIT(16'h07f7))
    _al_u403 (
    .a(u194_sel_is_0_o),
    .b(_al_u102_o),
    .c(_al_u103_o),
    .d(n2[16]),
    .o(_al_u403_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u404 (
    .a(_al_u103_o),
    .b(n1[17]),
    .o(_al_u404_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(A*~(D*~(B)*~(E)+D*B*~(E)+~(D)*B*E+D*B*E)))"),
    .INIT(32'h0d0d0f05))
    _al_u405 (
    .a(_al_u401_o),
    .b(_al_u268_o),
    .c(_al_u404_o),
    .d(_al_u248_o),
    .e(exp_diff[2]),
    .o(_al_u405_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u406 (
    .a(_al_u281_o),
    .b(_al_u317_o),
    .c(_al_u103_o),
    .d(n2[17]),
    .o(_al_u406_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*(~(B)*(D@C)*~(E)+B*~((D@C))*E))"),
    .INIT(32'h40040110))
    _al_u407 (
    .a(_al_u402_o),
    .b(_al_u403_o),
    .c(_al_u405_o),
    .d(_al_u406_o),
    .e(_al_u212_o),
    .o(_al_u407_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C@B))"),
    .INIT(8'h41))
    _al_u408 (
    .a(_al_u405_o),
    .b(_al_u406_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD03/ADD01/g1 ));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'ha3))
    _al_u409 (
    .a(_al_u160_o),
    .b(_al_u153_o),
    .c(exp_diff[2]),
    .o(_al_u409_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*A))"),
    .INIT(16'h7077))
    _al_u410 (
    .a(_al_u401_o),
    .b(_al_u409_o),
    .c(_al_u103_o),
    .d(n1[18]),
    .o(_al_u410_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'ha3))
    _al_u411 (
    .a(_al_u307_o),
    .b(_al_u172_o),
    .c(exp_diff[2]),
    .o(_al_u411_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u412 (
    .a(_al_u384_o),
    .b(_al_u411_o),
    .c(_al_u103_o),
    .d(n2[18]),
    .o(_al_u412_o));
  AL_MAP_LUT5 #(
    .EQN("(~((~B*~A))*~(C)*~((E@D))+(~B*~A)*~(C)*~((E@D))+~((~B*~A))*C*~((E@D))+~((~B*~A))*~(C)*(E@D))"),
    .INIT(32'hef0e0eef))
    _al_u413 (
    .a(_al_u407_o),
    .b(\ADD02/ADD03/ADD01/g1 ),
    .c(_al_u410_o),
    .d(_al_u412_o),
    .e(_al_u212_o),
    .o(_al_u413_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*~B))"),
    .INIT(8'h54))
    _al_u414 (
    .a(_al_u294_o),
    .b(_al_u180_o),
    .c(exp_diff[2]),
    .o(_al_u414_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(~B*A))"),
    .INIT(16'h0ddd))
    _al_u415 (
    .a(_al_u384_o),
    .b(_al_u414_o),
    .c(_al_u103_o),
    .d(n2[19]),
    .o(_al_u415_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*~D)*~(~C*~B*A))"),
    .INIT(32'hfd00fdfd))
    _al_u416 (
    .a(_al_u150_o),
    .b(_al_u365_o),
    .c(exp_diff[3]),
    .d(_al_u103_o),
    .e(n1[19]),
    .o(_al_u416_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(C)*~((D@B))+A*~(C)*~((D@B))+A*C*~((D@B))+A*~(C)*(D@B))"),
    .INIT(16'h8e2b))
    _al_u417 (
    .a(_al_u413_o),
    .b(_al_u415_o),
    .c(_al_u416_o),
    .d(_al_u212_o),
    .o(_al_u417_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u418 (
    .a(_al_u395_o),
    .b(_al_u396_o),
    .o(\ADD02/ADD03/ADD02/p0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u419 (
    .a(\ADD02/ADD03/ADD02/p0_lutinv ),
    .b(\ADD02/ADD03/ADD02/p1_lutinv ),
    .o(\ADD02/ADD03/ADD02/n3 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u420 (
    .a(\ADD02/ADD03/ADD02/p3_lutinv ),
    .b(\ADD02/ADD03/ADD02/n3 ),
    .c(\ADD02/ADD03/ADD02/p2_lutinv ),
    .o(_al_u420_o));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u421 (
    .a(_al_u410_o),
    .b(_al_u412_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD03/ADD01/p2_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u422 (
    .a(_al_u402_o),
    .b(_al_u403_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD03/ADD01/p0_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u423 (
    .a(_al_u405_o),
    .b(_al_u406_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD03/ADD01/p1_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u424 (
    .a(_al_u415_o),
    .b(_al_u416_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD03/ADD01/p3_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u425 (
    .a(\ADD02/ADD03/ADD01/p2_lutinv ),
    .b(\ADD02/ADD03/ADD01/p0_lutinv ),
    .c(\ADD02/ADD03/ADD01/p1_lutinv ),
    .d(\ADD02/ADD03/ADD01/p3_lutinv ),
    .o(_al_u425_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(D*~(~C*~(E*~A))))"),
    .INIT(32'h08cc0ccc))
    _al_u426 (
    .a(_al_u380_o),
    .b(_al_u400_o),
    .c(_al_u417_o),
    .d(_al_u420_o),
    .e(_al_u425_o),
    .o(_al_u426_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u427 (
    .a(_al_u119_o),
    .b(_al_u151_o),
    .o(_al_u427_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~((C@B))*~(D)*~(E)+A*~((C@B))*~(D)*~(E)+A*(C@B)*~(D)*~(E)+~(A)*~((C@B))*D*~(E)+~(A)*(C@B)*D*~(E)+A*(C@B)*D*~(E)+A*~((C@B))*~(D)*E+~(A)*(C@B)*~(D)*E+A*(C@B)*~(D)*E+~(A)*~((C@B))*D*E+~(A)*(C@B)*D*E+A*(C@B)*D*E)"),
    .INIT(32'h7dbe7deb))
    _al_u428 (
    .a(_al_u427_o),
    .b(_al_u275_o),
    .c(_al_u283_o),
    .d(_al_u266_o),
    .e(_al_u212_o),
    .o(_al_u428_o));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u429 (
    .a(_al_u289_o),
    .b(_al_u310_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD01/ADD01/p2_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u430 (
    .a(_al_u297_o),
    .b(_al_u303_o),
    .c(_al_u212_o),
    .o(\ADD02/ADD01/ADD01/p3_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u431 (
    .a(_al_u428_o),
    .b(\ADD02/ADD01/ADD01/p2_lutinv ),
    .c(\ADD02/ADD01/ADD01/p3_lutinv ),
    .o(_al_u431_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u432 (
    .a(_al_u264_o),
    .b(_al_u225_o),
    .o(_al_u432_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*~B*A)"),
    .INIT(16'h0020))
    _al_u433 (
    .a(_al_u431_o),
    .b(_al_u432_o),
    .c(\ADD02/ADD01/ADD02/p1_lutinv ),
    .d(\ADD02/ADD01/ADD02/g0 ),
    .o(_al_u433_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u434 (
    .a(_al_u283_o),
    .b(_al_u212_o),
    .o(_al_u434_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~B*(~(C)*~(D)*~(E)+~(C)*D*~(E)+C*D*~(E)+~(C)*D*E)))"),
    .INIT(32'ha8aa88a8))
    _al_u435 (
    .a(_al_u311_o),
    .b(_al_u312_o),
    .c(_al_u434_o),
    .d(\ADD02/ADD01/ADD01/c0_lutinv ),
    .e(_al_u275_o),
    .o(_al_u435_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(~(A)*~(C)*~(D)+A*~(C)*~(D)+A*C*~(D)+A*~(C)*D)*~(E)*~(B)+~(~(A)*~(C)*~(D)+A*~(C)*~(D)+A*C*~(D)+A*~(C)*D)*E*~(B)+~(~(~(A)*~(C)*~(D)+A*~(C)*~(D)+A*C*~(D)+A*~(C)*D))*E*B+~(~(A)*~(C)*~(D)+A*~(C)*~(D)+A*C*~(D)+A*~(C)*D)*E*B)"),
    .INIT(32'h0223ceef))
    _al_u436 (
    .a(\ADD02/ADD01/ADD02/g0 ),
    .b(_al_u259_o),
    .c(_al_u244_o),
    .d(_al_u256_o),
    .e(_al_u164_o),
    .o(_al_u436_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u437 (
    .a(\ADD02/ADD01/ADD02/p1_lutinv ),
    .b(_al_u259_o),
    .o(\ADD02/ADD01/ADD02/n7 ));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u438 (
    .a(_al_u264_o),
    .b(_al_u225_o),
    .o(_al_u438_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(~B*~(~D*C*~A)))"),
    .INIT(32'hccdc3323))
    _al_u439 (
    .a(_al_u435_o),
    .b(_al_u436_o),
    .c(\ADD02/ADD01/ADD02/n7 ),
    .d(_al_u438_o),
    .e(_al_u261_o),
    .o(_al_u439_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*B*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'hd4))
    _al_u440 (
    .a(\ADD02/ADD01/ADD02/g0 ),
    .b(_al_u244_o),
    .c(_al_u256_o),
    .o(_al_u440_o));
  AL_MAP_LUT5 #(
    .EQN("(~((C@A))*~((D@B))*~(E)+(C@A)*~((D@B))*~(E)+~((C@A))*(D@B)*~(E)+(C@A)*~((D@B))*E+~((C@A))*(D@B)*E+(C@A)*(D@B)*E)"),
    .INIT(32'h7bdeedb7))
    _al_u441 (
    .a(_al_u256_o),
    .b(_al_u225_o),
    .c(_al_u243_o),
    .d(_al_u230_o),
    .e(_al_u212_o),
    .o(_al_u441_o));
  AL_MAP_LUT4 #(
    .EQN("~(D@(B*~(~C*~A)))"),
    .INIT(16'hc837))
    _al_u442 (
    .a(_al_u435_o),
    .b(_al_u440_o),
    .c(_al_u441_o),
    .d(_al_u259_o),
    .o(_al_u442_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u443 (
    .a(_al_u433_o),
    .b(_al_u439_o),
    .c(_al_u442_o),
    .d(\ADD02/ADD02/ADD01/p0_lutinv ),
    .o(_al_u443_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u444 (
    .a(\ADD02/ADD02/ADD01/p1_lutinv ),
    .b(\ADD02/ADD02/ADD01/p0_lutinv ),
    .o(\ADD02/ADD02/ADD01/n3 ));
  AL_MAP_LUT5 #(
    .EQN("(E*~(D*~(B*~(C*~A))))"),
    .INIT(32'h8cff0000))
    _al_u445 (
    .a(_al_u435_o),
    .b(_al_u257_o),
    .c(_al_u265_o),
    .d(\ADD02/ADD02/ADD01/n3 ),
    .e(_al_u360_o),
    .o(_al_u445_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u446 (
    .a(_al_u370_o),
    .b(_al_u374_o),
    .o(\ADD02/ADD02/ADD01/p2_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u447 (
    .a(_al_u445_o),
    .b(\ADD02/ADD02/ADD01/p2_lutinv ),
    .o(_al_u447_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(E*~(B*~(D*~A))))"),
    .INIT(32'h080c0f0f))
    _al_u448 (
    .a(_al_u435_o),
    .b(_al_u257_o),
    .c(_al_u375_o),
    .d(_al_u265_o),
    .e(\ADD02/ADD02/ADD01/n20 ),
    .o(_al_u448_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u449 (
    .a(_al_u448_o),
    .b(\ADD02/ADD02/ADD02/p0_lutinv ),
    .o(_al_u449_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u450 (
    .a(\ADD02/ADD02/ADD01/p1_lutinv ),
    .b(\ADD02/ADD02/ADD01/p3_lutinv ),
    .o(_al_u450_o));
  AL_MAP_LUT5 #(
    .EQN("(D@(A*~(E*C*B)))"),
    .INIT(32'hd52a55aa))
    _al_u451 (
    .a(_al_u426_o),
    .b(_al_u443_o),
    .c(_al_u447_o),
    .d(_al_u449_o),
    .e(_al_u450_o),
    .o(M_result2[12]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u452 (
    .a(_al_u355_o),
    .b(_al_u359_o),
    .o(\ADD02/ADD02/ADD01/g0 ));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(E*~(B*~(C*~A))))"),
    .INIT(32'h008c00ff))
    _al_u453 (
    .a(_al_u435_o),
    .b(_al_u257_o),
    .c(_al_u265_o),
    .d(\ADD02/ADD02/ADD01/g0 ),
    .e(\ADD02/ADD02/ADD01/p0_lutinv ),
    .o(_al_u453_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u454 (
    .a(_al_u453_o),
    .b(\ADD02/ADD02/ADD01/p1_lutinv ),
    .o(_al_u454_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(C)*~((~D*~B))+~(A)*C*~((~D*~B))+A*C*~((~D*~B))+A*C*(~D*~B))"),
    .INIT(16'hfae8))
    _al_u455 (
    .a(_al_u370_o),
    .b(_al_u349_o),
    .c(_al_u374_o),
    .d(_al_u352_o),
    .o(_al_u455_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@(C*~(D*B*~A)))"),
    .INIT(32'hb0f04f0f))
    _al_u456 (
    .a(_al_u453_o),
    .b(\ADD02/ADD02/ADD01/p2_lutinv ),
    .c(_al_u455_o),
    .d(\ADD02/ADD02/ADD01/p1_lutinv ),
    .e(\ADD02/ADD02/ADD01/p3_lutinv ),
    .o(_al_u456_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(A*~(D*C*B)))"),
    .INIT(32'hd5552aaa))
    _al_u457 (
    .a(_al_u426_o),
    .b(_al_u443_o),
    .c(_al_u447_o),
    .d(_al_u454_o),
    .e(_al_u456_o),
    .o(M_result2[11]));
  AL_MAP_LUT4 #(
    .EQN("~(C@(A*~(D*B)))"),
    .INIT(16'h2da5))
    _al_u458 (
    .a(_al_u426_o),
    .b(_al_u443_o),
    .c(_al_u447_o),
    .d(_al_u454_o),
    .o(M_result2[10]));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(E*~(C*~(D*~A))))"),
    .INIT(32'h20303333))
    _al_u459 (
    .a(_al_u448_o),
    .b(_al_u417_o),
    .c(_al_u341_o),
    .d(_al_u344_o),
    .e(_al_u425_o),
    .o(_al_u459_o));
  AL_MAP_LUT5 #(
    .EQN("~(C@(D*~A*~(E*~B)))"),
    .INIT(32'h4b0f5a0f))
    _al_u460 (
    .a(_al_u443_o),
    .b(_al_u459_o),
    .c(_al_u454_o),
    .d(_al_u400_o),
    .e(_al_u420_o),
    .o(M_result2[9]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*~B*A))"),
    .INIT(16'hdf00))
    _al_u461 (
    .a(_al_u433_o),
    .b(_al_u439_o),
    .c(_al_u442_o),
    .d(_al_u212_o),
    .o(_al_u461_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u462 (
    .a(_al_u313_o),
    .b(\ADD02/ADD02/ADD01/p0_lutinv ),
    .o(_al_u462_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u463 (
    .a(\ADD02/ADD03/ADD02/n16_lutinv ),
    .b(\ADD02/ADD03/ADD02/p3_lutinv ),
    .c(\ADD02/ADD03/ADD02/n1 ),
    .d(\ADD02/ADD03/ADD02/p2_lutinv ),
    .o(_al_u463_o));
  AL_MAP_LUT5 #(
    .EQN("(C@(D*A*~(E*~B)))"),
    .INIT(32'h78f05af0))
    _al_u464 (
    .a(_al_u461_o),
    .b(_al_u459_o),
    .c(_al_u462_o),
    .d(_al_u463_o),
    .e(_al_u420_o),
    .o(M_result2[8]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u465 (
    .a(_al_u259_o),
    .b(_al_u433_o),
    .o(_al_u465_o));
  AL_MAP_LUT5 #(
    .EQN("(C@(D*~B*~(E*~A)))"),
    .INIT(32'hd2f0c3f0))
    _al_u466 (
    .a(_al_u459_o),
    .b(_al_u465_o),
    .c(_al_u439_o),
    .d(_al_u400_o),
    .e(_al_u420_o),
    .o(M_result2[7]));
  AL_MAP_LUT5 #(
    .EQN("~(C@(D*~B*~(E*~A)))"),
    .INIT(32'h2d0f3c0f))
    _al_u467 (
    .a(_al_u459_o),
    .b(_al_u433_o),
    .c(_al_u442_o),
    .d(_al_u400_o),
    .e(_al_u420_o),
    .o(M_result2[6]));
  AL_MAP_LUT4 #(
    .EQN("~(D@(B*~(~C*A)))"),
    .INIT(16'hc43b))
    _al_u468 (
    .a(_al_u284_o),
    .b(_al_u311_o),
    .c(_al_u312_o),
    .d(_al_u438_o),
    .o(_al_u468_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u469 (
    .a(_al_u431_o),
    .b(_al_u468_o),
    .o(_al_u469_o));
  AL_MAP_LUT4 #(
    .EQN("~(C@(~D*~(~B*~A)))"),
    .INIT(16'h0fe1))
    _al_u470 (
    .a(_al_u435_o),
    .b(_al_u438_o),
    .c(\ADD02/ADD01/ADD02/p1_lutinv ),
    .d(\ADD02/ADD01/ADD02/g0 ),
    .o(_al_u470_o));
  AL_MAP_LUT5 #(
    .EQN("(C@(D*~B*~(E*~A)))"),
    .INIT(32'hd2f0c3f0))
    _al_u471 (
    .a(_al_u459_o),
    .b(_al_u469_o),
    .c(_al_u470_o),
    .d(_al_u400_o),
    .e(_al_u420_o),
    .o(M_result2[5]));
  AL_MAP_LUT5 #(
    .EQN("~(E@(~D*B*~(C*~A)))"),
    .INIT(32'h008cff73))
    _al_u472 (
    .a(_al_u459_o),
    .b(_al_u400_o),
    .c(_al_u420_o),
    .d(_al_u431_o),
    .e(_al_u468_o),
    .o(M_result2[4]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u473 (
    .a(_al_u284_o),
    .b(\ADD02/ADD01/ADD01/p2_lutinv ),
    .o(_al_u473_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*~A))"),
    .INIT(8'he0))
    _al_u474 (
    .a(_al_u473_o),
    .b(_al_u428_o),
    .c(_al_u212_o),
    .o(_al_u474_o));
  AL_MAP_LUT4 #(
    .EQN("(C@~(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B))"),
    .INIT(16'h87b4))
    _al_u475 (
    .a(_al_u284_o),
    .b(\ADD02/ADD01/ADD01/p2_lutinv ),
    .c(\ADD02/ADD01/ADD01/p3_lutinv ),
    .d(_al_u289_o),
    .o(_al_u475_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@(C*B*~(D*~A)))"),
    .INIT(32'h80c07f3f))
    _al_u476 (
    .a(_al_u459_o),
    .b(_al_u474_o),
    .c(_al_u463_o),
    .d(_al_u420_o),
    .e(_al_u475_o),
    .o(M_result2[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u477 (
    .a(_al_u428_o),
    .b(_al_u212_o),
    .o(_al_u477_o));
  AL_MAP_LUT5 #(
    .EQN("(D@(E*B*~(C*~A)))"),
    .INIT(32'h738cff00))
    _al_u478 (
    .a(_al_u459_o),
    .b(_al_u463_o),
    .c(_al_u420_o),
    .d(_al_u473_o),
    .e(_al_u477_o),
    .o(M_result2[2]));
  AL_MAP_LUT5 #(
    .EQN("~(C@B@(~A*~(E@D)))"),
    .INIT(32'h96c3c396))
    _al_u479 (
    .a(_al_u427_o),
    .b(_al_u275_o),
    .c(_al_u283_o),
    .d(_al_u266_o),
    .e(_al_u212_o),
    .o(\C03/outtemp [1]));
  AL_MAP_LUT5 #(
    .EQN("~(D@(E*B*~(C*~A)))"),
    .INIT(32'h8c7300ff))
    _al_u480 (
    .a(_al_u459_o),
    .b(_al_u400_o),
    .c(_al_u420_o),
    .d(\C03/outtemp [1]),
    .e(M_result[0]),
    .o(M_result2[1]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u481 (
    .a(_al_u439_o),
    .b(_al_u259_o),
    .c(\ADD02/ADD02/ADD01/p0_lutinv ),
    .o(_al_u481_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u482 (
    .a(_al_u481_o),
    .b(_al_u450_o),
    .c(_al_u433_o),
    .d(\ADD02/ADD02/ADD01/p2_lutinv ),
    .o(_al_u482_o));
  AL_MAP_LUT4 #(
    .EQN("(B@(~C*~(D*~A)))"),
    .INIT(16'hc6c3))
    _al_u483 (
    .a(_al_u448_o),
    .b(\ADD02/ADD02/ADD02/p1_lutinv ),
    .c(\ADD02/ADD02/ADD02/g0 ),
    .d(\ADD02/ADD02/ADD02/p0_lutinv ),
    .o(_al_u483_o));
  AL_MAP_LUT4 #(
    .EQN("~(D@(B*~(~C*A)))"),
    .INIT(16'hc43b))
    _al_u484 (
    .a(_al_u482_o),
    .b(_al_u426_o),
    .c(_al_u449_o),
    .d(_al_u483_o),
    .o(M_result2[13]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u485 (
    .a(\ADD02/ADD02/ADD02/p2_lutinv ),
    .b(\ADD02/ADD02/ADD02/p1_lutinv ),
    .c(\ADD02/ADD02/ADD02/p0_lutinv ),
    .o(_al_u485_o));
  AL_MAP_LUT3 #(
    .EQN("(A*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'he8))
    _al_u486 (
    .a(_al_u327_o),
    .b(_al_u330_o),
    .c(_al_u332_o),
    .o(_al_u486_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B*~A)))"),
    .INIT(16'h4fb0))
    _al_u487 (
    .a(_al_u448_o),
    .b(_al_u485_o),
    .c(_al_u486_o),
    .d(\ADD02/ADD02/ADD02/p3_lutinv ),
    .o(_al_u487_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u488 (
    .a(\ADD02/ADD02/ADD02/p1_lutinv ),
    .b(\ADD02/ADD02/ADD02/p0_lutinv ),
    .o(\ADD02/ADD02/ADD02/n3 ));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B*~A)))"),
    .INIT(16'h4fb0))
    _al_u489 (
    .a(_al_u448_o),
    .b(\ADD02/ADD02/ADD02/n3 ),
    .c(_al_u327_o),
    .d(\ADD02/ADD02/ADD02/p2_lutinv ),
    .o(_al_u489_o));
  AL_MAP_LUT5 #(
    .EQN("~(C@(B*~(E*D*A)))"),
    .INIT(32'h4bc3c3c3))
    _al_u490 (
    .a(_al_u482_o),
    .b(_al_u426_o),
    .c(_al_u487_o),
    .d(_al_u489_o),
    .e(\ADD02/ADD02/ADD02/n3 ),
    .o(M_result2[15]));
  AL_MAP_LUT5 #(
    .EQN("~(E@(B*~(D*~C*A)))"),
    .INIT(32'hc4cc3b33))
    _al_u491 (
    .a(_al_u482_o),
    .b(_al_u426_o),
    .c(_al_u449_o),
    .d(_al_u483_o),
    .e(_al_u489_o),
    .o(M_result2[14]));
  AL_MAP_LUT5 #(
    .EQN("(D*~(E)*~((~(C*~A)*B))+D*E*~((~(C*~A)*B))+~(D)*E*(~(C*~A)*B)+D*E*(~(C*~A)*B))"),
    .INIT(32'hff8c7300))
    _al_u492 (
    .a(_al_u459_o),
    .b(_al_u463_o),
    .c(_al_u420_o),
    .d(n1[31]),
    .e(n2[31]),
    .o(result[31]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u493 (
    .a(_al_u450_o),
    .b(\ADD02/ADD02/ADD01/p2_lutinv ),
    .o(\ADD02/ADD02/ADD01/n17 ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u494 (
    .a(\ADD02/ADD02/ADD01/n17 ),
    .b(\ADD02/ADD02/ADD02/n3 ),
    .c(_al_u433_o),
    .d(_al_u481_o),
    .o(_al_u494_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u495 (
    .a(_al_u487_o),
    .b(\ADD02/ADD02/ADD02/p2_lutinv ),
    .o(_al_u495_o));
  AL_MAP_LUT4 #(
    .EQN("~(D@(B*~(C*~A)))"),
    .INIT(16'h8c73))
    _al_u496 (
    .a(_al_u448_o),
    .b(_al_u341_o),
    .c(_al_u344_o),
    .d(\ADD02/ADD03/ADD01/p0_lutinv ),
    .o(_al_u496_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*~(B*A)))"),
    .INIT(16'h8f70))
    _al_u497 (
    .a(_al_u494_o),
    .b(_al_u495_o),
    .c(_al_u426_o),
    .d(_al_u496_o),
    .o(M_result2[16]));
  AL_MAP_LUT5 #(
    .EQN("(B@(A*C*~((E@D))+A*~(C)*(E@D)+~(A)*C*(E@D)+A*C*(E@D)))"),
    .INIT(32'h6c36366c))
    _al_u498 (
    .a(_al_u380_o),
    .b(\ADD02/ADD03/ADD01/p1_lutinv ),
    .c(_al_u402_o),
    .d(_al_u403_o),
    .e(_al_u212_o),
    .o(_al_u498_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@(C*~(~E*B*A)))"),
    .INIT(32'hf00f708f))
    _al_u499 (
    .a(_al_u494_o),
    .b(_al_u495_o),
    .c(_al_u426_o),
    .d(_al_u498_o),
    .e(_al_u496_o),
    .o(M_result2[17]));
  AL_MAP_LUT4 #(
    .EQN("~(A@(B*(D@C)))"),
    .INIT(16'h5995))
    _al_u500 (
    .a(\ADD02/ADD03/ADD01/p1_lutinv ),
    .b(_al_u402_o),
    .c(_al_u403_o),
    .d(_al_u212_o),
    .o(_al_u500_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u501 (
    .a(_al_u500_o),
    .b(\ADD02/ADD03/ADD01/p2_lutinv ),
    .c(\ADD02/ADD03/ADD01/p0_lutinv ),
    .o(_al_u501_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u502 (
    .a(\ADD02/ADD03/ADD01/p0_lutinv ),
    .b(\ADD02/ADD03/ADD01/p1_lutinv ),
    .o(\ADD02/ADD03/ADD01/n3 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u503 (
    .a(\ADD02/ADD03/ADD01/n3 ),
    .b(\ADD02/ADD03/ADD01/p2_lutinv ),
    .o(_al_u503_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(~C*~(B*~A)))"),
    .INIT(16'hf40b))
    _al_u504 (
    .a(_al_u380_o),
    .b(_al_u503_o),
    .c(_al_u413_o),
    .d(\ADD02/ADD03/ADD01/p3_lutinv ),
    .o(_al_u504_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@(D*~(C*B*A)))"),
    .INIT(32'h7f0080ff))
    _al_u505 (
    .a(_al_u494_o),
    .b(_al_u495_o),
    .c(_al_u501_o),
    .d(_al_u426_o),
    .e(_al_u504_o),
    .o(M_result2[19]));
  AL_MAP_LUT5 #(
    .EQN("(D@(~E*~C*~(B*~A)))"),
    .INIT(32'hff00f40b))
    _al_u506 (
    .a(_al_u380_o),
    .b(\ADD02/ADD03/ADD01/n3 ),
    .c(_al_u407_o),
    .d(\ADD02/ADD03/ADD01/p2_lutinv ),
    .e(\ADD02/ADD03/ADD01/g1 ),
    .o(_al_u506_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u507 (
    .a(_al_u500_o),
    .b(\ADD02/ADD03/ADD01/p0_lutinv ),
    .o(_al_u507_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@(C*~(E*B*A)))"),
    .INIT(32'h708ff00f))
    _al_u508 (
    .a(_al_u494_o),
    .b(_al_u495_o),
    .c(_al_u426_o),
    .d(_al_u506_o),
    .e(_al_u507_o),
    .o(M_result2[18]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u509 (
    .a(_al_u507_o),
    .b(\ADD02/ADD03/ADD01/p2_lutinv ),
    .c(\ADD02/ADD03/ADD01/p3_lutinv ),
    .o(_al_u509_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@(~B*~(D*C*~A)))"),
    .INIT(32'h2333dccc))
    _al_u510 (
    .a(_al_u380_o),
    .b(_al_u417_o),
    .c(_al_u503_o),
    .d(\ADD02/ADD03/ADD01/p3_lutinv ),
    .e(\ADD02/ADD03/ADD02/p0_lutinv ),
    .o(_al_u510_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*~(C*B*A)))"),
    .INIT(32'h80ff7f00))
    _al_u511 (
    .a(_al_u509_o),
    .b(_al_u494_o),
    .c(_al_u495_o),
    .d(_al_u426_o),
    .e(_al_u510_o),
    .o(M_result2[20]));
  AL_MAP_LUT4 #(
    .EQN("(D@(~B*~(C*~A)))"),
    .INIT(16'hdc23))
    _al_u512 (
    .a(_al_u459_o),
    .b(\ADD02/ADD03/ADD02/g0 ),
    .c(\ADD02/ADD03/ADD02/p0_lutinv ),
    .d(\ADD02/ADD03/ADD02/p1_lutinv ),
    .o(_al_u512_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u513 (
    .a(\ADD02/ADD02/ADD01/n17 ),
    .b(_al_u481_o),
    .c(_al_u507_o),
    .d(\ADD02/ADD02/ADD02/n3 ),
    .e(_al_u433_o),
    .o(_al_u513_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u514 (
    .a(\ADD02/ADD03/ADD01/p2_lutinv ),
    .b(\ADD02/ADD03/ADD01/p3_lutinv ),
    .o(\ADD02/ADD03/ADD01/n14 ));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u515 (
    .a(_al_u513_o),
    .b(\ADD02/ADD03/ADD01/n14 ),
    .c(_al_u495_o),
    .d(_al_u426_o),
    .o(_al_u515_o));
  AL_MAP_LUT4 #(
    .EQN("~(A@(B*~(~D*~C)))"),
    .INIT(16'h9995))
    _al_u516 (
    .a(_al_u512_o),
    .b(_al_u426_o),
    .c(_al_u510_o),
    .d(_al_u515_o),
    .o(M_result2[21]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u517 (
    .a(\ADD02/ADD03/ADD02/n1 ),
    .b(\ADD02/ADD03/ADD02/g1 ),
    .o(_al_u517_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(B*~(C*~A)))"),
    .INIT(16'h738c))
    _al_u518 (
    .a(_al_u459_o),
    .b(_al_u517_o),
    .c(\ADD02/ADD03/ADD02/n3 ),
    .d(\ADD02/ADD03/ADD02/p2_lutinv ),
    .o(_al_u518_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u519 (
    .a(_al_u509_o),
    .b(_al_u494_o),
    .c(_al_u495_o),
    .d(_al_u518_o),
    .e(\ADD02/ADD03/ADD02/n3 ),
    .o(_al_u519_o));
  AL_MAP_LUT4 #(
    .EQN("~(A@(~B*~(D*C)))"),
    .INIT(16'h5666))
    _al_u520 (
    .a(\ADD02/ADD03/ADD02/p3_lutinv ),
    .b(\ADD02/ADD03/ADD02/g2 ),
    .c(\ADD02/ADD03/ADD02/p2_lutinv ),
    .d(_al_u518_o),
    .o(_al_u520_o));
  AL_MAP_LUT3 #(
    .EQN("(B@(C*~A))"),
    .INIT(8'h9c))
    _al_u521 (
    .a(_al_u519_o),
    .b(_al_u520_o),
    .c(_al_u426_o),
    .o(M_result2[23]));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u522 (
    .a(\ADD02/ADD03/ADD02/n3 ),
    .b(_al_u443_o),
    .c(_al_u447_o),
    .d(_al_u450_o),
    .e(\ADD02/ADD02/ADD02/n3 ),
    .o(_al_u522_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@(E*~(C*B*A)))"),
    .INIT(32'h7f8000ff))
    _al_u523 (
    .a(_al_u522_o),
    .b(_al_u509_o),
    .c(_al_u495_o),
    .d(_al_u518_o),
    .e(_al_u426_o),
    .o(M_result2[22]));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u524 (
    .a(_al_u459_o),
    .b(_al_u463_o),
    .c(_al_u420_o),
    .o(_al_u524_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u525 (
    .a(_al_u524_o),
    .b(_al_u212_o),
    .o(_al_u525_o));
  AL_MAP_LUT4 #(
    .EQN("((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'haca0))
    _al_u526 (
    .a(\NM/n4 [0]),
    .b(M_result2[23]),
    .c(_al_u525_o),
    .d(M_result[0]),
    .o(result[0]));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u527 (
    .a(_al_u522_o),
    .b(_al_u509_o),
    .c(_al_u495_o),
    .o(_al_u527_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb7fc))
    _al_u528 (
    .a(_al_u527_o),
    .b(_al_u520_o),
    .c(_al_u518_o),
    .d(_al_u426_o),
    .o(_al_u528_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u529 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[1]),
    .d(M_result[0]),
    .o(_al_u529_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'ha3))
    _al_u530 (
    .a(\NM/n4 [1]),
    .b(_al_u529_o),
    .c(_al_u525_o),
    .o(result[1]));
  AL_MAP_LUT5 #(
    .EQN("(~(B)*~(D)*~((E*C*~A))+B*~(D)*~((E*C*~A))+B*D*~((E*C*~A))+~(B)*~(D)*(E*C*~A)+~(B)*D*(E*C*~A)+B*D*(E*C*~A))"),
    .INIT(32'hdcbfccff))
    _al_u531 (
    .a(_al_u527_o),
    .b(_al_u520_o),
    .c(_al_u524_o),
    .d(_al_u518_o),
    .e(_al_u212_o),
    .o(_al_u531_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u532 (
    .a(_al_u531_o),
    .b(M_result2[21]),
    .o(_al_u532_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u533 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[2]),
    .d(M_result2[1]),
    .o(_al_u533_o));
  AL_MAP_LUT5 #(
    .EQN("(~(C*~(E*B))*~(A)*~(D)+~(C*~(E*B))*A*~(D)+~(~(C*~(E*B)))*A*D+~(C*~(E*B))*A*D)"),
    .INIT(32'haacfaa0f))
    _al_u534 (
    .a(\NM/n4 [2]),
    .b(_al_u532_o),
    .c(_al_u533_o),
    .d(_al_u525_o),
    .e(M_result[0]),
    .o(result[2]));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u535 (
    .a(_al_u531_o),
    .b(M_result2[21]),
    .c(M_result2[20]),
    .o(_al_u535_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u536 (
    .a(_al_u532_o),
    .b(_al_u535_o),
    .c(M_result2[1]),
    .d(M_result[0]),
    .o(_al_u536_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u537 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[3]),
    .d(M_result2[2]),
    .o(_al_u537_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(A)*~(D)+~(C*B)*A*~(D)+~(~(C*B))*A*D+~(C*B)*A*D)"),
    .INIT(16'haa3f))
    _al_u538 (
    .a(\NM/n4 [3]),
    .b(_al_u536_o),
    .c(_al_u537_o),
    .d(_al_u525_o),
    .o(result[3]));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*~(B)*~(C)+A*B*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'hdb))
    _al_u539 (
    .a(_al_u515_o),
    .b(_al_u512_o),
    .c(_al_u510_o),
    .o(_al_u539_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u540 (
    .a(_al_u531_o),
    .b(_al_u539_o),
    .o(_al_u540_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u541 (
    .a(_al_u540_o),
    .b(M_result2[19]),
    .o(_al_u541_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*B)*~(E*~A))"),
    .INIT(32'h020a030f))
    _al_u542 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(_al_u525_o),
    .d(M_result2[4]),
    .e(M_result2[3]),
    .o(_al_u542_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D*B)*~(E*A))"),
    .INIT(32'h105030f0))
    _al_u543 (
    .a(_al_u541_o),
    .b(_al_u532_o),
    .c(_al_u542_o),
    .d(M_result2[2]),
    .e(M_result[0]),
    .o(_al_u543_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~(E*C)*B)*~(D*~A))"),
    .INIT(32'ha2f32233))
    _al_u544 (
    .a(\NM/n4 [4]),
    .b(_al_u543_o),
    .c(_al_u535_o),
    .d(_al_u525_o),
    .e(M_result2[1]),
    .o(result[4]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u545 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[5]),
    .d(M_result2[4]),
    .o(_al_u545_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u546 (
    .a(_al_u532_o),
    .b(_al_u545_o),
    .c(M_result2[3]),
    .o(_al_u546_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u547 (
    .a(_al_u546_o),
    .b(_al_u541_o),
    .c(_al_u535_o),
    .d(M_result2[2]),
    .e(M_result2[1]),
    .o(_al_u547_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u548 (
    .a(_al_u531_o),
    .b(M_result2[21]),
    .o(_al_u548_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*~(B)*~(C)+A*B*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'hdb))
    _al_u549 (
    .a(_al_u426_o),
    .b(_al_u504_o),
    .c(_al_u510_o),
    .o(_al_u549_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u550 (
    .a(_al_u548_o),
    .b(_al_u549_o),
    .c(M_result2[18]),
    .o(_al_u550_o));
  AL_MAP_LUT5 #(
    .EQN("(~(B*~(E*C))*~(A)*~(D)+~(B*~(E*C))*A*~(D)+~(~(B*~(E*C)))*A*D+~(B*~(E*C))*A*D)"),
    .INIT(32'haaf3aa33))
    _al_u551 (
    .a(\NM/n4 [5]),
    .b(_al_u547_o),
    .c(_al_u550_o),
    .d(_al_u525_o),
    .e(M_result[0]),
    .o(result[5]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u552 (
    .a(_al_u532_o),
    .b(_al_u535_o),
    .c(M_result2[4]),
    .d(M_result2[3]),
    .o(_al_u552_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'heff7))
    _al_u553 (
    .a(_al_u512_o),
    .b(_al_u504_o),
    .c(_al_u510_o),
    .d(_al_u426_o),
    .o(_al_u553_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u554 (
    .a(_al_u531_o),
    .b(_al_u553_o),
    .c(M_result2[18]),
    .o(_al_u554_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u555 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[6]),
    .d(M_result2[5]),
    .o(_al_u555_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u556 (
    .a(_al_u552_o),
    .b(_al_u554_o),
    .c(_al_u555_o),
    .d(M_result2[1]),
    .o(_al_u556_o));
  AL_MAP_LUT5 #(
    .EQN("(~((C*~(B*A)))*~(D)*~(E)+~((C*~(B*A)))*D*~(E)+(C*~(B*A))*D*~(E)+~((C*~(B*A)))*~(D)*E+(C*~(B*A))*~(D)*E+(C*~(B*A))*D*E)"),
    .INIT(32'h70ffff8f))
    _al_u557 (
    .a(_al_u513_o),
    .b(_al_u495_o),
    .c(_al_u426_o),
    .d(_al_u506_o),
    .e(_al_u504_o),
    .o(_al_u557_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(~(B)*C*~(D)+B*~(C)*D))"),
    .INIT(16'h0410))
    _al_u558 (
    .a(_al_u557_o),
    .b(_al_u515_o),
    .c(_al_u512_o),
    .d(_al_u510_o),
    .o(_al_u558_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u559 (
    .a(_al_u531_o),
    .b(_al_u558_o),
    .o(_al_u559_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u560 (
    .a(_al_u559_o),
    .b(M_result2[17]),
    .o(_al_u560_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u561 (
    .a(_al_u541_o),
    .b(_al_u560_o),
    .c(M_result2[2]),
    .d(M_result[0]),
    .o(_al_u561_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(A)*~(D)+~(C*B)*A*~(D)+~(~(C*B))*A*D+~(C*B)*A*D)"),
    .INIT(16'haa3f))
    _al_u562 (
    .a(\NM/n4 [6]),
    .b(_al_u556_o),
    .c(_al_u561_o),
    .d(_al_u525_o),
    .o(result[6]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u563 (
    .a(_al_u541_o),
    .b(_al_u560_o),
    .c(M_result2[4]),
    .d(M_result2[2]),
    .o(_al_u563_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*(D@C))"),
    .INIT(16'h0110))
    _al_u564 (
    .a(M_result2[19]),
    .b(M_result2[17]),
    .c(_al_u506_o),
    .d(_al_u426_o),
    .o(_al_u564_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u565 (
    .a(_al_u540_o),
    .b(_al_u564_o),
    .c(M_result2[16]),
    .o(_al_u565_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u566 (
    .a(_al_u531_o),
    .b(_al_u553_o),
    .o(_al_u566_o));
  AL_MAP_LUT5 #(
    .EQN("(~((C*~(B*A)))*~(D)*~(E)+(C*~(B*A))*~(D)*~(E)+(C*~(B*A))*D*~(E)+~((C*~(B*A)))*~(D)*E+~((C*~(B*A)))*D*E+(C*~(B*A))*D*E)"),
    .INIT(32'hff8f70ff))
    _al_u567 (
    .a(_al_u494_o),
    .b(_al_u495_o),
    .c(_al_u426_o),
    .d(_al_u498_o),
    .e(_al_u496_o),
    .o(_al_u567_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u568 (
    .a(M_result2[18]),
    .b(_al_u567_o),
    .c(M_result2[15]),
    .o(_al_u568_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u569 (
    .a(_al_u566_o),
    .b(_al_u568_o),
    .o(_al_u569_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u570 (
    .a(_al_u563_o),
    .b(_al_u565_o),
    .c(_al_u569_o),
    .d(M_result2[1]),
    .e(M_result[0]),
    .o(_al_u570_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u571 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[8]),
    .d(M_result2[7]),
    .o(_al_u571_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(D*A))"),
    .INIT(16'h040c))
    _al_u572 (
    .a(_al_u554_o),
    .b(_al_u571_o),
    .c(_al_u525_o),
    .d(M_result2[3]),
    .o(_al_u572_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u573 (
    .a(_al_u572_o),
    .b(_al_u532_o),
    .c(_al_u535_o),
    .d(M_result2[6]),
    .e(M_result2[5]),
    .o(_al_u573_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u574 (
    .a(\NM/n4 [8]),
    .b(_al_u570_o),
    .c(_al_u573_o),
    .d(_al_u525_o),
    .o(result[8]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u575 (
    .a(_al_u532_o),
    .b(_al_u554_o),
    .c(M_result2[5]),
    .d(M_result2[2]),
    .o(_al_u575_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u576 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[7]),
    .d(M_result2[6]),
    .o(_al_u576_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u577 (
    .a(_al_u575_o),
    .b(_al_u535_o),
    .c(_al_u576_o),
    .d(M_result2[4]),
    .o(_al_u577_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u578 (
    .a(_al_u541_o),
    .b(_al_u560_o),
    .c(M_result2[3]),
    .d(M_result2[1]),
    .o(_al_u578_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u579 (
    .a(_al_u577_o),
    .b(_al_u578_o),
    .c(_al_u565_o),
    .d(M_result[0]),
    .o(_al_u579_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'ha3))
    _al_u580 (
    .a(\NM/n4 [7]),
    .b(_al_u579_o),
    .c(_al_u525_o),
    .o(result[7]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u581 (
    .a(_al_u541_o),
    .b(M_result2[5]),
    .o(_al_u581_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u582 (
    .a(_al_u566_o),
    .b(M_result2[18]),
    .o(_al_u582_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*C)*~(D*B))"),
    .INIT(32'h01051155))
    _al_u583 (
    .a(_al_u581_o),
    .b(_al_u582_o),
    .c(_al_u565_o),
    .d(M_result2[4]),
    .e(M_result2[2]),
    .o(_al_u583_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hfdbf))
    _al_u584 (
    .a(_al_u426_o),
    .b(_al_u498_o),
    .c(_al_u506_o),
    .d(_al_u496_o),
    .o(_al_u584_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u585 (
    .a(_al_u584_o),
    .b(M_result2[15]),
    .c(M_result2[14]),
    .o(_al_u585_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u586 (
    .a(_al_u566_o),
    .b(_al_u585_o),
    .o(_al_u586_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u587 (
    .a(_al_u569_o),
    .b(_al_u586_o),
    .c(M_result2[1]),
    .d(M_result[0]),
    .o(_al_u587_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u588 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[9]),
    .d(M_result2[8]),
    .o(_al_u588_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E*B)*~(D*A))"),
    .INIT(32'h103050f0))
    _al_u589 (
    .a(_al_u532_o),
    .b(_al_u535_o),
    .c(_al_u588_o),
    .d(M_result2[7]),
    .e(M_result2[6]),
    .o(_al_u589_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u590 (
    .a(_al_u583_o),
    .b(_al_u587_o),
    .c(_al_u589_o),
    .d(_al_u525_o),
    .o(_al_u590_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~(E*C)*B)*~(D*~A))"),
    .INIT(32'ha2f32233))
    _al_u591 (
    .a(\NM/n4 [9]),
    .b(_al_u590_o),
    .c(_al_u560_o),
    .d(_al_u525_o),
    .e(M_result2[3]),
    .o(result[9]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u592 (
    .a(_al_u567_o),
    .b(M_result2[15]),
    .o(_al_u592_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hcfffff7b))
    _al_u593 (
    .a(_al_u482_o),
    .b(_al_u426_o),
    .c(_al_u449_o),
    .d(_al_u483_o),
    .e(_al_u489_o),
    .o(_al_u593_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u594 (
    .a(_al_u559_o),
    .b(_al_u592_o),
    .c(_al_u593_o),
    .o(_al_u594_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u595 (
    .a(_al_u594_o),
    .b(M_result[0]),
    .o(_al_u595_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*C)*~(D*B))"),
    .INIT(32'h01051155))
    _al_u596 (
    .a(_al_u595_o),
    .b(_al_u569_o),
    .c(_al_u586_o),
    .d(M_result2[3]),
    .e(M_result2[2]),
    .o(_al_u596_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u597 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[11]),
    .d(M_result2[10]),
    .o(_al_u597_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E*B)*~(D*A))"),
    .INIT(32'h103050f0))
    _al_u598 (
    .a(_al_u532_o),
    .b(_al_u535_o),
    .c(_al_u597_o),
    .d(M_result2[9]),
    .e(M_result2[8]),
    .o(_al_u598_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u599 (
    .a(_al_u426_o),
    .b(_al_u489_o),
    .o(_al_u599_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u600 (
    .a(_al_u559_o),
    .b(_al_u592_o),
    .c(M_result2[13]),
    .d(_al_u599_o),
    .o(_al_u600_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*B*A*~(E*C))"),
    .INIT(32'h00080088))
    _al_u601 (
    .a(_al_u596_o),
    .b(_al_u598_o),
    .c(_al_u600_o),
    .d(_al_u525_o),
    .e(M_result2[1]),
    .o(_al_u601_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u602 (
    .a(_al_u601_o),
    .b(_al_u541_o),
    .c(_al_u565_o),
    .d(M_result2[7]),
    .e(M_result2[4]),
    .o(_al_u602_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u603 (
    .a(_al_u582_o),
    .b(_al_u560_o),
    .c(M_result2[6]),
    .d(M_result2[5]),
    .o(_al_u603_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u604 (
    .a(\NM/n4 [11]),
    .b(_al_u602_o),
    .c(_al_u603_o),
    .d(_al_u525_o),
    .o(result[11]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u605 (
    .a(_al_u541_o),
    .b(M_result2[6]),
    .o(_al_u605_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*C)*~(D*B))"),
    .INIT(32'h01051155))
    _al_u606 (
    .a(_al_u605_o),
    .b(_al_u582_o),
    .c(_al_u560_o),
    .d(M_result2[5]),
    .e(M_result2[4]),
    .o(_al_u606_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u607 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[10]),
    .d(M_result2[9]),
    .o(_al_u607_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E*B)*~(D*A))"),
    .INIT(32'h103050f0))
    _al_u608 (
    .a(_al_u532_o),
    .b(_al_u535_o),
    .c(_al_u607_o),
    .d(M_result2[8]),
    .e(M_result2[7]),
    .o(_al_u608_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u609 (
    .a(_al_u608_o),
    .b(_al_u586_o),
    .c(_al_u525_o),
    .d(M_result2[1]),
    .o(_al_u609_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u610 (
    .a(_al_u600_o),
    .b(M_result[0]),
    .o(_al_u610_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*A*~(E*D))"),
    .INIT(32'h00080808))
    _al_u611 (
    .a(_al_u606_o),
    .b(_al_u609_o),
    .c(_al_u610_o),
    .d(_al_u569_o),
    .e(M_result2[2]),
    .o(_al_u611_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~(E*C)*B)*~(D*~A))"),
    .INIT(32'ha2f32233))
    _al_u612 (
    .a(\NM/n4 [10]),
    .b(_al_u611_o),
    .c(_al_u565_o),
    .d(_al_u525_o),
    .e(M_result2[3]),
    .o(result[10]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u613 (
    .a(_al_u541_o),
    .b(M_result2[8]),
    .o(_al_u613_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*C)*~(D*B))"),
    .INIT(32'h01051155))
    _al_u614 (
    .a(_al_u613_o),
    .b(_al_u550_o),
    .c(_al_u565_o),
    .d(M_result2[7]),
    .e(M_result2[5]),
    .o(_al_u614_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u615 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[12]),
    .d(M_result2[11]),
    .o(_al_u615_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E*B)*~(D*A))"),
    .INIT(32'h103050f0))
    _al_u616 (
    .a(_al_u532_o),
    .b(_al_u535_o),
    .c(_al_u615_o),
    .d(M_result2[10]),
    .e(M_result2[9]),
    .o(_al_u616_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u617 (
    .a(_al_u616_o),
    .b(_al_u560_o),
    .c(M_result2[6]),
    .o(_al_u617_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u618 (
    .a(_al_u614_o),
    .b(_al_u617_o),
    .c(_al_u586_o),
    .d(M_result2[3]),
    .o(_al_u618_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u619 (
    .a(_al_u600_o),
    .b(_al_u594_o),
    .c(M_result2[2]),
    .d(M_result2[1]),
    .o(_al_u619_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u620 (
    .a(_al_u564_o),
    .b(_al_u539_o),
    .o(_al_u620_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u621 (
    .a(_al_u620_o),
    .b(_al_u531_o),
    .o(_al_u621_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'heff7))
    _al_u622 (
    .a(_al_u426_o),
    .b(_al_u449_o),
    .c(_al_u483_o),
    .d(_al_u489_o),
    .o(_al_u622_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u623 (
    .a(M_result2[16]),
    .b(M_result2[15]),
    .c(_al_u622_o),
    .d(M_result2[11]),
    .o(_al_u623_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u624 (
    .a(_al_u621_o),
    .b(_al_u623_o),
    .o(_al_u624_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u625 (
    .a(_al_u619_o),
    .b(_al_u624_o),
    .c(_al_u569_o),
    .d(M_result2[4]),
    .e(M_result[0]),
    .o(_al_u625_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(A)*~(D)+~(C*B)*A*~(D)+~(~(C*B))*A*D+~(C*B)*A*D)"),
    .INIT(16'haa3f))
    _al_u626 (
    .a(\NM/n4 [12]),
    .b(_al_u618_o),
    .c(_al_u625_o),
    .d(_al_u525_o),
    .o(result[12]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*B)*~(C*~A))"),
    .INIT(32'h000023af))
    _al_u627 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[13]),
    .d(M_result2[14]),
    .e(_al_u525_o),
    .o(_al_u627_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D*B)*~(E*A))"),
    .INIT(32'h105030f0))
    _al_u628 (
    .a(_al_u624_o),
    .b(_al_u535_o),
    .c(_al_u627_o),
    .d(M_result2[11]),
    .e(M_result2[2]),
    .o(_al_u628_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u629 (
    .a(_al_u628_o),
    .b(_al_u541_o),
    .c(_al_u569_o),
    .d(M_result2[10]),
    .e(M_result2[6]),
    .o(_al_u629_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u630 (
    .a(_al_u565_o),
    .b(M_result2[7]),
    .o(_al_u630_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u631 (
    .a(M_result2[16]),
    .b(M_result2[15]),
    .o(_al_u631_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C)"),
    .INIT(8'hbd))
    _al_u632 (
    .a(_al_u426_o),
    .b(_al_u483_o),
    .c(_al_u489_o),
    .o(_al_u632_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C+~(A)*B*C)"),
    .INIT(8'h7e))
    _al_u633 (
    .a(_al_u426_o),
    .b(_al_u449_o),
    .c(_al_u456_o),
    .o(_al_u633_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u634 (
    .a(_al_u631_o),
    .b(_al_u632_o),
    .c(_al_u633_o),
    .d(M_result2[10]),
    .o(_al_u634_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u635 (
    .a(_al_u621_o),
    .b(_al_u634_o),
    .o(_al_u635_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u636 (
    .a(_al_u630_o),
    .b(_al_u635_o),
    .c(M_result2[1]),
    .o(_al_u636_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u637 (
    .a(_al_u629_o),
    .b(_al_u636_o),
    .c(_al_u560_o),
    .d(M_result2[8]),
    .o(_al_u637_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*(D@C))"),
    .INIT(16'h0110))
    _al_u638 (
    .a(_al_u549_o),
    .b(_al_u584_o),
    .c(_al_u512_o),
    .d(_al_u426_o),
    .o(_al_u638_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u639 (
    .a(M_result2[15]),
    .b(_al_u622_o),
    .o(_al_u639_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u64 (
    .a(n1[23]),
    .b(n2[23]),
    .o(_al_u64_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfdf7ffaf))
    _al_u640 (
    .a(_al_u426_o),
    .b(_al_u443_o),
    .c(_al_u447_o),
    .d(_al_u454_o),
    .e(_al_u456_o),
    .o(_al_u640_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u641 (
    .a(_al_u639_o),
    .b(_al_u640_o),
    .o(_al_u641_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u642 (
    .a(_al_u638_o),
    .b(_al_u641_o),
    .c(_al_u531_o),
    .o(_al_u642_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u643 (
    .a(_al_u642_o),
    .b(_al_u554_o),
    .c(M_result2[9]),
    .d(M_result[0]),
    .o(_al_u643_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u644 (
    .a(_al_u643_o),
    .b(_al_u594_o),
    .c(_al_u532_o),
    .d(M_result2[12]),
    .e(M_result2[3]),
    .o(_al_u644_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u645 (
    .a(_al_u638_o),
    .b(_al_u531_o),
    .c(M_result2[15]),
    .d(M_result2[14]),
    .o(_al_u645_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u646 (
    .a(_al_u644_o),
    .b(_al_u600_o),
    .c(_al_u645_o),
    .d(M_result2[5]),
    .e(M_result2[4]),
    .o(_al_u646_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u647 (
    .a(\NM/n4 [14]),
    .b(_al_u637_o),
    .c(_al_u646_o),
    .d(_al_u525_o),
    .o(result[14]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u648 (
    .a(_al_u541_o),
    .b(_al_u550_o),
    .c(M_result2[9]),
    .d(M_result2[8]),
    .o(_al_u648_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u649 (
    .a(_al_u648_o),
    .b(_al_u565_o),
    .c(M_result2[6]),
    .o(_al_u649_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u65 (
    .a(_al_u64_o),
    .b(n2[15]),
    .c(n2[14]),
    .o(n227_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u650 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[13]),
    .d(M_result2[12]),
    .o(_al_u650_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E*B)*~(D*A))"),
    .INIT(32'h103050f0))
    _al_u651 (
    .a(_al_u532_o),
    .b(_al_u535_o),
    .c(_al_u650_o),
    .d(M_result2[11]),
    .e(M_result2[10]),
    .o(_al_u651_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u652 (
    .a(_al_u651_o),
    .b(_al_u560_o),
    .c(_al_u586_o),
    .d(M_result2[7]),
    .e(M_result2[4]),
    .o(_al_u652_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u653 (
    .a(_al_u649_o),
    .b(_al_u652_o),
    .c(_al_u635_o),
    .d(M_result[0]),
    .o(_al_u653_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u654 (
    .a(_al_u600_o),
    .b(_al_u594_o),
    .c(M_result2[3]),
    .d(M_result2[2]),
    .o(_al_u654_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u655 (
    .a(_al_u654_o),
    .b(_al_u624_o),
    .c(_al_u569_o),
    .d(M_result2[5]),
    .e(M_result2[1]),
    .o(_al_u655_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(A)*~(D)+~(C*B)*A*~(D)+~(~(C*B))*A*D+~(C*B)*A*D)"),
    .INIT(16'haa3f))
    _al_u656 (
    .a(\NM/n4 [13]),
    .b(_al_u653_o),
    .c(_al_u655_o),
    .d(_al_u525_o),
    .o(result[13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u657 (
    .a(_al_u532_o),
    .b(M_result2[13]),
    .o(_al_u657_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*B)*~(D*~A))"),
    .INIT(32'h00002a3f))
    _al_u658 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[15]),
    .d(M_result2[14]),
    .e(_al_u525_o),
    .o(_al_u658_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~B*~(D*A))"),
    .INIT(16'h1030))
    _al_u659 (
    .a(_al_u560_o),
    .b(_al_u657_o),
    .c(_al_u658_o),
    .d(M_result2[9]),
    .o(_al_u659_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u66 (
    .a(_al_u64_o),
    .b(n2[13]),
    .c(n2[12]),
    .o(n229_lutinv));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u660 (
    .a(_al_u659_o),
    .b(_al_u624_o),
    .c(_al_u541_o),
    .d(M_result2[11]),
    .e(M_result2[3]),
    .o(_al_u660_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u661 (
    .a(_al_u535_o),
    .b(M_result2[12]),
    .o(_al_u661_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*C)*~(E*B))"),
    .INIT(32'h01110555))
    _al_u662 (
    .a(_al_u661_o),
    .b(_al_u642_o),
    .c(_al_u554_o),
    .d(M_result2[10]),
    .e(M_result2[1]),
    .o(_al_u662_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u663 (
    .a(_al_u660_o),
    .b(_al_u662_o),
    .c(_al_u594_o),
    .d(M_result2[4]),
    .o(_al_u663_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u664 (
    .a(_al_u600_o),
    .b(_al_u645_o),
    .c(M_result2[6]),
    .d(M_result2[5]),
    .o(_al_u664_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u665 (
    .a(M_result2[9]),
    .b(M_result2[8]),
    .o(_al_u665_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*~(B)*~(C)+A*B*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'hdb))
    _al_u666 (
    .a(_al_u426_o),
    .b(_al_u447_o),
    .c(_al_u456_o),
    .o(_al_u666_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*A)"),
    .INIT(16'h0002))
    _al_u667 (
    .a(_al_u665_o),
    .b(M_result2[15]),
    .c(_al_u622_o),
    .d(_al_u666_o),
    .o(_al_u667_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u668 (
    .a(_al_u638_o),
    .b(_al_u531_o),
    .c(_al_u667_o),
    .o(_al_u668_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u669 (
    .a(_al_u664_o),
    .b(_al_u668_o),
    .c(M_result[0]),
    .o(_al_u669_o));
  AL_MAP_LUT4 #(
    .EQN("(C@A@(D*~B))"),
    .INIT(16'h695a))
    _al_u67 (
    .a(n1[24]),
    .b(n1[23]),
    .c(n2[24]),
    .d(n2[23]),
    .o(_al_u67_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u670 (
    .a(_al_u565_o),
    .b(M_result2[8]),
    .o(_al_u670_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*C)*~(E*B))"),
    .INIT(32'h01110555))
    _al_u671 (
    .a(_al_u670_o),
    .b(_al_u635_o),
    .c(_al_u569_o),
    .d(M_result2[7]),
    .e(M_result2[2]),
    .o(_al_u671_o));
  AL_MAP_LUT5 #(
    .EQN("(~(D*C*B)*~(E*~A))"),
    .INIT(32'h2aaa3fff))
    _al_u672 (
    .a(\NM/n4 [15]),
    .b(_al_u663_o),
    .c(_al_u669_o),
    .d(_al_u671_o),
    .e(_al_u525_o),
    .o(result[15]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u673 (
    .a(_al_u621_o),
    .b(_al_u631_o),
    .o(_al_u673_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u674 (
    .a(_al_u633_o),
    .b(M_result2[10]),
    .o(_al_u674_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    _al_u675 (
    .a(_al_u674_o),
    .b(_al_u632_o),
    .c(M_result2[9]),
    .d(M_result2[8]),
    .e(M_result2[7]),
    .o(_al_u675_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u676 (
    .a(_al_u673_o),
    .b(_al_u675_o),
    .o(_al_u676_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*B)*~(D*~A))"),
    .INIT(32'h00002a3f))
    _al_u677 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[16]),
    .d(M_result2[15]),
    .e(_al_u525_o),
    .o(_al_u677_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(D*B)*~(E*A))"),
    .INIT(32'h105030f0))
    _al_u678 (
    .a(_al_u569_o),
    .b(_al_u535_o),
    .c(_al_u677_o),
    .d(M_result2[13]),
    .e(M_result2[8]),
    .o(_al_u678_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(D*C)*~(E*A))"),
    .INIT(32'h04440ccc))
    _al_u679 (
    .a(_al_u676_o),
    .b(_al_u678_o),
    .c(_al_u624_o),
    .d(M_result2[4]),
    .e(M_result[0]),
    .o(_al_u679_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u68 (
    .a(n227_lutinv),
    .b(n229_lutinv),
    .c(_al_u67_o),
    .o(_al_u68_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u680 (
    .a(_al_u541_o),
    .b(_al_u565_o),
    .c(M_result2[12]),
    .d(M_result2[9]),
    .o(_al_u680_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u681 (
    .a(_al_u680_o),
    .b(_al_u635_o),
    .c(_al_u560_o),
    .d(M_result2[10]),
    .e(M_result2[3]),
    .o(_al_u681_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u682 (
    .a(_al_u532_o),
    .b(M_result2[14]),
    .o(_al_u682_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*C)*~(E*B))"),
    .INIT(32'h01110555))
    _al_u683 (
    .a(_al_u682_o),
    .b(_al_u642_o),
    .c(_al_u554_o),
    .d(M_result2[11]),
    .e(M_result2[2]),
    .o(_al_u683_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E*D))"),
    .INIT(32'h00808080))
    _al_u684 (
    .a(_al_u679_o),
    .b(_al_u681_o),
    .c(_al_u683_o),
    .d(_al_u668_o),
    .e(M_result2[1]),
    .o(_al_u684_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u685 (
    .a(_al_u600_o),
    .b(_al_u594_o),
    .c(M_result2[6]),
    .d(M_result2[5]),
    .o(_al_u685_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u686 (
    .a(_al_u685_o),
    .b(_al_u645_o),
    .c(M_result2[7]),
    .o(_al_u686_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u687 (
    .a(\NM/n4 [16]),
    .b(_al_u684_o),
    .c(_al_u686_o),
    .d(_al_u525_o),
    .o(result[16]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u688 (
    .a(_al_u565_o),
    .b(M_result2[10]),
    .o(_al_u688_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u689 (
    .a(_al_u676_o),
    .b(_al_u688_o),
    .c(M_result2[1]),
    .o(_al_u689_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u69 (
    .a(_al_u64_o),
    .b(n2[11]),
    .c(n2[10]),
    .o(n231_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u690 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[17]),
    .d(M_result2[16]),
    .o(_al_u690_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*B*~(D*A))"),
    .INIT(16'h040c))
    _al_u691 (
    .a(_al_u642_o),
    .b(_al_u690_o),
    .c(_al_u525_o),
    .d(M_result2[3]),
    .o(_al_u691_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u692 (
    .a(_al_u689_o),
    .b(_al_u624_o),
    .c(_al_u691_o),
    .d(M_result2[5]),
    .o(_al_u692_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u693 (
    .a(_al_u560_o),
    .b(_al_u569_o),
    .c(M_result2[11]),
    .d(M_result2[9]),
    .o(_al_u693_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u694 (
    .a(_al_u693_o),
    .b(_al_u635_o),
    .c(_al_u541_o),
    .d(M_result2[13]),
    .e(M_result2[4]),
    .o(_al_u694_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u695 (
    .a(_al_u532_o),
    .b(M_result2[15]),
    .o(_al_u695_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*C)*~(D*B))"),
    .INIT(32'h01051155))
    _al_u696 (
    .a(_al_u695_o),
    .b(_al_u535_o),
    .c(_al_u554_o),
    .d(M_result2[14]),
    .e(M_result2[12]),
    .o(_al_u696_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u697 (
    .a(_al_u557_o),
    .b(_al_u567_o),
    .c(M_result2[15]),
    .d(_al_u622_o),
    .o(_al_u697_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u698 (
    .a(_al_u697_o),
    .b(_al_u539_o),
    .o(_al_u698_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u699 (
    .a(_al_u698_o),
    .b(_al_u531_o),
    .o(_al_u699_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u70 (
    .a(_al_u64_o),
    .b(n2[9]),
    .c(n2[8]),
    .o(n233_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(~C*B*A)"),
    .INIT(8'h08))
    _al_u700 (
    .a(_al_u641_o),
    .b(_al_u558_o),
    .c(_al_u567_o),
    .o(_al_u700_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u701 (
    .a(_al_u666_o),
    .b(M_result2[8]),
    .c(M_result2[7]),
    .d(M_result2[6]),
    .o(_al_u701_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u702 (
    .a(_al_u699_o),
    .b(_al_u700_o),
    .c(_al_u701_o),
    .d(M_result[0]),
    .o(_al_u702_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u703 (
    .a(_al_u692_o),
    .b(_al_u694_o),
    .c(_al_u696_o),
    .d(_al_u702_o),
    .o(_al_u703_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u704 (
    .a(_al_u594_o),
    .b(_al_u645_o),
    .c(M_result2[8]),
    .d(M_result2[6]),
    .o(_al_u704_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u705 (
    .a(_al_u704_o),
    .b(_al_u600_o),
    .c(_al_u668_o),
    .d(M_result2[7]),
    .e(M_result2[2]),
    .o(_al_u705_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u706 (
    .a(\NM/n4 [17]),
    .b(_al_u703_o),
    .c(_al_u705_o),
    .d(_al_u525_o),
    .o(result[17]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u707 (
    .a(_al_u624_o),
    .b(M_result2[7]),
    .o(_al_u707_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u708 (
    .a(_al_u707_o),
    .b(_al_u635_o),
    .c(M_result2[6]),
    .o(_al_u708_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u709 (
    .a(_al_u708_o),
    .b(_al_u586_o),
    .c(_al_u535_o),
    .d(M_result2[16]),
    .e(M_result2[10]),
    .o(_al_u709_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u71 (
    .a(n231_lutinv),
    .b(n233_lutinv),
    .c(_al_u67_o),
    .o(_al_u71_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u710 (
    .a(_al_u700_o),
    .b(_al_u531_o),
    .o(_al_u710_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u711 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[19]),
    .d(M_result2[18]),
    .o(_al_u711_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(C*A))"),
    .INIT(16'h004c))
    _al_u712 (
    .a(_al_u532_o),
    .b(_al_u711_o),
    .c(M_result2[17]),
    .d(_al_u525_o),
    .o(_al_u712_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u713 (
    .a(_al_u709_o),
    .b(_al_u710_o),
    .c(_al_u712_o),
    .d(M_result2[5]),
    .o(_al_u713_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u714 (
    .a(_al_u673_o),
    .b(_al_u701_o),
    .c(_al_u622_o),
    .d(M_result2[9]),
    .o(_al_u714_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u715 (
    .a(_al_u668_o),
    .b(M_result2[4]),
    .o(_al_u715_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(E*B)*~(D*A))"),
    .INIT(32'h0103050f))
    _al_u716 (
    .a(_al_u676_o),
    .b(_al_u714_o),
    .c(_al_u715_o),
    .d(M_result2[3]),
    .e(M_result2[2]),
    .o(_al_u716_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u717 (
    .a(_al_u569_o),
    .b(_al_u594_o),
    .c(M_result2[11]),
    .d(M_result2[8]),
    .o(_al_u717_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u718 (
    .a(_al_u716_o),
    .b(_al_u717_o),
    .c(_al_u600_o),
    .d(M_result2[9]),
    .o(_al_u718_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u719 (
    .a(M_result2[5]),
    .b(_al_u449_o),
    .c(_al_u483_o),
    .o(_al_u719_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u72 (
    .a(_al_u64_o),
    .b(n2[7]),
    .c(n2[6]),
    .o(n235_lutinv));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*(A*~(D)*~(E)+~(A)*D*E))"),
    .INIT(32'h04000008))
    _al_u720 (
    .a(_al_u426_o),
    .b(_al_u719_o),
    .c(M_result2[12]),
    .d(_al_u487_o),
    .e(_al_u489_o),
    .o(_al_u720_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*~A)"),
    .INIT(32'h00000001))
    _al_u721 (
    .a(_al_u666_o),
    .b(M_result2[9]),
    .c(M_result2[8]),
    .d(M_result2[7]),
    .e(M_result2[6]),
    .o(_al_u721_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*~A)"),
    .INIT(32'h00100000))
    _al_u722 (
    .a(_al_u531_o),
    .b(_al_u553_o),
    .c(_al_u720_o),
    .d(_al_u584_o),
    .e(_al_u721_o),
    .o(_al_u722_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u723 (
    .a(_al_u722_o),
    .b(_al_u565_o),
    .c(M_result2[12]),
    .d(M_result2[1]),
    .o(_al_u723_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u724 (
    .a(_al_u582_o),
    .b(_al_u560_o),
    .c(M_result2[13]),
    .d(M_result2[14]),
    .o(_al_u724_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u725 (
    .a(_al_u723_o),
    .b(_al_u724_o),
    .c(_al_u541_o),
    .d(M_result2[15]),
    .o(_al_u725_o));
  AL_MAP_LUT5 #(
    .EQN("(~(D*C*B)*~(E*~A))"),
    .INIT(32'h2aaa3fff))
    _al_u726 (
    .a(\NM/n4 [19]),
    .b(_al_u713_o),
    .c(_al_u718_o),
    .d(_al_u725_o),
    .e(_al_u525_o),
    .o(result[19]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u727 (
    .a(_al_u676_o),
    .b(M_result2[2]),
    .o(_al_u727_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u728 (
    .a(_al_u668_o),
    .b(M_result2[3]),
    .o(_al_u728_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*B))"),
    .INIT(16'h0105))
    _al_u729 (
    .a(_al_u727_o),
    .b(_al_u714_o),
    .c(_al_u728_o),
    .d(M_result2[1]),
    .o(_al_u729_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u73 (
    .a(_al_u64_o),
    .b(n2[5]),
    .c(n2[4]),
    .o(n237_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u730 (
    .a(_al_u722_o),
    .b(_al_u565_o),
    .c(M_result2[11]),
    .d(M_result[0]),
    .o(_al_u730_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u731 (
    .a(_al_u541_o),
    .b(_al_u560_o),
    .c(M_result2[14]),
    .d(M_result2[12]),
    .o(_al_u731_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u732 (
    .a(_al_u730_o),
    .b(_al_u731_o),
    .c(_al_u582_o),
    .d(M_result2[13]),
    .o(_al_u732_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u733 (
    .a(_al_u569_o),
    .b(_al_u594_o),
    .c(M_result2[10]),
    .d(M_result2[7]),
    .o(_al_u733_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E*D))"),
    .INIT(32'h00808080))
    _al_u734 (
    .a(_al_u729_o),
    .b(_al_u732_o),
    .c(_al_u733_o),
    .d(_al_u600_o),
    .e(M_result2[8]),
    .o(_al_u734_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u735 (
    .a(_al_u710_o),
    .b(_al_u586_o),
    .c(M_result2[9]),
    .d(M_result2[4]),
    .o(_al_u735_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u736 (
    .a(_al_u735_o),
    .b(_al_u624_o),
    .c(_al_u635_o),
    .d(M_result2[6]),
    .e(M_result2[5]),
    .o(_al_u736_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u737 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[17]),
    .d(M_result2[18]),
    .o(_al_u737_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(C*A))"),
    .INIT(16'h004c))
    _al_u738 (
    .a(_al_u532_o),
    .b(_al_u737_o),
    .c(M_result2[16]),
    .d(_al_u525_o),
    .o(_al_u738_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u739 (
    .a(_al_u736_o),
    .b(_al_u738_o),
    .c(_al_u535_o),
    .d(M_result2[15]),
    .o(_al_u739_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u74 (
    .a(n235_lutinv),
    .b(n237_lutinv),
    .c(_al_u67_o),
    .o(_al_u74_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u740 (
    .a(\NM/n4 [18]),
    .b(_al_u734_o),
    .c(_al_u739_o),
    .d(_al_u525_o),
    .o(result[18]));
  AL_MAP_LUT4 #(
    .EQN("(~B*(A*~(C)*~(D)+~(A)*C*D))"),
    .INIT(16'h1002))
    _al_u741 (
    .a(_al_u426_o),
    .b(M_result2[15]),
    .c(_al_u483_o),
    .d(_al_u489_o),
    .o(_al_u741_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u742 (
    .a(_al_u539_o),
    .b(_al_u741_o),
    .c(_al_u557_o),
    .d(_al_u567_o),
    .o(_al_u742_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u743 (
    .a(_al_u742_o),
    .b(_al_u531_o),
    .o(_al_u743_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u744 (
    .a(M_result2[9]),
    .b(M_result2[8]),
    .c(M_result2[7]),
    .d(M_result2[6]),
    .o(_al_u744_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u745 (
    .a(M_result2[5]),
    .b(M_result2[4]),
    .o(_al_u745_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u746 (
    .a(_al_u744_o),
    .b(_al_u745_o),
    .o(_al_u746_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u747 (
    .a(_al_u743_o),
    .b(_al_u746_o),
    .c(_al_u674_o),
    .d(M_result2[3]),
    .o(_al_u747_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u748 (
    .a(_al_u747_o),
    .b(_al_u722_o),
    .c(M_result2[2]),
    .d(M_result[0]),
    .o(_al_u748_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(D*C)*~(E*A))"),
    .INIT(32'h04440ccc))
    _al_u749 (
    .a(_al_u714_o),
    .b(_al_u748_o),
    .c(_al_u668_o),
    .d(M_result2[5]),
    .e(M_result2[3]),
    .o(_al_u749_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u75 (
    .a(n1[25]),
    .b(n2[25]),
    .o(\ADD01/ADD01/p2_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u750 (
    .a(_al_u624_o),
    .b(_al_u600_o),
    .c(M_result2[10]),
    .d(M_result2[8]),
    .o(_al_u750_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u751 (
    .a(_al_u750_o),
    .b(_al_u635_o),
    .c(M_result2[7]),
    .o(_al_u751_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u752 (
    .a(_al_u541_o),
    .b(_al_u565_o),
    .c(M_result2[16]),
    .d(M_result2[13]),
    .o(_al_u752_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*A))"),
    .INIT(8'h4c))
    _al_u753 (
    .a(_al_u676_o),
    .b(_al_u752_o),
    .c(M_result2[4]),
    .o(_al_u753_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E*D))"),
    .INIT(32'h00808080))
    _al_u754 (
    .a(_al_u749_o),
    .b(_al_u751_o),
    .c(_al_u753_o),
    .d(_al_u569_o),
    .e(M_result2[12]),
    .o(_al_u754_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u755 (
    .a(_al_u582_o),
    .b(_al_u560_o),
    .c(M_result2[15]),
    .d(M_result2[14]),
    .o(_al_u755_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u756 (
    .a(_al_u755_o),
    .b(_al_u535_o),
    .c(M_result2[17]),
    .o(_al_u756_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u757 (
    .a(_al_u586_o),
    .b(_al_u594_o),
    .c(M_result2[11]),
    .d(M_result2[9]),
    .o(_al_u757_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*~A))"),
    .INIT(16'h23af))
    _al_u758 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[19]),
    .d(M_result2[20]),
    .o(_al_u758_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(C*A))"),
    .INIT(16'h004c))
    _al_u759 (
    .a(_al_u532_o),
    .b(_al_u758_o),
    .c(M_result2[18]),
    .d(_al_u525_o),
    .o(_al_u759_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u76 (
    .a(\ADD01/ADD01/p2_lutinv ),
    .b(_al_u64_o),
    .c(n1[24]),
    .d(n2[24]),
    .o(\ADD01/ADD01/n10 ));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u760 (
    .a(_al_u757_o),
    .b(_al_u710_o),
    .c(_al_u759_o),
    .d(M_result2[6]),
    .o(_al_u760_o));
  AL_MAP_LUT5 #(
    .EQN("(~(D*C*B)*~(E*~A))"),
    .INIT(32'h2aaa3fff))
    _al_u761 (
    .a(\NM/n4 [20]),
    .b(_al_u754_o),
    .c(_al_u756_o),
    .d(_al_u760_o),
    .e(_al_u525_o),
    .o(result[20]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u762 (
    .a(_al_u624_o),
    .b(_al_u569_o),
    .c(M_result2[13]),
    .d(M_result2[9]),
    .o(_al_u762_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u763 (
    .a(_al_u762_o),
    .b(_al_u600_o),
    .c(_al_u594_o),
    .d(M_result2[11]),
    .e(M_result2[10]),
    .o(_al_u763_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hbd9f))
    _al_u764 (
    .a(_al_u426_o),
    .b(_al_u475_o),
    .c(_al_u473_o),
    .d(_al_u428_o),
    .o(_al_u764_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*A)"),
    .INIT(16'h0080))
    _al_u765 (
    .a(_al_u743_o),
    .b(_al_u746_o),
    .c(_al_u674_o),
    .d(_al_u764_o),
    .o(_al_u765_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u766 (
    .a(_al_u747_o),
    .b(_al_u765_o),
    .c(M_result2[1]),
    .d(M_result[0]),
    .o(_al_u766_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u767 (
    .a(_al_u763_o),
    .b(_al_u766_o),
    .c(_al_u722_o),
    .d(M_result2[3]),
    .o(_al_u767_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u768 (
    .a(_al_u676_o),
    .b(_al_u714_o),
    .c(M_result2[5]),
    .d(M_result2[4]),
    .o(_al_u768_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u769 (
    .a(_al_u582_o),
    .b(_al_u565_o),
    .c(M_result2[16]),
    .d(M_result2[14]),
    .o(_al_u769_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(C)*~((~D*B))+~(A)*C*~((~D*B))+A*C*~((~D*B))+~(A)*C*(~D*B))"),
    .INIT(16'hf571))
    _al_u77 (
    .a(n1[29]),
    .b(n1[28]),
    .c(n2[29]),
    .d(n2[28]),
    .o(_al_u77_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(E*D))"),
    .INIT(32'h00808080))
    _al_u770 (
    .a(_al_u767_o),
    .b(_al_u768_o),
    .c(_al_u769_o),
    .d(_al_u668_o),
    .e(M_result2[6]),
    .o(_al_u770_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~A*~(D*B)))"),
    .INIT(16'he0a0))
    _al_u771 (
    .a(_al_u541_o),
    .b(_al_u559_o),
    .c(M_result2[17]),
    .d(M_result2[15]),
    .o(_al_u771_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u772 (
    .a(_al_u528_o),
    .b(M_result2[23]),
    .c(M_result2[21]),
    .d(M_result2[20]),
    .o(_al_u772_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(C*A))"),
    .INIT(16'h004c))
    _al_u773 (
    .a(_al_u532_o),
    .b(_al_u772_o),
    .c(M_result2[19]),
    .d(_al_u525_o),
    .o(_al_u773_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(D*B))"),
    .INIT(16'h1050))
    _al_u774 (
    .a(_al_u771_o),
    .b(_al_u710_o),
    .c(_al_u773_o),
    .d(M_result2[7]),
    .o(_al_u774_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u775 (
    .a(_al_u635_o),
    .b(_al_u586_o),
    .c(M_result2[12]),
    .d(M_result2[8]),
    .o(_al_u775_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u776 (
    .a(_al_u774_o),
    .b(_al_u775_o),
    .c(_al_u535_o),
    .d(M_result2[18]),
    .o(_al_u776_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u777 (
    .a(\NM/n4 [21]),
    .b(_al_u770_o),
    .c(_al_u776_o),
    .d(_al_u525_o),
    .o(result[21]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u778 (
    .a(M_result2[3]),
    .b(M_result2[2]),
    .o(_al_u778_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u779 (
    .a(_al_u721_o),
    .b(_al_u745_o),
    .c(_al_u778_o),
    .d(M_result2[1]),
    .e(M_result[0]),
    .o(_al_u779_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*B*~(C)+~(A)*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'hd4))
    _al_u78 (
    .a(n1[30]),
    .b(n2[30]),
    .c(_al_u77_o),
    .o(_al_u78_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u780 (
    .a(_al_u699_o),
    .b(_al_u535_o),
    .c(_al_u779_o),
    .d(M_result2[19]),
    .o(_al_u780_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*~(~B*~(D*C))))"),
    .INIT(32'h0222aaaa))
    _al_u781 (
    .a(_al_u780_o),
    .b(_al_u541_o),
    .c(_al_u566_o),
    .d(M_result2[17]),
    .e(M_result2[18]),
    .o(_al_u781_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u782 (
    .a(_al_u600_o),
    .b(_al_u594_o),
    .c(M_result2[12]),
    .d(M_result2[11]),
    .o(_al_u782_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D))"),
    .INIT(32'h00001b1f))
    _al_u783 (
    .a(M_result2[23]),
    .b(M_result2[21]),
    .c(M_result2[22]),
    .d(M_result2[20]),
    .e(_al_u525_o),
    .o(_al_u783_o));
  AL_MAP_LUT5 #(
    .EQN("(D*B*A*~(E*C))"),
    .INIT(32'h08008800))
    _al_u784 (
    .a(_al_u781_o),
    .b(_al_u782_o),
    .c(_al_u710_o),
    .d(_al_u783_o),
    .e(M_result2[8]),
    .o(_al_u784_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u785 (
    .a(_al_u624_o),
    .b(_al_u569_o),
    .c(M_result2[14]),
    .d(M_result2[10]),
    .o(_al_u785_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u786 (
    .a(_al_u785_o),
    .b(_al_u635_o),
    .c(_al_u586_o),
    .d(M_result2[13]),
    .e(M_result2[9]),
    .o(_al_u786_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u787 (
    .a(_al_u714_o),
    .b(_al_u722_o),
    .c(M_result2[5]),
    .d(M_result2[4]),
    .o(_al_u787_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u788 (
    .a(_al_u747_o),
    .b(_al_u765_o),
    .c(M_result2[2]),
    .d(M_result2[1]),
    .o(_al_u788_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u789 (
    .a(_al_u784_o),
    .b(_al_u786_o),
    .c(_al_u787_o),
    .d(_al_u788_o),
    .o(_al_u789_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u79 (
    .a(n1[29]),
    .b(n1[28]),
    .c(n2[29]),
    .d(n2[28]),
    .o(\ADD01/ADD02/n7 ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u790 (
    .a(_al_u560_o),
    .b(_al_u565_o),
    .c(M_result2[16]),
    .d(M_result2[15]),
    .o(_al_u790_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(D*C)*~(E*A))"),
    .INIT(32'h04440ccc))
    _al_u791 (
    .a(_al_u676_o),
    .b(_al_u790_o),
    .c(_al_u668_o),
    .d(M_result2[7]),
    .e(M_result2[6]),
    .o(_al_u791_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u792 (
    .a(\NM/n4 [22]),
    .b(_al_u789_o),
    .c(_al_u791_o),
    .d(_al_u525_o),
    .o(result[22]));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(~C*~(D*~B)))"),
    .INIT(16'h5150))
    _al_u793 (
    .a(M_result2[21]),
    .b(_al_u549_o),
    .c(M_result2[20]),
    .d(M_result2[18]),
    .o(_al_u793_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~C*~(~E*~D*~A)))"),
    .INIT(32'hc0c0c0c4))
    _al_u794 (
    .a(_al_u793_o),
    .b(_al_u528_o),
    .c(_al_u531_o),
    .d(_al_u565_o),
    .e(_al_u586_o),
    .o(_al_u794_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*~(~E*~D*~C))"),
    .INIT(32'h22222220))
    _al_u795 (
    .a(_al_u638_o),
    .b(_al_u531_o),
    .c(_al_u667_o),
    .d(_al_u634_o),
    .e(_al_u594_o),
    .o(_al_u795_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u796 (
    .a(_al_u745_o),
    .b(_al_u778_o),
    .c(M_result2[1]),
    .d(M_result[0]),
    .o(_al_u796_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*~C*B*~A)"),
    .INIT(32'h04000000))
    _al_u797 (
    .a(_al_u531_o),
    .b(_al_u697_o),
    .c(_al_u539_o),
    .d(_al_u796_o),
    .e(_al_u721_o),
    .o(_al_u797_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*~B*A)"),
    .INIT(32'h00000002))
    _al_u798 (
    .a(_al_u794_o),
    .b(_al_u795_o),
    .c(_al_u797_o),
    .d(_al_u714_o),
    .e(_al_u765_o),
    .o(_al_u798_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u799 (
    .a(_al_u103_o),
    .b(n1[23]),
    .c(n2[23]),
    .o(E[0]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u80 (
    .a(n1[30]),
    .b(n2[30]),
    .o(\ADD01/ADD02/p3_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("~(C@(~B*A))"),
    .INIT(8'h2d))
    _al_u800 (
    .a(_al_u798_o),
    .b(_al_u525_o),
    .c(E[0]),
    .o(\ADD03/ADD01/p0_neg ));
  AL_MAP_LUT5 #(
    .EQN("(~C*~B*~(D*~(~E*A)))"),
    .INIT(32'h00030203))
    _al_u801 (
    .a(_al_u665_o),
    .b(M_result2[15]),
    .c(_al_u622_o),
    .d(_al_u640_o),
    .e(_al_u666_o),
    .o(_al_u801_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u802 (
    .a(_al_u638_o),
    .b(_al_u531_o),
    .c(_al_u801_o),
    .o(_al_u802_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~A*~(D*~(~E*B)))"),
    .INIT(32'h00050405))
    _al_u803 (
    .a(_al_u567_o),
    .b(M_result2[13]),
    .c(M_result2[15]),
    .d(_al_u593_o),
    .e(_al_u599_o),
    .o(_al_u803_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~C*~(~D*~(~E*~B))))"),
    .INIT(32'h50555054))
    _al_u804 (
    .a(_al_u531_o),
    .b(_al_u803_o),
    .c(_al_u539_o),
    .d(_al_u557_o),
    .e(_al_u567_o),
    .o(_al_u804_o));
  AL_MAP_LUT5 #(
    .EQN("(C*B*A*~(~E*~D))"),
    .INIT(32'h80808000))
    _al_u805 (
    .a(_al_u721_o),
    .b(_al_u745_o),
    .c(_al_u778_o),
    .d(M_result2[1]),
    .e(M_result[0]),
    .o(_al_u805_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u806 (
    .a(_al_u531_o),
    .b(_al_u805_o),
    .c(_al_u697_o),
    .o(_al_u806_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~D*~C*~B*~A))"),
    .INIT(32'h0000fffe))
    _al_u807 (
    .a(_al_u802_o),
    .b(_al_u804_o),
    .c(_al_u806_o),
    .d(_al_u722_o),
    .e(_al_u525_o),
    .o(_al_u807_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u808 (
    .a(_al_u525_o),
    .b(E[0]),
    .o(_al_u808_o));
  AL_MAP_LUT5 #(
    .EQN("((D*~(E)*~(C)+D*E*~(C)+~(D)*E*C+D*E*C)@(B*A))"),
    .INIT(32'h77788788))
    _al_u809 (
    .a(_al_u525_o),
    .b(E[0]),
    .c(_al_u103_o),
    .d(n1[24]),
    .e(n2[24]),
    .o(_al_u809_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u81 (
    .a(n1[27]),
    .b(n2[27]),
    .o(\ADD01/ADD02/g0 ));
  AL_MAP_LUT4 #(
    .EQN("(D@B@(C*~A))"),
    .INIT(16'h639c))
    _al_u810 (
    .a(_al_u798_o),
    .b(_al_u807_o),
    .c(_al_u808_o),
    .d(_al_u809_o),
    .o(result[24]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u811 (
    .a(_al_u721_o),
    .b(_al_u745_o),
    .c(_al_u778_o),
    .d(M_result2[12]),
    .o(_al_u811_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(~D*~C))"),
    .INIT(16'h2220))
    _al_u812 (
    .a(_al_u698_o),
    .b(_al_u531_o),
    .c(_al_u805_o),
    .d(_al_u811_o),
    .o(_al_u812_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~B*~(~D*~A))"),
    .INIT(16'h0302))
    _al_u813 (
    .a(_al_u634_o),
    .b(_al_u531_o),
    .c(_al_u539_o),
    .d(_al_u623_o),
    .o(_al_u813_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~A*~(~E*~D*~B))"),
    .INIT(32'h05050504))
    _al_u814 (
    .a(_al_u531_o),
    .b(_al_u801_o),
    .c(_al_u539_o),
    .d(_al_u557_o),
    .e(_al_u567_o),
    .o(_al_u814_o));
  AL_MAP_LUT4 #(
    .EQN("(A*(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'ha820))
    _al_u815 (
    .a(E[0]),
    .b(_al_u103_o),
    .c(n1[24]),
    .d(n2[24]),
    .o(\ADD0212/ADD01/n1 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u816 (
    .a(_al_u103_o),
    .b(n1[25]),
    .c(n2[25]),
    .o(E[2]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'h78))
    _al_u817 (
    .a(_al_u525_o),
    .b(\ADD0212/ADD01/n1 ),
    .c(E[2]),
    .o(_al_u817_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@(~E*~(~C*~B*~A)))"),
    .INIT(32'h00fffe01))
    _al_u818 (
    .a(_al_u812_o),
    .b(_al_u813_o),
    .c(_al_u814_o),
    .d(_al_u817_o),
    .e(_al_u525_o),
    .o(_al_u818_o));
  AL_MAP_LUT5 #(
    .EQN("(B@(~(C)*~((D*~A))*~(E)+~(C)*~((D*~A))*E+C*~((D*~A))*E+~(C)*(D*~A)*E))"),
    .INIT(32'h6333c6c3))
    _al_u819 (
    .a(_al_u798_o),
    .b(_al_u818_o),
    .c(_al_u807_o),
    .d(_al_u808_o),
    .e(_al_u809_o),
    .o(result[25]));
  AL_MAP_LUT5 #(
    .EQN("(B*~A*~(E*D*C))"),
    .INIT(32'h04444444))
    _al_u82 (
    .a(\ADD01/ADD01/n10 ),
    .b(_al_u78_o),
    .c(\ADD01/ADD02/n7 ),
    .d(\ADD01/ADD02/p3_lutinv ),
    .e(\ADD01/ADD02/g0 ),
    .o(_al_u82_o));
  AL_MAP_LUT4 #(
    .EQN("(~(B)*~((C*~A))*~(D)+~(B)*~((C*~A))*D+B*~((C*~A))*D+~(B)*(C*~A)*D)"),
    .INIT(16'hbf23))
    _al_u820 (
    .a(_al_u798_o),
    .b(_al_u807_o),
    .c(_al_u808_o),
    .d(_al_u809_o),
    .o(_al_u820_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u821 (
    .a(_al_u634_o),
    .b(_al_u623_o),
    .o(_al_u821_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~A*~(C*~B)))"),
    .INIT(16'h00ba))
    _al_u822 (
    .a(_al_u700_o),
    .b(_al_u821_o),
    .c(_al_u620_o),
    .d(_al_u531_o),
    .o(_al_u822_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*~B))"),
    .INIT(16'h4555))
    _al_u823 (
    .a(_al_u668_o),
    .b(_al_u531_o),
    .c(_al_u558_o),
    .d(_al_u803_o),
    .o(_al_u823_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*~B))"),
    .INIT(8'ha8))
    _al_u824 (
    .a(_al_u566_o),
    .b(_al_u585_o),
    .c(_al_u568_o),
    .o(_al_u824_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u825 (
    .a(\ADD0212/ADD01/n1 ),
    .b(E[2]),
    .o(\ADD0212/ADD01/n8 ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u826 (
    .a(_al_u103_o),
    .b(n1[26]),
    .c(n2[26]),
    .o(E[3]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'h78))
    _al_u827 (
    .a(_al_u525_o),
    .b(\ADD0212/ADD01/n8 ),
    .c(E[3]),
    .o(_al_u827_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@(~E*~(~C*B*~A)))"),
    .INIT(32'h00fffb04))
    _al_u828 (
    .a(_al_u822_o),
    .b(_al_u823_o),
    .c(_al_u824_o),
    .d(_al_u827_o),
    .e(_al_u525_o),
    .o(_al_u828_o));
  AL_MAP_LUT5 #(
    .EQN("(D*~(~E*~(~C*~B*~A)))"),
    .INIT(32'hff000100))
    _al_u829 (
    .a(_al_u812_o),
    .b(_al_u813_o),
    .c(_al_u814_o),
    .d(_al_u817_o),
    .e(_al_u525_o),
    .o(_al_u829_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(C)*~((D*~B))+A*~(C)*~((D*~B))+A*C*~((D*~B))+A*~(C)*(D*~B))"),
    .INIT(16'h8eaf))
    _al_u83 (
    .a(n1[24]),
    .b(n1[23]),
    .c(n2[24]),
    .d(n2[23]),
    .o(\ADD01/ADD01/c1_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~(~C*~B*~A))"),
    .INIT(32'h000000fe))
    _al_u830 (
    .a(_al_u812_o),
    .b(_al_u813_o),
    .c(_al_u814_o),
    .d(_al_u525_o),
    .e(E[2]),
    .o(_al_u830_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(~C*~(~D*A)))"),
    .INIT(16'h3c36))
    _al_u831 (
    .a(_al_u820_o),
    .b(_al_u828_o),
    .c(_al_u829_o),
    .d(_al_u830_o),
    .o(result[26]));
  AL_MAP_LUT5 #(
    .EQN("(B*(~(C)*~((D*~A))*~(E)+~(C)*~((D*~A))*E+C*~((D*~A))*E+~(C)*(D*~A)*E))"),
    .INIT(32'h8ccc080c))
    _al_u832 (
    .a(_al_u798_o),
    .b(_al_u818_o),
    .c(_al_u807_o),
    .d(_al_u808_o),
    .e(_al_u809_o),
    .o(_al_u832_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*~(~D*~(~E*~A)))"),
    .INIT(32'h30003010))
    _al_u833 (
    .a(_al_u821_o),
    .b(_al_u531_o),
    .c(_al_u558_o),
    .d(_al_u803_o),
    .e(M_result2[17]),
    .o(_al_u833_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~D*~C*~A))"),
    .INIT(16'h3332))
    _al_u834 (
    .a(_al_u833_o),
    .b(_al_u525_o),
    .c(_al_u824_o),
    .d(_al_u802_o),
    .o(_al_u834_o));
  AL_MAP_LUT5 #(
    .EQN("(D*C*~B*~(~E*~A))"),
    .INIT(32'h30002000))
    _al_u835 (
    .a(_al_u675_o),
    .b(_al_u531_o),
    .c(_al_u558_o),
    .d(_al_u592_o),
    .e(_al_u714_o),
    .o(_al_u835_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u836 (
    .a(_al_u103_o),
    .b(n1[27]),
    .c(n2[27]),
    .o(E[4]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*B*A))"),
    .INIT(16'h7f80))
    _al_u837 (
    .a(_al_u525_o),
    .b(\ADD0212/ADD01/n8 ),
    .c(E[3]),
    .d(E[4]),
    .o(_al_u837_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@(~E*~(~C*~B*~A)))"),
    .INIT(32'h00fffe01))
    _al_u838 (
    .a(_al_u812_o),
    .b(_al_u835_o),
    .c(_al_u722_o),
    .d(_al_u837_o),
    .e(_al_u525_o),
    .o(_al_u838_o));
  AL_MAP_LUT5 #(
    .EQN("(D@(~(B)*~((~C*~A))*~(E)+~(B)*~((~C*~A))*E+B*~((~C*~A))*E+~(B)*(~C*~A)*E))"),
    .INIT(32'h04fbcd32))
    _al_u839 (
    .a(_al_u832_o),
    .b(_al_u834_o),
    .c(_al_u829_o),
    .d(_al_u838_o),
    .e(_al_u827_o),
    .o(result[27]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u84 (
    .a(n1[26]),
    .b(n2[26]),
    .o(\ADD01/ADD01/p3_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(D*(~(B)*~((~C*~A))*~(E)+~(B)*~((~C*~A))*E+B*~((~C*~A))*E+~(B)*(~C*~A)*E))"),
    .INIT(32'hfb003200))
    _al_u840 (
    .a(_al_u832_o),
    .b(_al_u834_o),
    .c(_al_u829_o),
    .d(_al_u838_o),
    .e(_al_u827_o),
    .o(_al_u840_o));
  AL_MAP_LUT5 #(
    .EQN("(D*~(~E*~(~C*~B*~A)))"),
    .INIT(32'hff000100))
    _al_u841 (
    .a(_al_u812_o),
    .b(_al_u835_o),
    .c(_al_u722_o),
    .d(_al_u837_o),
    .e(_al_u525_o),
    .o(_al_u841_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u842 (
    .a(E[3]),
    .b(E[4]),
    .o(_al_u842_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u843 (
    .a(_al_u103_o),
    .b(n1[28]),
    .c(n2[28]),
    .o(E[5]));
  AL_MAP_LUT4 #(
    .EQN("(D@(C*B*A))"),
    .INIT(16'h7f80))
    _al_u844 (
    .a(_al_u525_o),
    .b(\ADD0212/ADD01/n8 ),
    .c(_al_u842_o),
    .d(E[5]),
    .o(_al_u844_o));
  AL_MAP_LUT3 #(
    .EQN("(C@(~B*~A))"),
    .INIT(8'he1))
    _al_u845 (
    .a(_al_u840_o),
    .b(_al_u841_o),
    .c(_al_u844_o),
    .o(result[28]));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u846 (
    .a(_al_u525_o),
    .b(\ADD0212/ADD01/n8 ),
    .c(_al_u842_o),
    .d(E[5]),
    .o(_al_u846_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u847 (
    .a(_al_u846_o),
    .b(n2[29]),
    .o(_al_u847_o));
  AL_MAP_LUT3 #(
    .EQN("~(A@(~C*~B))"),
    .INIT(8'h56))
    _al_u848 (
    .a(_al_u847_o),
    .b(n1[30]),
    .c(n2[30]),
    .o(_al_u848_o));
  AL_MAP_LUT4 #(
    .EQN("(A@(C*~(D)*~(B)+C*D*~(B)+~(C)*D*B+C*D*B))"),
    .INIT(16'h569a))
    _al_u849 (
    .a(_al_u846_o),
    .b(_al_u103_o),
    .c(n1[29]),
    .d(n2[29]),
    .o(_al_u849_o));
  AL_MAP_LUT4 #(
    .EQN("(B@(~(A)*~(C)*~(D)+~(A)*~(C)*D+A*~(C)*D+~(A)*C*D))"),
    .INIT(16'h93c9))
    _al_u85 (
    .a(\ADD01/ADD01/c1_lutinv ),
    .b(\ADD01/ADD01/p3_lutinv ),
    .c(n1[25]),
    .d(n2[25]),
    .o(\C023/outtemp [3]));
  AL_MAP_LUT5 #(
    .EQN("(C@(~E*~D*~B*~A))"),
    .INIT(32'hf0f0f0e1))
    _al_u850 (
    .a(_al_u840_o),
    .b(_al_u841_o),
    .c(_al_u848_o),
    .d(_al_u849_o),
    .e(_al_u844_o),
    .o(result[30]));
  AL_MAP_LUT4 #(
    .EQN("(C@(~D*~B*~A))"),
    .INIT(16'hf0e1))
    _al_u851 (
    .a(_al_u840_o),
    .b(_al_u841_o),
    .c(_al_u849_o),
    .d(_al_u844_o),
    .o(result[29]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*B*C*D*E)"),
    .INIT(32'h80ecc8fe))
    _al_u86 (
    .a(\ADD01/ADD01/c1_lutinv ),
    .b(n1[26]),
    .c(n1[25]),
    .d(n2[26]),
    .e(n2[25]),
    .o(\ADD01/ctemp_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u87 (
    .a(n1[28]),
    .b(n2[28]),
    .o(\ADD01/ADD02/p1_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u88 (
    .a(\ADD01/ADD02/p1_lutinv ),
    .b(n1[30]),
    .c(n1[29]),
    .d(n2[30]),
    .e(n2[29]),
    .o(\ADD01/ADD02/n17 ));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u89 (
    .a(n1[27]),
    .b(n2[27]),
    .o(\ADD01/ADD02/p0_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("~(B@(A*~(E*D*C)))"),
    .INIT(32'h39999999))
    _al_u90 (
    .a(_al_u82_o),
    .b(\C023/outtemp [3]),
    .c(\ADD01/ctemp_lutinv ),
    .d(\ADD01/ADD02/n17 ),
    .e(\ADD01/ADD02/p0_lutinv ),
    .o(exp_diff[3]));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u91 (
    .a(n1[24]),
    .b(n1[23]),
    .c(n2[24]),
    .d(n2[23]),
    .o(\ADD01/ADD01/n3 ));
  AL_MAP_LUT5 #(
    .EQN("(~C*A*~(E*D*B))"),
    .INIT(32'h020a0a0a))
    _al_u92 (
    .a(_al_u78_o),
    .b(\ADD01/ADD02/n7 ),
    .c(\ADD01/ADD01/n3 ),
    .d(\ADD01/ADD02/p3_lutinv ),
    .e(\ADD01/ADD02/g0 ),
    .o(_al_u92_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u93 (
    .a(\ADD01/ADD01/c1_lutinv ),
    .b(\ADD01/ADD01/p2_lutinv ),
    .o(_al_u93_o));
  AL_MAP_LUT5 #(
    .EQN("(C@(A*~(E*D*B)))"),
    .INIT(32'hd25a5a5a))
    _al_u94 (
    .a(_al_u92_o),
    .b(\ADD01/ctemp_lutinv ),
    .c(_al_u93_o),
    .d(\ADD01/ADD02/n17 ),
    .e(\ADD01/ADD02/p0_lutinv ),
    .o(exp_diff[2]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haaf0ccff))
    _al_u95 (
    .a(_al_u68_o),
    .b(_al_u71_o),
    .c(_al_u74_o),
    .d(exp_diff[3]),
    .e(exp_diff[2]),
    .o(_al_u95_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u96 (
    .a(_al_u64_o),
    .b(n2[22]),
    .o(_al_u96_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u97 (
    .a(_al_u64_o),
    .b(n2[21]),
    .c(n2[20]),
    .o(n221_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u98 (
    .a(_al_u96_o),
    .b(n221_lutinv),
    .c(_al_u67_o),
    .o(_al_u98_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u99 (
    .a(_al_u64_o),
    .b(n2[19]),
    .c(n2[18]),
    .o(n223_lutinv));

endmodule 

module add_sub  // ../RTL/core/fpu.v(83)
  (
  n1,
  n2,
  sub,
  Exception,
  Overflow,
  Underflow,
  result
  );

  input [31:0] n1;  // ../RTL/core/fpu.v(84)
  input [31:0] n2;  // ../RTL/core/fpu.v(85)
  input sub;  // ../RTL/core/fpu.v(87)
  output Exception;  // ../RTL/core/fpu.v(90)
  output Overflow;  // ../RTL/core/fpu.v(88)
  output Underflow;  // ../RTL/core/fpu.v(89)
  output [31:0] result;  // ../RTL/core/fpu.v(86)

  wire [7:0] \C023/outtemp ;  // ../RTL/core/fpu_utils.v(93)
  wire [7:0] E;  // ../RTL/core/fpu.v(95)
  wire [23:0] M1;  // ../RTL/core/fpu.v(97)
  wire [23:0] M_result;  // ../RTL/core/fpu.v(97)
  wire [23:0] M_result2;  // ../RTL/core/fpu.v(97)
  wire [22:0] \NM/n4 ;
  wire [7:0] exp_diff;  // ../RTL/core/fpu.v(95)
  wire [23:0] new_M2;  // ../RTL/core/fpu.v(97)
  wire \ADD01/ADD01/c1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD01/n20 ;
  wire \ADD01/ADD01/n3 ;
  wire \ADD01/ADD01/n7 ;
  wire \ADD01/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/n17 ;
  wire \ADD01/ADD02/n3 ;
  wire \ADD01/ADD02/p0_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ADD02/p1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD01/ctemp_lutinv ;  // ../RTL/core/fpu_utils.v(76)
  wire \ADD02/ADD01/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD01/p3_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/n3 ;
  wire \ADD02/ADD01/ADD02/p0_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/p1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD01/ADD02/p2_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/g2 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/n1 ;
  wire \ADD02/ADD02/ADD01/n3 ;
  wire \ADD02/ADD02/ADD01/p0_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/p1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD01/p2_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/n10 ;
  wire \ADD02/ADD02/ADD02/p0_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/p1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/p2_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD02/ADD02/p3_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/n14 ;
  wire \ADD02/ADD03/ADD01/n3 ;
  wire \ADD02/ADD03/ADD01/p0_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/p1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/p2_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD01/p3_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g0 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g1 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/g3 ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/n18 ;
  wire \ADD02/ADD03/ADD02/n20 ;
  wire \ADD02/ADD03/ADD02/n3 ;
  wire \ADD02/ADD03/ADD02/n6_lutinv ;
  wire \ADD02/ADD03/ADD02/p0_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/p1_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/p2_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD02/ADD03/ADD02/p3_lutinv ;  // ../RTL/core/fpu_utils.v(54)
  wire \ADD03/ADD01/p0_neg ;
  wire \C023/ADD01/ADD02/n0 ;
  wire \M04/M01/M01/invSL_lutinv ;  // ../RTL/core/fpu_utils.v(105)
  wire \NM/add0/c11 ;  // ../RTL/core/fpu_utils.v(158)
  wire \NM/add0/c15 ;  // ../RTL/core/fpu_utils.v(158)
  wire \NM/add0/c19 ;  // ../RTL/core/fpu_utils.v(158)
  wire \NM/add0/c3 ;  // ../RTL/core/fpu_utils.v(158)
  wire \NM/add0/c7 ;  // ../RTL/core/fpu_utils.v(158)
  wire _al_u102_o;
  wire _al_u103_o;
  wire _al_u104_o;
  wire _al_u105_o;
  wire _al_u108_o;
  wire _al_u109_o;
  wire _al_u110_o;
  wire _al_u112_o;
  wire _al_u114_o;
  wire _al_u115_o;
  wire _al_u116_o;
  wire _al_u117_o;
  wire _al_u120_o;
  wire _al_u123_o;
  wire _al_u124_o;
  wire _al_u127_o;
  wire _al_u129_o;
  wire _al_u130_o;
  wire _al_u131_o;
  wire _al_u132_o;
  wire _al_u134_o;
  wire _al_u137_o;
  wire _al_u138_o;
  wire _al_u139_o;
  wire _al_u140_o;
  wire _al_u141_o;
  wire _al_u142_o;
  wire _al_u144_o;
  wire _al_u145_o;
  wire _al_u148_o;
  wire _al_u150_o;
  wire _al_u151_o;
  wire _al_u152_o;
  wire _al_u155_o;
  wire _al_u156_o;
  wire _al_u159_o;
  wire _al_u160_o;
  wire _al_u163_o;
  wire _al_u166_o;
  wire _al_u167_o;
  wire _al_u168_o;
  wire _al_u169_o;
  wire _al_u170_o;
  wire _al_u171_o;
  wire _al_u173_o;
  wire _al_u174_o;
  wire _al_u177_o;
  wire _al_u178_o;
  wire _al_u180_o;
  wire _al_u183_o;
  wire _al_u184_o;
  wire _al_u187_o;
  wire _al_u190_o;
  wire _al_u191_o;
  wire _al_u192_o;
  wire _al_u193_o;
  wire _al_u195_o;
  wire _al_u196_o;
  wire _al_u197_o;
  wire _al_u198_o;
  wire _al_u199_o;
  wire _al_u200_o;
  wire _al_u201_o;
  wire _al_u202_o;
  wire _al_u203_o;
  wire _al_u205_o;
  wire _al_u206_o;
  wire _al_u207_o;
  wire _al_u209_o;
  wire _al_u210_o;
  wire _al_u211_o;
  wire _al_u212_o;
  wire _al_u213_o;
  wire _al_u214_o;
  wire _al_u215_o;
  wire _al_u216_o;
  wire _al_u217_o;
  wire _al_u218_o;
  wire _al_u220_o;
  wire _al_u221_o;
  wire _al_u222_o;
  wire _al_u223_o;
  wire _al_u224_o;
  wire _al_u225_o;
  wire _al_u226_o;
  wire _al_u227_o;
  wire _al_u228_o;
  wire _al_u229_o;
  wire _al_u231_o;
  wire _al_u232_o;
  wire _al_u233_o;
  wire _al_u234_o;
  wire _al_u235_o;
  wire _al_u236_o;
  wire _al_u237_o;
  wire _al_u238_o;
  wire _al_u239_o;
  wire _al_u240_o;
  wire _al_u241_o;
  wire _al_u242_o;
  wire _al_u243_o;
  wire _al_u244_o;
  wire _al_u245_o;
  wire _al_u246_o;
  wire _al_u247_o;
  wire _al_u248_o;
  wire _al_u249_o;
  wire _al_u250_o;
  wire _al_u251_o;
  wire _al_u253_o;
  wire _al_u254_o;
  wire _al_u255_o;
  wire _al_u257_o;
  wire _al_u258_o;
  wire _al_u259_o;
  wire _al_u261_o;
  wire _al_u262_o;
  wire _al_u263_o;
  wire _al_u264_o;
  wire _al_u265_o;
  wire _al_u266_o;
  wire _al_u267_o;
  wire _al_u268_o;
  wire _al_u269_o;
  wire _al_u270_o;
  wire _al_u271_o;
  wire _al_u272_o;
  wire _al_u274_o;
  wire _al_u275_o;
  wire _al_u276_o;
  wire _al_u277_o;
  wire _al_u278_o;
  wire _al_u279_o;
  wire _al_u281_o;
  wire _al_u282_o;
  wire _al_u284_o;
  wire _al_u285_o;
  wire _al_u286_o;
  wire _al_u287_o;
  wire _al_u288_o;
  wire _al_u289_o;
  wire _al_u290_o;
  wire _al_u291_o;
  wire _al_u292_o;
  wire _al_u294_o;
  wire _al_u296_o;
  wire _al_u297_o;
  wire _al_u298_o;
  wire _al_u299_o;
  wire _al_u300_o;
  wire _al_u301_o;
  wire _al_u302_o;
  wire _al_u303_o;
  wire _al_u304_o;
  wire _al_u306_o;
  wire _al_u307_o;
  wire _al_u308_o;
  wire _al_u310_o;
  wire _al_u311_o;
  wire _al_u315_o;
  wire _al_u316_o;
  wire _al_u317_o;
  wire _al_u318_o;
  wire _al_u319_o;
  wire _al_u320_o;
  wire _al_u321_o;
  wire _al_u322_o;
  wire _al_u323_o;
  wire _al_u328_o;
  wire _al_u329_o;
  wire _al_u330_o;
  wire _al_u331_o;
  wire _al_u332_o;
  wire _al_u333_o;
  wire _al_u334_o;
  wire _al_u335_o;
  wire _al_u336_o;
  wire _al_u337_o;
  wire _al_u338_o;
  wire _al_u339_o;
  wire _al_u341_o;
  wire _al_u342_o;
  wire _al_u343_o;
  wire _al_u345_o;
  wire _al_u347_o;
  wire _al_u348_o;
  wire _al_u349_o;
  wire _al_u350_o;
  wire _al_u351_o;
  wire _al_u352_o;
  wire _al_u353_o;
  wire _al_u354_o;
  wire _al_u355_o;
  wire _al_u356_o;
  wire _al_u358_o;
  wire _al_u359_o;
  wire _al_u360_o;
  wire _al_u362_o;
  wire _al_u363_o;
  wire _al_u364_o;
  wire _al_u365_o;
  wire _al_u366_o;
  wire _al_u368_o;
  wire _al_u369_o;
  wire _al_u370_o;
  wire _al_u371_o;
  wire _al_u374_o;
  wire _al_u375_o;
  wire _al_u377_o;
  wire _al_u378_o;
  wire _al_u380_o;
  wire _al_u381_o;
  wire _al_u382_o;
  wire _al_u384_o;
  wire _al_u386_o;
  wire _al_u387_o;
  wire _al_u388_o;
  wire _al_u390_o;
  wire _al_u391_o;
  wire _al_u393_o;
  wire _al_u395_o;
  wire _al_u397_o;
  wire _al_u400_o;
  wire _al_u401_o;
  wire _al_u403_o;
  wire _al_u404_o;
  wire _al_u406_o;
  wire _al_u407_o;
  wire _al_u408_o;
  wire _al_u409_o;
  wire _al_u410_o;
  wire _al_u412_o;
  wire _al_u413_o;
  wire _al_u415_o;
  wire _al_u416_o;
  wire _al_u423_o;
  wire _al_u427_o;
  wire _al_u428_o;
  wire _al_u430_o;
  wire _al_u431_o;
  wire _al_u432_o;
  wire _al_u433_o;
  wire _al_u434_o;
  wire _al_u435_o;
  wire _al_u438_o;
  wire _al_u440_o;
  wire _al_u442_o;
  wire _al_u443_o;
  wire _al_u444_o;
  wire _al_u446_o;
  wire _al_u448_o;
  wire _al_u449_o;
  wire _al_u451_o;
  wire _al_u452_o;
  wire _al_u454_o;
  wire _al_u455_o;
  wire _al_u456_o;
  wire _al_u457_o;
  wire _al_u459_o;
  wire _al_u461_o;
  wire _al_u462_o;
  wire _al_u464_o;
  wire _al_u465_o;
  wire _al_u467_o;
  wire _al_u468_o;
  wire _al_u469_o;
  wire _al_u470_o;
  wire _al_u471_o;
  wire _al_u472_o;
  wire _al_u475_o;
  wire _al_u476_o;
  wire _al_u478_o;
  wire _al_u479_o;
  wire _al_u481_o;
  wire _al_u482_o;
  wire _al_u485_o;
  wire _al_u486_o;
  wire _al_u487_o;
  wire _al_u489_o;
  wire _al_u490_o;
  wire _al_u493_o;
  wire _al_u494_o;
  wire _al_u496_o;
  wire _al_u497_o;
  wire _al_u499_o;
  wire _al_u500_o;
  wire _al_u501_o;
  wire _al_u502_o;
  wire _al_u505_o;
  wire _al_u507_o;
  wire _al_u508_o;
  wire _al_u510_o;
  wire _al_u511_o;
  wire _al_u512_o;
  wire _al_u514_o;
  wire _al_u515_o;
  wire _al_u516_o;
  wire _al_u517_o;
  wire _al_u519_o;
  wire _al_u520_o;
  wire _al_u521_o;
  wire _al_u522_o;
  wire _al_u523_o;
  wire _al_u524_o;
  wire _al_u526_o;
  wire _al_u527_o;
  wire _al_u528_o;
  wire _al_u529_o;
  wire _al_u530_o;
  wire _al_u531_o;
  wire _al_u533_o;
  wire _al_u534_o;
  wire _al_u535_o;
  wire _al_u536_o;
  wire _al_u537_o;
  wire _al_u538_o;
  wire _al_u540_o;
  wire _al_u541_o;
  wire _al_u542_o;
  wire _al_u543_o;
  wire _al_u544_o;
  wire _al_u545_o;
  wire _al_u546_o;
  wire _al_u547_o;
  wire _al_u548_o;
  wire _al_u549_o;
  wire _al_u550_o;
  wire _al_u551_o;
  wire _al_u553_o;
  wire _al_u554_o;
  wire _al_u555_o;
  wire _al_u556_o;
  wire _al_u557_o;
  wire _al_u558_o;
  wire _al_u559_o;
  wire _al_u560_o;
  wire _al_u562_o;
  wire _al_u563_o;
  wire _al_u564_o;
  wire _al_u565_o;
  wire _al_u566_o;
  wire _al_u567_o;
  wire _al_u568_o;
  wire _al_u569_o;
  wire _al_u570_o;
  wire _al_u571_o;
  wire _al_u572_o;
  wire _al_u573_o;
  wire _al_u575_o;
  wire _al_u576_o;
  wire _al_u577_o;
  wire _al_u578_o;
  wire _al_u579_o;
  wire _al_u580_o;
  wire _al_u581_o;
  wire _al_u582_o;
  wire _al_u583_o;
  wire _al_u584_o;
  wire _al_u585_o;
  wire _al_u586_o;
  wire _al_u587_o;
  wire _al_u588_o;
  wire _al_u589_o;
  wire _al_u590_o;
  wire _al_u592_o;
  wire _al_u593_o;
  wire _al_u594_o;
  wire _al_u595_o;
  wire _al_u596_o;
  wire _al_u597_o;
  wire _al_u599_o;
  wire _al_u600_o;
  wire _al_u601_o;
  wire _al_u602_o;
  wire _al_u603_o;
  wire _al_u604_o;
  wire _al_u605_o;
  wire _al_u606_o;
  wire _al_u607_o;
  wire _al_u608_o;
  wire _al_u610_o;
  wire _al_u611_o;
  wire _al_u612_o;
  wire _al_u613_o;
  wire _al_u614_o;
  wire _al_u615_o;
  wire _al_u616_o;
  wire _al_u617_o;
  wire _al_u618_o;
  wire _al_u619_o;
  wire _al_u620_o;
  wire _al_u621_o;
  wire _al_u622_o;
  wire _al_u623_o;
  wire _al_u624_o;
  wire _al_u625_o;
  wire _al_u627_o;
  wire _al_u628_o;
  wire _al_u629_o;
  wire _al_u630_o;
  wire _al_u631_o;
  wire _al_u632_o;
  wire _al_u633_o;
  wire _al_u634_o;
  wire _al_u636_o;
  wire _al_u637_o;
  wire _al_u638_o;
  wire _al_u639_o;
  wire _al_u640_o;
  wire _al_u641_o;
  wire _al_u642_o;
  wire _al_u643_o;
  wire _al_u644_o;
  wire _al_u645_o;
  wire _al_u646_o;
  wire _al_u647_o;
  wire _al_u648_o;
  wire _al_u649_o;
  wire _al_u64_o;
  wire _al_u651_o;
  wire _al_u652_o;
  wire _al_u653_o;
  wire _al_u654_o;
  wire _al_u655_o;
  wire _al_u656_o;
  wire _al_u657_o;
  wire _al_u658_o;
  wire _al_u659_o;
  wire _al_u65_o;
  wire _al_u660_o;
  wire _al_u661_o;
  wire _al_u662_o;
  wire _al_u663_o;
  wire _al_u664_o;
  wire _al_u665_o;
  wire _al_u666_o;
  wire _al_u667_o;
  wire _al_u668_o;
  wire _al_u66_o;
  wire _al_u670_o;
  wire _al_u671_o;
  wire _al_u672_o;
  wire _al_u673_o;
  wire _al_u674_o;
  wire _al_u675_o;
  wire _al_u676_o;
  wire _al_u677_o;
  wire _al_u678_o;
  wire _al_u679_o;
  wire _al_u67_o;
  wire _al_u680_o;
  wire _al_u681_o;
  wire _al_u682_o;
  wire _al_u683_o;
  wire _al_u685_o;
  wire _al_u686_o;
  wire _al_u687_o;
  wire _al_u688_o;
  wire _al_u689_o;
  wire _al_u690_o;
  wire _al_u691_o;
  wire _al_u692_o;
  wire _al_u693_o;
  wire _al_u694_o;
  wire _al_u695_o;
  wire _al_u696_o;
  wire _al_u697_o;
  wire _al_u698_o;
  wire _al_u699_o;
  wire _al_u700_o;
  wire _al_u702_o;
  wire _al_u703_o;
  wire _al_u704_o;
  wire _al_u705_o;
  wire _al_u706_o;
  wire _al_u707_o;
  wire _al_u708_o;
  wire _al_u709_o;
  wire _al_u70_o;
  wire _al_u710_o;
  wire _al_u711_o;
  wire _al_u712_o;
  wire _al_u713_o;
  wire _al_u714_o;
  wire _al_u716_o;
  wire _al_u717_o;
  wire _al_u718_o;
  wire _al_u719_o;
  wire _al_u71_o;
  wire _al_u720_o;
  wire _al_u721_o;
  wire _al_u722_o;
  wire _al_u723_o;
  wire _al_u724_o;
  wire _al_u725_o;
  wire _al_u726_o;
  wire _al_u727_o;
  wire _al_u728_o;
  wire _al_u729_o;
  wire _al_u730_o;
  wire _al_u731_o;
  wire _al_u732_o;
  wire _al_u733_o;
  wire _al_u735_o;
  wire _al_u736_o;
  wire _al_u737_o;
  wire _al_u738_o;
  wire _al_u739_o;
  wire _al_u740_o;
  wire _al_u741_o;
  wire _al_u742_o;
  wire _al_u743_o;
  wire _al_u744_o;
  wire _al_u745_o;
  wire _al_u746_o;
  wire _al_u747_o;
  wire _al_u748_o;
  wire _al_u749_o;
  wire _al_u750_o;
  wire _al_u751_o;
  wire _al_u753_o;
  wire _al_u754_o;
  wire _al_u755_o;
  wire _al_u756_o;
  wire _al_u757_o;
  wire _al_u758_o;
  wire _al_u759_o;
  wire _al_u75_o;
  wire _al_u760_o;
  wire _al_u761_o;
  wire _al_u762_o;
  wire _al_u763_o;
  wire _al_u764_o;
  wire _al_u765_o;
  wire _al_u766_o;
  wire _al_u767_o;
  wire _al_u768_o;
  wire _al_u769_o;
  wire _al_u770_o;
  wire _al_u771_o;
  wire _al_u773_o;
  wire _al_u774_o;
  wire _al_u775_o;
  wire _al_u776_o;
  wire _al_u777_o;
  wire _al_u778_o;
  wire _al_u779_o;
  wire _al_u780_o;
  wire _al_u781_o;
  wire _al_u784_o;
  wire _al_u785_o;
  wire _al_u786_o;
  wire _al_u787_o;
  wire _al_u788_o;
  wire _al_u789_o;
  wire _al_u78_o;
  wire _al_u790_o;
  wire _al_u791_o;
  wire _al_u792_o;
  wire _al_u793_o;
  wire _al_u795_o;
  wire _al_u797_o;
  wire _al_u798_o;
  wire _al_u799_o;
  wire _al_u79_o;
  wire _al_u800_o;
  wire _al_u801_o;
  wire _al_u802_o;
  wire _al_u804_o;
  wire _al_u805_o;
  wire _al_u806_o;
  wire _al_u808_o;
  wire _al_u809_o;
  wire _al_u810_o;
  wire _al_u811_o;
  wire _al_u812_o;
  wire _al_u813_o;
  wire _al_u814_o;
  wire _al_u815_o;
  wire _al_u816_o;
  wire _al_u817_o;
  wire _al_u818_o;
  wire _al_u820_o;
  wire _al_u821_o;
  wire _al_u823_o;
  wire _al_u824_o;
  wire _al_u825_o;
  wire _al_u826_o;
  wire _al_u827_o;
  wire _al_u829_o;
  wire _al_u830_o;
  wire _al_u832_o;
  wire _al_u833_o;
  wire _al_u834_o;
  wire _al_u835_o;
  wire _al_u837_o;
  wire _al_u839_o;
  wire _al_u840_o;
  wire _al_u842_o;
  wire _al_u843_o;
  wire _al_u844_o;
  wire _al_u845_o;
  wire _al_u86_o;
  wire _al_u87_o;
  wire _al_u92_o;
  wire _al_u93_o;
  wire _al_u96_o;
  wire _al_u98_o;
  wire _al_u99_o;
  wire \exp_diff[4]_neg_lutinv ;
  wire n100_lutinv;
  wire n101_lutinv;
  wire n102_lutinv;
  wire n103_lutinv;
  wire n104_lutinv;
  wire n105_lutinv;
  wire n106_lutinv;
  wire n107_lutinv;
  wire n112_lutinv;
  wire n165_lutinv;
  wire n198_lutinv;
  wire n221_lutinv;
  wire n222_lutinv;
  wire n223_lutinv;
  wire n224_lutinv;
  wire n225_lutinv;
  wire n226_lutinv;
  wire n227_lutinv;
  wire n228_lutinv;
  wire n229_lutinv;
  wire n230_lutinv;
  wire n231_lutinv;
  wire n232_lutinv;
  wire n233_lutinv;
  wire n234_lutinv;
  wire n235_lutinv;
  wire n236_lutinv;
  wire n237_lutinv;
  wire n238_lutinv;
  wire n239_lutinv;
  wire n5_lutinv;
  wire n63_lutinv;
  wire n86_lutinv;
  wire n87_lutinv;
  wire n88_lutinv;
  wire n89_lutinv;
  wire n90_lutinv;
  wire n91_lutinv;
  wire n92_lutinv;
  wire n93_lutinv;
  wire n94_lutinv;
  wire n95_lutinv;
  wire n96_lutinv;
  wire n97_lutinv;
  wire n98_lutinv;
  wire n99_lutinv;
  wire u194_sel_is_0_o;

  assign result[23] = \ADD03/ADD01/p0_neg ;
  EG_PHY_LSLICE #(
    //.MACRO("NM/add0/ucin_al_u848"),
    //.R_POSITION("X0Y1Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \NM/add0/u11_al_u851  (
    .a({M_result2[14],M_result2[12]}),
    .b({M_result2[15],M_result2[13]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\NM/add0/c11 ),
    .f({\NM/n4 [13],\NM/n4 [11]}),
    .fco(\NM/add0/c15 ),
    .fx({\NM/n4 [14],\NM/n4 [12]}));
  EG_PHY_LSLICE #(
    //.MACRO("NM/add0/ucin_al_u848"),
    //.R_POSITION("X0Y2Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \NM/add0/u15_al_u852  (
    .a({M_result2[18],M_result2[16]}),
    .b({M_result2[19],M_result2[17]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\NM/add0/c15 ),
    .f({\NM/n4 [17],\NM/n4 [15]}),
    .fco(\NM/add0/c19 ),
    .fx({\NM/n4 [18],\NM/n4 [16]}));
  EG_PHY_LSLICE #(
    //.MACRO("NM/add0/ucin_al_u848"),
    //.R_POSITION("X0Y2Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \NM/add0/u19_al_u853  (
    .a({M_result2[22],M_result2[20]}),
    .b({M_result2[23],M_result2[21]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\NM/add0/c19 ),
    .f({\NM/n4 [21],\NM/n4 [19]}),
    .fx({\NM/n4 [22],\NM/n4 [20]}));
  EG_PHY_LSLICE #(
    //.MACRO("NM/add0/ucin_al_u848"),
    //.R_POSITION("X0Y0Z1"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \NM/add0/u3_al_u849  (
    .a({M_result2[6],M_result2[4]}),
    .b({M_result2[7],M_result2[5]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\NM/add0/c3 ),
    .f({\NM/n4 [5],\NM/n4 [3]}),
    .fco(\NM/add0/c7 ),
    .fx({\NM/n4 [6],\NM/n4 [4]}));
  EG_PHY_LSLICE #(
    //.MACRO("NM/add0/ucin_al_u848"),
    //.R_POSITION("X0Y1Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'hA55A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \NM/add0/u7_al_u850  (
    .a({M_result2[10],M_result2[8]}),
    .b({M_result2[11],M_result2[9]}),
    .c(2'b00),
    .d(2'b00),
    .e(2'b00),
    .fci(\NM/add0/c7 ),
    .f({\NM/n4 [9],\NM/n4 [7]}),
    .fco(\NM/add0/c11 ),
    .fx({\NM/n4 [10],\NM/n4 [8]}));
  EG_PHY_LSLICE #(
    //.MACRO("NM/add0/ucin_al_u848"),
    //.R_POSITION("X0Y0Z0"),
    .DEMUX0("E"),
    .DEMUX1("E"),
    .INIT_LUTF0(16'h000A),
    .INIT_LUTF1(16'hA55A),
    .INIT_LUTG0(16'hC33C),
    .INIT_LUTG1(16'hC33C),
    .LSFMUX0("SUM"),
    .LSFMUX1("SUM"),
    .LSFXMUX0("SUM"),
    .LSFXMUX1("SUM"),
    .MODE("RIPPLE"))
    \NM/add0/ucin_al_u848  (
    .a({M_result2[2],1'b0}),
    .b({M_result2[3],M_result2[1]}),
    .c(2'b00),
    .d(2'b01),
    .e({1'b0,M_result[0]}),
    .f({\NM/n4 [1],open_n108}),
    .fco(\NM/add0/c3 ),
    .fx({\NM/n4 [2],\NM/n4 [0]}));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u100 (
    .a(_al_u67_o),
    .b(n1[11]),
    .c(n1[10]),
    .o(n99_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u101 (
    .a(_al_u67_o),
    .b(n1[9]),
    .c(n1[8]),
    .o(n101_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u102 (
    .a(n99_lutinv),
    .b(n101_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u102_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hdc7e))
    _al_u103 (
    .a(_al_u78_o),
    .b(_al_u79_o),
    .c(\C023/outtemp [3]),
    .d(\ADD01/ADD01/n3 ),
    .o(_al_u103_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(~C*B))"),
    .INIT(8'ha2))
    _al_u104 (
    .a(\exp_diff[4]_neg_lutinv ),
    .b(_al_u102_o),
    .c(_al_u103_o),
    .o(_al_u104_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*A))"),
    .INIT(8'hc4))
    _al_u105 (
    .a(_al_u79_o),
    .b(\C023/outtemp [3]),
    .c(\ADD01/ADD01/n3 ),
    .o(_al_u105_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u106 (
    .a(_al_u67_o),
    .b(n1[15]),
    .c(n1[14]),
    .o(n95_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u107 (
    .a(_al_u67_o),
    .b(n1[13]),
    .c(n1[12]),
    .o(n97_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u108 (
    .a(n95_lutinv),
    .b(n97_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u108_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u109 (
    .a(_al_u105_o),
    .b(_al_u108_o),
    .o(_al_u109_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C)"),
    .INIT(8'hb2))
    _al_u110 (
    .a(_al_u86_o),
    .b(n1[29]),
    .c(n2[29]),
    .o(_al_u110_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u111 (
    .a(\ADD01/ADD02/p1_lutinv ),
    .b(\ADD01/ADD02/p0_lutinv ),
    .o(\ADD01/ADD02/n3 ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h43f4c33c))
    _al_u112 (
    .a(\ADD01/ctemp_lutinv ),
    .b(_al_u110_o),
    .c(n1[30]),
    .d(n2[30]),
    .e(\ADD01/ADD02/n3 ),
    .o(_al_u112_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u113 (
    .a(\ADD01/ADD01/n20 ),
    .b(n1[27]),
    .c(n2[27]),
    .o(\C023/ADD01/ADD02/n0 ));
  AL_MAP_LUT4 #(
    .EQN("(B@(A*~(C)*~(D)+~(A)*C*~(D)+A*C*~(D)+A*C*D))"),
    .INIT(16'h6c36))
    _al_u114 (
    .a(\ADD01/ctemp_lutinv ),
    .b(\ADD01/ADD02/p1_lutinv ),
    .c(n1[27]),
    .d(n2[27]),
    .o(_al_u114_o));
  AL_MAP_LUT5 #(
    .EQN("(E@D@(C*~(B*A)))"),
    .INIT(32'h708f8f70))
    _al_u115 (
    .a(\ADD01/ctemp_lutinv ),
    .b(\ADD01/ADD02/n3 ),
    .c(_al_u86_o),
    .d(n1[29]),
    .e(n2[29]),
    .o(_al_u115_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*~B*A)"),
    .INIT(32'h20000000))
    _al_u116 (
    .a(_al_u112_o),
    .b(\C023/ADD01/ADD02/n0 ),
    .c(_al_u114_o),
    .d(_al_u78_o),
    .e(_al_u115_o),
    .o(_al_u116_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~A*~(~D*C*~B)))"),
    .INIT(32'haaba0000))
    _al_u117 (
    .a(_al_u93_o),
    .b(_al_u99_o),
    .c(_al_u104_o),
    .d(_al_u109_o),
    .e(_al_u116_o),
    .o(_al_u117_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u118 (
    .a(_al_u67_o),
    .b(n2[15]),
    .c(n2[14]),
    .o(n227_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u119 (
    .a(_al_u67_o),
    .b(n2[13]),
    .c(n2[12]),
    .o(n229_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u120 (
    .a(n227_lutinv),
    .b(n229_lutinv),
    .c(_al_u70_o),
    .o(_al_u120_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u121 (
    .a(_al_u67_o),
    .b(n2[11]),
    .c(n2[10]),
    .o(n231_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u122 (
    .a(_al_u67_o),
    .b(n2[9]),
    .c(n2[8]),
    .o(n233_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u123 (
    .a(n231_lutinv),
    .b(n233_lutinv),
    .c(_al_u70_o),
    .o(_al_u123_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u124 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u120_o),
    .d(_al_u123_o),
    .o(_al_u124_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u125 (
    .a(_al_u67_o),
    .b(n2[7]),
    .c(n2[6]),
    .o(n235_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u126 (
    .a(_al_u67_o),
    .b(n2[5]),
    .c(n2[4]),
    .o(n237_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u127 (
    .a(n235_lutinv),
    .b(n237_lutinv),
    .c(_al_u70_o),
    .o(_al_u127_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u128 (
    .a(_al_u67_o),
    .b(n2[3]),
    .c(n2[2]),
    .o(n239_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u129 (
    .a(_al_u67_o),
    .b(n2[1]),
    .c(n2[0]),
    .o(_al_u129_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'ha3))
    _al_u130 (
    .a(n239_lutinv),
    .b(_al_u129_o),
    .c(_al_u70_o),
    .o(_al_u130_o));
  AL_MAP_LUT4 #(
    .EQN("(D*(~C*~(B)*~(A)+~C*B*~(A)+~(~C)*B*A+~C*B*A))"),
    .INIT(16'h8d00))
    _al_u131 (
    .a(exp_diff[2]),
    .b(_al_u127_o),
    .c(_al_u130_o),
    .d(\C023/outtemp [3]),
    .o(_al_u131_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u132 (
    .a(_al_u67_o),
    .b(n2[22]),
    .o(_al_u132_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u133 (
    .a(_al_u67_o),
    .b(n2[21]),
    .c(n2[20]),
    .o(n221_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u134 (
    .a(_al_u132_o),
    .b(n221_lutinv),
    .c(_al_u70_o),
    .o(_al_u134_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u135 (
    .a(_al_u67_o),
    .b(n2[19]),
    .c(n2[18]),
    .o(n223_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u136 (
    .a(_al_u67_o),
    .b(n2[17]),
    .c(n2[16]),
    .o(n225_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u137 (
    .a(n223_lutinv),
    .b(n225_lutinv),
    .c(_al_u70_o),
    .o(_al_u137_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'h5c))
    _al_u138 (
    .a(_al_u134_o),
    .b(_al_u137_o),
    .c(_al_u79_o),
    .o(_al_u138_o));
  AL_MAP_LUT5 #(
    .EQN("~((~D*~C)*~((~B*~A))*~(E)+(~D*~C)*(~B*~A)*~(E)+~((~D*~C))*(~B*~A)*E+(~D*~C)*(~B*~A)*E)"),
    .INIT(32'heeeefff0))
    _al_u139 (
    .a(_al_u124_o),
    .b(_al_u131_o),
    .c(_al_u138_o),
    .d(exp_diff[3]),
    .e(\exp_diff[4]_neg_lutinv ),
    .o(_al_u139_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u140 (
    .a(_al_u112_o),
    .b(_al_u78_o),
    .c(_al_u115_o),
    .d(_al_u114_o),
    .o(_al_u140_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u141 (
    .a(_al_u78_o),
    .b(n1[0]),
    .o(_al_u141_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u142 (
    .a(_al_u78_o),
    .b(n2[0]),
    .o(_al_u142_o));
  AL_MAP_LUT5 #(
    .EQN("((~E*~(C*~B))@(~D*~A))"),
    .INIT(32'h0055cf9a))
    _al_u143 (
    .a(_al_u117_o),
    .b(_al_u139_o),
    .c(_al_u140_o),
    .d(_al_u141_o),
    .e(_al_u142_o),
    .o(M_result[0]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u144 (
    .a(_al_u117_o),
    .b(_al_u141_o),
    .o(_al_u144_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B*~A))"),
    .INIT(8'h0b))
    _al_u145 (
    .a(_al_u139_o),
    .b(_al_u140_o),
    .c(_al_u142_o),
    .o(_al_u145_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u146 (
    .a(_al_u67_o),
    .b(n1[14]),
    .c(n1[13]),
    .o(n96_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u147 (
    .a(_al_u67_o),
    .b(n1[16]),
    .c(n1[15]),
    .o(n94_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(A)*~((D@C))+B*A*~((D@C))+~(B)*A*(D@C)+B*A*(D@C))"),
    .INIT(16'h3553))
    _al_u148 (
    .a(n96_lutinv),
    .b(n94_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u148_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u149 (
    .a(_al_u67_o),
    .b(n1[4]),
    .c(n1[3]),
    .o(n106_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h717d))
    _al_u150 (
    .a(n106_lutinv),
    .b(_al_u70_o),
    .c(_al_u67_o),
    .d(n1[2]),
    .o(_al_u150_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hddfa))
    _al_u151 (
    .a(exp_diff[2]),
    .b(_al_u148_o),
    .c(_al_u150_o),
    .d(\C023/outtemp [3]),
    .o(_al_u151_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hb7bd))
    _al_u152 (
    .a(_al_u78_o),
    .b(_al_u79_o),
    .c(\C023/outtemp [3]),
    .d(\ADD01/ADD01/n3 ),
    .o(_al_u152_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u153 (
    .a(_al_u67_o),
    .b(n1[8]),
    .c(n1[7]),
    .o(n102_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u154 (
    .a(_al_u67_o),
    .b(n1[6]),
    .c(n1[5]),
    .o(n104_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u155 (
    .a(n102_lutinv),
    .b(n104_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u155_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u156 (
    .a(_al_u152_o),
    .b(_al_u155_o),
    .o(_al_u156_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u157 (
    .a(_al_u67_o),
    .b(n1[10]),
    .c(n1[9]),
    .o(n100_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u158 (
    .a(_al_u67_o),
    .b(n1[12]),
    .c(n1[11]),
    .o(n98_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(A)*~((D@C))+B*A*~((D@C))+~(B)*A*(D@C)+B*A*(D@C))"),
    .INIT(16'h3553))
    _al_u159 (
    .a(n100_lutinv),
    .b(n98_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u159_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*A*~(~E*~D))"),
    .INIT(32'h20202000))
    _al_u160 (
    .a(_al_u151_o),
    .b(_al_u156_o),
    .c(\exp_diff[4]_neg_lutinv ),
    .d(_al_u103_o),
    .e(_al_u159_o),
    .o(_al_u160_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u161 (
    .a(_al_u67_o),
    .b(n1[20]),
    .c(n1[19]),
    .o(n90_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u162 (
    .a(_al_u67_o),
    .b(n1[18]),
    .c(n1[17]),
    .o(n92_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u163 (
    .a(n90_lutinv),
    .b(n92_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u163_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(~E*~D*C*A))"),
    .INIT(32'hcccccc4c))
    _al_u164 (
    .a(_al_u64_o),
    .b(_al_u67_o),
    .c(_al_u65_o),
    .d(n1[30]),
    .e(n1[29]),
    .o(n86_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u165 (
    .a(_al_u67_o),
    .b(n1[22]),
    .c(n1[21]),
    .o(n88_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hace8))
    _al_u166 (
    .a(n86_lutinv),
    .b(n88_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u166_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A))"),
    .INIT(16'h2301))
    _al_u167 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u163_o),
    .d(_al_u166_o),
    .o(_al_u167_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u168 (
    .a(_al_u78_o),
    .b(n1[1]),
    .o(_al_u168_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*~A*~(~D*~B)))"),
    .INIT(32'h0000afbf))
    _al_u169 (
    .a(_al_u160_o),
    .b(_al_u167_o),
    .c(_al_u116_o),
    .d(\exp_diff[4]_neg_lutinv ),
    .e(_al_u168_o),
    .o(_al_u169_o));
  AL_MAP_LUT3 #(
    .EQN("~(B@(~C*A))"),
    .INIT(8'h39))
    _al_u170 (
    .a(_al_u78_o),
    .b(_al_u70_o),
    .c(_al_u67_o),
    .o(_al_u170_o));
  AL_MAP_LUT4 #(
    .EQN("(~(B)*~(C)*~((~D*A))+B*~(C)*~((~D*A))+B*C*~((~D*A))+~(B)*~(C)*(~D*A)+~(B)*C*(~D*A)+B*C*(~D*A))"),
    .INIT(16'hcfe7))
    _al_u171 (
    .a(_al_u78_o),
    .b(_al_u79_o),
    .c(\C023/outtemp [3]),
    .d(\ADD01/ADD01/n3 ),
    .o(_al_u171_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u172 (
    .a(_al_u67_o),
    .b(n2[4]),
    .c(n2[3]),
    .o(n238_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u173 (
    .a(_al_u67_o),
    .b(n2[2]),
    .c(n2[1]),
    .o(_al_u173_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A))"),
    .INIT(16'h1032))
    _al_u174 (
    .a(_al_u170_o),
    .b(_al_u171_o),
    .c(n238_lutinv),
    .d(_al_u173_o),
    .o(_al_u174_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u175 (
    .a(_al_u67_o),
    .b(n2[8]),
    .c(n2[7]),
    .o(n234_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u176 (
    .a(_al_u67_o),
    .b(n2[6]),
    .c(n2[5]),
    .o(n236_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u177 (
    .a(n234_lutinv),
    .b(n236_lutinv),
    .c(_al_u70_o),
    .o(_al_u177_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~A*~(~D*~B))"),
    .INIT(16'h5040))
    _al_u178 (
    .a(_al_u174_o),
    .b(_al_u152_o),
    .c(\exp_diff[4]_neg_lutinv ),
    .d(_al_u177_o),
    .o(_al_u178_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u179 (
    .a(_al_u67_o),
    .b(n2[22]),
    .c(n2[21]),
    .o(n165_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C)*~(B)+A*C*~(B)+~(A)*C*B+A*C*B)"),
    .INIT(8'he2))
    _al_u180 (
    .a(n165_lutinv),
    .b(_al_u70_o),
    .c(_al_u67_o),
    .o(_al_u180_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u181 (
    .a(_al_u67_o),
    .b(n2[20]),
    .c(n2[19]),
    .o(n222_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u182 (
    .a(_al_u67_o),
    .b(n2[18]),
    .c(n2[17]),
    .o(n224_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u183 (
    .a(n222_lutinv),
    .b(n224_lutinv),
    .c(_al_u70_o),
    .o(_al_u183_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(~B*(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)))"),
    .INIT(32'h0d0f0c0e))
    _al_u184 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(\exp_diff[4]_neg_lutinv ),
    .d(_al_u180_o),
    .e(_al_u183_o),
    .o(_al_u184_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u185 (
    .a(_al_u67_o),
    .b(n2[10]),
    .c(n2[9]),
    .o(n232_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u186 (
    .a(_al_u67_o),
    .b(n2[12]),
    .c(n2[11]),
    .o(n230_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u187 (
    .a(n232_lutinv),
    .b(n230_lutinv),
    .c(_al_u70_o),
    .o(_al_u187_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u188 (
    .a(_al_u67_o),
    .b(n2[14]),
    .c(n2[13]),
    .o(n228_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u189 (
    .a(_al_u67_o),
    .b(n2[16]),
    .c(n2[15]),
    .o(n226_lutinv));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u190 (
    .a(n228_lutinv),
    .b(n226_lutinv),
    .c(_al_u70_o),
    .o(_al_u190_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h048c))
    _al_u191 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u187_o),
    .d(_al_u190_o),
    .o(_al_u191_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u192 (
    .a(_al_u78_o),
    .b(n2[1]),
    .o(_al_u192_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*~B*~(~C*A)))"),
    .INIT(32'h0000ceff))
    _al_u193 (
    .a(_al_u178_o),
    .b(_al_u184_o),
    .c(_al_u191_o),
    .d(_al_u140_o),
    .e(_al_u192_o),
    .o(_al_u193_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u194 (
    .a(n1[31]),
    .b(n2[31]),
    .o(\M04/M01/M01/invSL_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*C*D*~(E)+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfee020f2))
    _al_u195 (
    .a(_al_u144_o),
    .b(_al_u145_o),
    .c(_al_u169_o),
    .d(_al_u193_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u195_o));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u196 (
    .a(n230_lutinv),
    .b(n228_lutinv),
    .c(_al_u70_o),
    .o(_al_u196_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u197 (
    .a(n224_lutinv),
    .b(n226_lutinv),
    .c(_al_u70_o),
    .o(_al_u197_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u198 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u196_o),
    .d(_al_u197_o),
    .o(_al_u198_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u199 (
    .a(n232_lutinv),
    .b(n234_lutinv),
    .c(_al_u70_o),
    .o(_al_u199_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C*~A))"),
    .INIT(8'h8c))
    _al_u200 (
    .a(_al_u152_o),
    .b(\exp_diff[4]_neg_lutinv ),
    .c(_al_u199_o),
    .o(_al_u200_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'hac))
    _al_u201 (
    .a(n236_lutinv),
    .b(n238_lutinv),
    .c(_al_u70_o),
    .o(_al_u201_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*~C))"),
    .INIT(16'h4440))
    _al_u202 (
    .a(_al_u198_o),
    .b(_al_u200_o),
    .c(_al_u171_o),
    .d(_al_u201_o),
    .o(_al_u202_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u203 (
    .a(n165_lutinv),
    .b(n222_lutinv),
    .c(_al_u70_o),
    .o(_al_u203_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u204 (
    .a(n86_lutinv),
    .b(_al_u70_o),
    .o(n112_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~C*~(D)*~(A)+~C*D*~(A)+~(~C)*D*A+~C*D*A))"),
    .INIT(16'h2301))
    _al_u205 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u203_o),
    .d(n112_lutinv),
    .o(_al_u205_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u206 (
    .a(_al_u205_o),
    .b(\exp_diff[4]_neg_lutinv ),
    .o(_al_u206_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u207 (
    .a(_al_u78_o),
    .b(n2[3]),
    .o(_al_u207_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~(C*~(~B*~A))))"),
    .INIT(32'hffe0001f))
    _al_u208 (
    .a(_al_u202_o),
    .b(_al_u206_o),
    .c(_al_u140_o),
    .d(_al_u207_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(new_M2[3]));
  AL_MAP_LUT3 #(
    .EQN("~(A*~(B)*~(C)+A*B*~(C)+~(A)*B*C+A*B*C)"),
    .INIT(8'h35))
    _al_u209 (
    .a(n227_lutinv),
    .b(n225_lutinv),
    .c(_al_u70_o),
    .o(_al_u209_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u210 (
    .a(n229_lutinv),
    .b(n231_lutinv),
    .c(_al_u70_o),
    .o(_al_u210_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))"),
    .INIT(16'h00d8))
    _al_u211 (
    .a(exp_diff[2]),
    .b(_al_u209_o),
    .c(_al_u210_o),
    .d(\C023/outtemp [3]),
    .o(_al_u211_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u212 (
    .a(_al_u170_o),
    .b(_al_u171_o),
    .c(n239_lutinv),
    .d(n237_lutinv),
    .o(_al_u212_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u213 (
    .a(n233_lutinv),
    .b(n235_lutinv),
    .c(_al_u70_o),
    .o(_al_u213_o));
  AL_MAP_LUT5 #(
    .EQN("(D*~B*~A*~(E*~C))"),
    .INIT(32'h10001100))
    _al_u214 (
    .a(_al_u211_o),
    .b(_al_u212_o),
    .c(_al_u152_o),
    .d(\exp_diff[4]_neg_lutinv ),
    .e(_al_u213_o),
    .o(_al_u214_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u215 (
    .a(_al_u132_o),
    .b(_al_u70_o),
    .o(_al_u215_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(A)*~(C)+B*A*~(C)+~(B)*A*C+B*A*C)"),
    .INIT(8'h53))
    _al_u216 (
    .a(n221_lutinv),
    .b(n223_lutinv),
    .c(_al_u70_o),
    .o(_al_u216_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~C*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B))"),
    .INIT(32'h0000080b))
    _al_u217 (
    .a(_al_u215_o),
    .b(exp_diff[2]),
    .c(exp_diff[3]),
    .d(_al_u216_o),
    .e(\exp_diff[4]_neg_lutinv ),
    .o(_al_u217_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u218 (
    .a(_al_u78_o),
    .b(n2[2]),
    .o(_al_u218_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~(C*~(~B*~A))))"),
    .INIT(32'hffe0001f))
    _al_u219 (
    .a(_al_u214_o),
    .b(_al_u217_o),
    .c(_al_u140_o),
    .d(_al_u218_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(new_M2[2]));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u220 (
    .a(n100_lutinv),
    .b(n102_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u220_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hafca))
    _al_u221 (
    .a(n104_lutinv),
    .b(n106_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u221_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~B*(~E*~(D)*~(A)+~E*D*~(A)+~(~E)*D*A+~E*D*A)))"),
    .INIT(32'hd0f0c0e0))
    _al_u222 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(\exp_diff[4]_neg_lutinv ),
    .d(_al_u220_o),
    .e(_al_u221_o),
    .o(_al_u222_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(A)*~((D@C))+B*A*~((D@C))+~(B)*A*(D@C)+B*A*(D@C))"),
    .INIT(16'h3553))
    _al_u223 (
    .a(n90_lutinv),
    .b(n88_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u223_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~B*(~D*~(E)*~(A)+~D*E*~(A)+~(~D)*E*A+~D*E*A))"),
    .INIT(32'h02030001))
    _al_u224 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(\exp_diff[4]_neg_lutinv ),
    .d(_al_u223_o),
    .e(n112_lutinv),
    .o(_al_u224_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u225 (
    .a(n96_lutinv),
    .b(n98_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u225_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u226 (
    .a(n92_lutinv),
    .b(n94_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u226_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u227 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u225_o),
    .d(_al_u226_o),
    .o(_al_u227_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u228 (
    .a(_al_u78_o),
    .b(n1[3]),
    .o(_al_u228_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*~(~B*~(~C*A))))"),
    .INIT(32'h000031ff))
    _al_u229 (
    .a(_al_u222_o),
    .b(_al_u224_o),
    .c(_al_u227_o),
    .d(_al_u116_o),
    .e(_al_u228_o),
    .o(_al_u229_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u230 (
    .a(_al_u170_o),
    .b(n87_lutinv),
    .o(n63_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(A)*~((D@C))+B*A*~((D@C))+~(B)*A*(D@C)+B*A*(D@C))"),
    .INIT(16'h3553))
    _al_u231 (
    .a(n91_lutinv),
    .b(n89_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u231_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(~E*~(A)*~(B)+~E*A*~(B)+~(~E)*A*B+~E*A*B))"),
    .INIT(32'h0008000b))
    _al_u232 (
    .a(n63_lutinv),
    .b(exp_diff[2]),
    .c(exp_diff[3]),
    .d(\exp_diff[4]_neg_lutinv ),
    .e(_al_u231_o),
    .o(_al_u232_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(A)*~((D@C))+B*A*~((D@C))+~(B)*A*(D@C)+B*A*(D@C))"),
    .INIT(16'h3553))
    _al_u233 (
    .a(n95_lutinv),
    .b(n93_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u233_o));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u234 (
    .a(n97_lutinv),
    .b(n99_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u234_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(B*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)))"),
    .INIT(32'h30b070f0))
    _al_u235 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(\exp_diff[4]_neg_lutinv ),
    .d(_al_u233_o),
    .e(_al_u234_o),
    .o(_al_u235_o));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(A)*~((D@C))+B*A*~((D@C))+~(B)*A*(D@C)+B*A*(D@C))"),
    .INIT(16'h3553))
    _al_u236 (
    .a(n103_lutinv),
    .b(n101_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u236_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h5135))
    _al_u237 (
    .a(n105_lutinv),
    .b(n107_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u237_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h3120))
    _al_u238 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u236_o),
    .d(_al_u237_o),
    .o(_al_u238_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u239 (
    .a(_al_u78_o),
    .b(n1[2]),
    .o(_al_u239_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*~(~A*~(~C*B))))"),
    .INIT(32'h000051ff))
    _al_u240 (
    .a(_al_u232_o),
    .b(_al_u235_o),
    .c(_al_u238_o),
    .d(_al_u116_o),
    .e(_al_u239_o),
    .o(_al_u240_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(C)*~((~D*B))+~(A)*C*~((~D*B))+A*C*~((~D*B))+~(A)*C*(~D*B))"),
    .INIT(16'hf571))
    _al_u241 (
    .a(new_M2[3]),
    .b(new_M2[2]),
    .c(_al_u229_o),
    .d(_al_u240_o),
    .o(_al_u241_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(~C*B)))"),
    .INIT(16'haa08))
    _al_u242 (
    .a(_al_u116_o),
    .b(_al_u71_o),
    .c(_al_u171_o),
    .d(\exp_diff[4]_neg_lutinv ),
    .o(_al_u242_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u243 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u108_o),
    .d(_al_u92_o),
    .o(_al_u243_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u244 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u96_o),
    .d(_al_u102_o),
    .o(_al_u244_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u245 (
    .a(_al_u78_o),
    .b(n1[4]),
    .o(_al_u245_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(A*~(D*~(~C*~B))))"),
    .INIT(32'h0000fd55))
    _al_u246 (
    .a(_al_u242_o),
    .b(_al_u243_o),
    .c(_al_u244_o),
    .d(\exp_diff[4]_neg_lutinv ),
    .e(_al_u245_o),
    .o(_al_u246_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~B*~(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)))"),
    .INIT(32'hf0d0e0c0))
    _al_u247 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(\exp_diff[4]_neg_lutinv ),
    .d(_al_u123_o),
    .e(_al_u127_o),
    .o(_al_u247_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(~C*B)))"),
    .INIT(16'haa08))
    _al_u248 (
    .a(_al_u140_o),
    .b(_al_u134_o),
    .c(_al_u171_o),
    .d(\exp_diff[4]_neg_lutinv ),
    .o(_al_u248_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A))"),
    .INIT(16'h0027))
    _al_u249 (
    .a(exp_diff[2]),
    .b(_al_u137_o),
    .c(_al_u120_o),
    .d(\C023/outtemp [3]),
    .o(_al_u249_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u250 (
    .a(_al_u78_o),
    .b(n2[4]),
    .o(_al_u250_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@(~D*~(B*~(~C*A))))"),
    .INIT(32'h003bffc4))
    _al_u251 (
    .a(_al_u247_o),
    .b(_al_u248_o),
    .c(_al_u249_o),
    .d(_al_u250_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u251_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u252 (
    .a(_al_u246_o),
    .b(_al_u251_o),
    .o(\ADD02/ADD01/ADD02/p0_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h3120))
    _al_u253 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u213_o),
    .d(_al_u212_o),
    .o(_al_u253_o));
  AL_MAP_LUT5 #(
    .EQN("(D*~(~A*~(E*~C*~B)))"),
    .INIT(32'hab00aa00))
    _al_u254 (
    .a(_al_u217_o),
    .b(_al_u253_o),
    .c(_al_u211_o),
    .d(_al_u140_o),
    .e(\exp_diff[4]_neg_lutinv ),
    .o(_al_u254_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@A@(~B*~(E*C)))"),
    .INIT(32'ha9569966))
    _al_u255 (
    .a(_al_u240_o),
    .b(_al_u254_o),
    .c(_al_u78_o),
    .d(\M04/M01/M01/invSL_lutinv ),
    .e(n2[2]),
    .o(_al_u255_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u256 (
    .a(_al_u229_o),
    .b(new_M2[3]),
    .o(\ADD02/ADD01/ADD01/p3_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(C*~(B*~(E*D*~A)))"),
    .INIT(32'h70303030))
    _al_u257 (
    .a(_al_u195_o),
    .b(_al_u241_o),
    .c(\ADD02/ADD01/ADD02/p0_lutinv ),
    .d(_al_u255_o),
    .e(\ADD02/ADD01/ADD01/p3_lutinv ),
    .o(_al_u257_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~B*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)))"),
    .INIT(32'hc0e0d0f0))
    _al_u258 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(\exp_diff[4]_neg_lutinv ),
    .d(_al_u196_o),
    .e(_al_u199_o),
    .o(_al_u258_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u259 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u203_o),
    .d(_al_u197_o),
    .o(_al_u259_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u260 (
    .a(n112_lutinv),
    .b(_al_u79_o),
    .o(n198_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u261 (
    .a(n198_lutinv),
    .b(exp_diff[3]),
    .c(\exp_diff[4]_neg_lutinv ),
    .o(_al_u261_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u262 (
    .a(_al_u78_o),
    .b(n2[7]),
    .o(_al_u262_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*~(~C*~(~B*A))))"),
    .INIT(32'h00000dff))
    _al_u263 (
    .a(_al_u258_o),
    .b(_al_u259_o),
    .c(_al_u261_o),
    .d(_al_u140_o),
    .e(_al_u262_o),
    .o(_al_u263_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~B*(E*~(D)*~(A)+E*D*~(A)+~(E)*D*A+E*D*A)))"),
    .INIT(32'hc0e0d0f0))
    _al_u264 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(\exp_diff[4]_neg_lutinv ),
    .d(_al_u225_o),
    .e(_al_u220_o),
    .o(_al_u264_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'hc480))
    _al_u265 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u223_o),
    .d(_al_u226_o),
    .o(_al_u265_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u266 (
    .a(_al_u78_o),
    .b(n1[7]),
    .o(_al_u266_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*~(~C*~(~B*A))))"),
    .INIT(32'h00000dff))
    _al_u267 (
    .a(_al_u264_o),
    .b(_al_u265_o),
    .c(_al_u261_o),
    .d(_al_u116_o),
    .e(_al_u266_o),
    .o(_al_u267_o));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u268 (
    .a(_al_u263_o),
    .b(_al_u267_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u268_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(~C*B)))"),
    .INIT(16'haa08))
    _al_u269 (
    .a(_al_u116_o),
    .b(_al_u166_o),
    .c(_al_u171_o),
    .d(\exp_diff[4]_neg_lutinv ),
    .o(_al_u269_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u270 (
    .a(_al_u78_o),
    .b(n1[5]),
    .o(_al_u270_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*C*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hf0ca))
    _al_u271 (
    .a(_al_u155_o),
    .b(_al_u159_o),
    .c(exp_diff[2]),
    .d(exp_diff[3]),
    .o(_al_u271_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*~(B)*~(C)*~(D)+~(A)*B*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h530f))
    _al_u272 (
    .a(_al_u163_o),
    .b(_al_u148_o),
    .c(_al_u271_o),
    .d(exp_diff[3]),
    .o(_al_u272_o));
  AL_MAP_LUT4 #(
    .EQN("~(~C*~((~D*B))*~(A)+~C*(~D*B)*~(A)+~(~C)*(~D*B)*A+~C*(~D*B)*A)"),
    .INIT(16'hfa72))
    _al_u273 (
    .a(_al_u269_o),
    .b(\exp_diff[4]_neg_lutinv ),
    .c(_al_u270_o),
    .d(_al_u272_o),
    .o(M1[5]));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h084c))
    _al_u274 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u183_o),
    .d(_al_u190_o),
    .o(_al_u274_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~C*~(D*~B)))"),
    .INIT(16'ha2a0))
    _al_u275 (
    .a(_al_u140_o),
    .b(_al_u171_o),
    .c(\exp_diff[4]_neg_lutinv ),
    .d(_al_u180_o),
    .o(_al_u275_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u276 (
    .a(_al_u171_o),
    .b(\exp_diff[4]_neg_lutinv ),
    .c(_al_u177_o),
    .o(_al_u276_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u277 (
    .a(_al_u152_o),
    .b(_al_u187_o),
    .o(_al_u277_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u278 (
    .a(_al_u78_o),
    .b(n2[5]),
    .o(_al_u278_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(B*~(~D*C*~A)))"),
    .INIT(32'h00003373))
    _al_u279 (
    .a(_al_u274_o),
    .b(_al_u275_o),
    .c(_al_u276_o),
    .d(_al_u277_o),
    .e(_al_u278_o),
    .o(_al_u279_o));
  AL_MAP_LUT3 #(
    .EQN("(A*(C@B))"),
    .INIT(8'h28))
    _al_u280 (
    .a(M1[5]),
    .b(_al_u279_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD01/ADD02/g1 ));
  AL_MAP_LUT4 #(
    .EQN("(B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'hc840))
    _al_u281 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u233_o),
    .d(_al_u231_o),
    .o(_al_u281_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h3120))
    _al_u282 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u234_o),
    .d(_al_u236_o),
    .o(_al_u282_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u283 (
    .a(_al_u170_o),
    .b(_al_u171_o),
    .c(n87_lutinv),
    .o(n5_lutinv));
  AL_MAP_LUT5 #(
    .EQN("(D*(C*~((~B*~A))*~(E)+C*(~B*~A)*~(E)+~(C)*(~B*~A)*E+C*(~B*~A)*E))"),
    .INIT(32'h1100f000))
    _al_u284 (
    .a(_al_u281_o),
    .b(_al_u282_o),
    .c(n5_lutinv),
    .d(_al_u116_o),
    .e(\exp_diff[4]_neg_lutinv ),
    .o(_al_u284_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*~B))"),
    .INIT(8'h45))
    _al_u285 (
    .a(_al_u284_o),
    .b(_al_u78_o),
    .c(n1[6]),
    .o(_al_u285_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hf7b3d591))
    _al_u286 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u216_o),
    .d(_al_u209_o),
    .e(_al_u210_o),
    .o(_al_u286_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(~D*~(~C*B)))"),
    .INIT(16'haa08))
    _al_u287 (
    .a(_al_u140_o),
    .b(_al_u215_o),
    .c(_al_u171_o),
    .d(\exp_diff[4]_neg_lutinv ),
    .o(_al_u287_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u288 (
    .a(_al_u171_o),
    .b(_al_u213_o),
    .o(_al_u288_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u289 (
    .a(_al_u78_o),
    .b(n2[6]),
    .o(_al_u289_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(B*~(D*~C*A)))"),
    .INIT(32'h00003b33))
    _al_u290 (
    .a(_al_u286_o),
    .b(_al_u287_o),
    .c(_al_u288_o),
    .d(\exp_diff[4]_neg_lutinv ),
    .e(_al_u289_o),
    .o(_al_u290_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u291 (
    .a(_al_u290_o),
    .b(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u291_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(~(B)*~(C)*~(D)+B*~(C)*~(D)+B*C*~(D)+B*~(C)*D)*~(E)*~(A)+~(~(B)*~(C)*~(D)+B*~(C)*~(D)+B*C*~(D)+B*~(C)*D)*E*~(A)+~(~(~(B)*~(C)*~(D)+B*~(C)*~(D)+B*C*~(D)+B*~(C)*D))*E*A+~(~(B)*~(C)*~(D)+B*~(C)*~(D)+B*C*~(D)+B*~(C)*D)*E*A)"),
    .INIT(32'h0445aeef))
    _al_u292 (
    .a(_al_u268_o),
    .b(\ADD02/ADD01/ADD02/g1 ),
    .c(_al_u285_o),
    .d(_al_u291_o),
    .e(_al_u267_o),
    .o(_al_u292_o));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u293 (
    .a(M1[5]),
    .b(_al_u279_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD01/ADD02/p1_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(B*~A*~(E@D@C))"),
    .INIT(32'h04404004))
    _al_u294 (
    .a(_al_u268_o),
    .b(\ADD02/ADD01/ADD02/p1_lutinv ),
    .c(_al_u285_o),
    .d(_al_u290_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u294_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u295 (
    .a(_al_u246_o),
    .b(_al_u251_o),
    .o(\ADD02/ADD01/ADD02/g0 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(C*~(~D*~A)))"),
    .INIT(16'h0313))
    _al_u296 (
    .a(_al_u257_o),
    .b(_al_u292_o),
    .c(_al_u294_o),
    .d(\ADD02/ADD01/ADD02/g0 ),
    .o(_al_u296_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u297 (
    .a(_al_u116_o),
    .b(\exp_diff[4]_neg_lutinv ),
    .o(_al_u297_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*~(B)*C*D+~(A)*B*C*D)"),
    .INIT(16'h62ea))
    _al_u298 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u163_o),
    .d(_al_u166_o),
    .o(_al_u298_o));
  AL_MAP_LUT5 #(
    .EQN("(A*(~(B)*~(C)*~(D)*~(E)+B*~(C)*~(D)*~(E)+~(B)*C*~(D)*~(E)+~(B)*~(C)*D*~(E)+~(B)*C*D*~(E)+B*~(C)*~(D)*E+~(B)*C*~(D)*E+~(B)*C*D*E))"),
    .INIT(32'h2028222a))
    _al_u299 (
    .a(_al_u297_o),
    .b(_al_u298_o),
    .c(exp_diff[3]),
    .d(_al_u148_o),
    .e(_al_u159_o),
    .o(_al_u299_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u300 (
    .a(_al_u140_o),
    .b(\exp_diff[4]_neg_lutinv ),
    .o(_al_u300_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(B)*~(A)+~C*B*~(A)+~(~C)*B*A+~C*B*A)"),
    .INIT(8'h8d))
    _al_u301 (
    .a(exp_diff[2]),
    .b(_al_u180_o),
    .c(_al_u183_o),
    .o(_al_u301_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u302 (
    .a(exp_diff[2]),
    .b(_al_u187_o),
    .c(_al_u190_o),
    .o(_al_u302_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u303 (
    .a(_al_u78_o),
    .b(n2[9]),
    .o(_al_u303_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)))"),
    .INIT(32'h0000775f))
    _al_u304 (
    .a(_al_u300_o),
    .b(_al_u301_o),
    .c(_al_u302_o),
    .d(exp_diff[3]),
    .e(_al_u303_o),
    .o(_al_u304_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@B@(~A*~(E*~C)))"),
    .INIT(32'h9c639966))
    _al_u305 (
    .a(_al_u299_o),
    .b(_al_u304_o),
    .c(_al_u78_o),
    .d(\M04/M01/M01/invSL_lutinv ),
    .e(n1[9]),
    .o(\ADD02/ADD02/ADD01/p1_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h3120))
    _al_u306 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u120_o),
    .d(_al_u123_o),
    .o(_al_u306_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B))"),
    .INIT(16'h0074))
    _al_u307 (
    .a(_al_u134_o),
    .b(exp_diff[2]),
    .c(_al_u137_o),
    .d(\C023/outtemp [3]),
    .o(_al_u307_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u308 (
    .a(_al_u78_o),
    .b(n2[8]),
    .o(_al_u308_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~(~C*~B*A)))"),
    .INIT(32'hff0200fd))
    _al_u309 (
    .a(_al_u300_o),
    .b(_al_u306_o),
    .c(_al_u307_o),
    .d(_al_u308_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(new_M2[8]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u310 (
    .a(_al_u71_o),
    .b(exp_diff[2]),
    .c(_al_u92_o),
    .o(_al_u310_o));
  AL_MAP_LUT5 #(
    .EQN("~(~(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(A)*~(C)+~(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*A*~(C)+~(~(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*A*C+~(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*A*C)"),
    .INIT(32'h5f535c50))
    _al_u311 (
    .a(_al_u310_o),
    .b(exp_diff[2]),
    .c(exp_diff[3]),
    .d(_al_u108_o),
    .e(_al_u102_o),
    .o(_al_u311_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(~(E*~D)*~(C*~B)))"),
    .INIT(32'h20aa2020))
    _al_u312 (
    .a(new_M2[8]),
    .b(_al_u311_o),
    .c(_al_u297_o),
    .d(_al_u78_o),
    .e(n1[8]),
    .o(\ADD02/ADD02/ADD01/g0 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u313 (
    .a(\ADD02/ADD02/ADD01/p1_lutinv ),
    .b(\ADD02/ADD02/ADD01/g0 ),
    .o(\ADD02/ADD02/ADD01/n1 ));
  AL_MAP_LUT5 #(
    .EQN("((D@B)*~(~(E*~C)*~A))"),
    .INIT(32'h238c2288))
    _al_u314 (
    .a(_al_u299_o),
    .b(_al_u304_o),
    .c(_al_u78_o),
    .d(\M04/M01/M01/invSL_lutinv ),
    .e(n1[9]),
    .o(\ADD02/ADD02/ADD01/g1 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u315 (
    .a(\ADD02/ADD02/ADD01/n1 ),
    .b(\ADD02/ADD02/ADD01/g1 ),
    .o(_al_u315_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h7f737c70))
    _al_u316 (
    .a(n63_lutinv),
    .b(exp_diff[2]),
    .c(exp_diff[3]),
    .d(_al_u233_o),
    .e(_al_u234_o),
    .o(_al_u316_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u317 (
    .a(_al_u103_o),
    .b(_al_u231_o),
    .o(_al_u317_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*~D)*~(B*~(~C*A)))"),
    .INIT(32'h3b003b3b))
    _al_u318 (
    .a(_al_u316_o),
    .b(_al_u297_o),
    .c(_al_u317_o),
    .d(_al_u78_o),
    .e(n1[10]),
    .o(_al_u318_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~(A)*~(B)+~C*A*~(B)+~(~C)*A*B+~C*A*B)"),
    .INIT(8'h8b))
    _al_u319 (
    .a(_al_u215_o),
    .b(exp_diff[2]),
    .c(_al_u216_o),
    .o(_al_u319_o));
  AL_MAP_LUT3 #(
    .EQN("~(C*~(B)*~(A)+C*B*~(A)+~(C)*B*A+C*B*A)"),
    .INIT(8'h27))
    _al_u320 (
    .a(exp_diff[2]),
    .b(_al_u209_o),
    .c(_al_u210_o),
    .o(_al_u320_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u321 (
    .a(_al_u78_o),
    .b(n2[10]),
    .o(_al_u321_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(A*(C*~(B)*~(D)+C*B*~(D)+~(C)*B*D+C*B*D)))"),
    .INIT(32'h0000775f))
    _al_u322 (
    .a(_al_u300_o),
    .b(_al_u319_o),
    .c(_al_u320_o),
    .d(exp_diff[3]),
    .e(_al_u321_o),
    .o(_al_u322_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u323 (
    .a(_al_u318_o),
    .b(_al_u322_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u323_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u324 (
    .a(_al_u318_o),
    .b(_al_u322_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD02/ADD01/g2 ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u325 (
    .a(_al_u323_o),
    .b(\ADD02/ADD02/ADD01/g2 ),
    .o(\ADD02/ADD02/ADD01/p2_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("~(A@(~(E*~D)*~(C*~B)))"),
    .INIT(32'h9a559a9a))
    _al_u326 (
    .a(new_M2[8]),
    .b(_al_u311_o),
    .c(_al_u297_o),
    .d(_al_u78_o),
    .e(n1[8]),
    .o(\ADD02/ADD02/ADD01/p0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u327 (
    .a(\ADD02/ADD02/ADD01/p1_lutinv ),
    .b(\ADD02/ADD02/ADD01/p0_lutinv ),
    .o(\ADD02/ADD02/ADD01/n3 ));
  AL_MAP_LUT4 #(
    .EQN("~(C@(B*~(D*~A)))"),
    .INIT(16'h87c3))
    _al_u328 (
    .a(_al_u296_o),
    .b(_al_u315_o),
    .c(\ADD02/ADD02/ADD01/p2_lutinv ),
    .d(\ADD02/ADD02/ADD01/n3 ),
    .o(_al_u328_o));
  AL_MAP_LUT3 #(
    .EQN("~(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'h1b))
    _al_u329 (
    .a(exp_diff[2]),
    .b(_al_u225_o),
    .c(_al_u226_o),
    .o(_al_u329_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'h4e))
    _al_u330 (
    .a(exp_diff[2]),
    .b(_al_u223_o),
    .c(n112_lutinv),
    .o(_al_u330_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u331 (
    .a(_al_u78_o),
    .b(n1[11]),
    .o(_al_u331_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(A*~(~B*~(C)*~(D)+~B*C*~(D)+~(~B)*C*D+~B*C*D)))"),
    .INIT(32'h0000f577))
    _al_u332 (
    .a(_al_u297_o),
    .b(_al_u329_o),
    .c(_al_u330_o),
    .d(exp_diff[3]),
    .e(_al_u331_o),
    .o(_al_u332_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(C*~(D)*~(A)+C*D*~(A)+~(C)*D*A+C*D*A))"),
    .INIT(16'h3210))
    _al_u333 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u196_o),
    .d(_al_u197_o),
    .o(_al_u333_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'h4e))
    _al_u334 (
    .a(exp_diff[2]),
    .b(_al_u203_o),
    .c(n112_lutinv),
    .o(_al_u334_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u335 (
    .a(_al_u78_o),
    .b(n2[11]),
    .o(_al_u335_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(~B*A*~(~E*C)))"),
    .INIT(32'h00dd00fd))
    _al_u336 (
    .a(_al_u300_o),
    .b(_al_u333_o),
    .c(_al_u334_o),
    .d(_al_u335_o),
    .e(\C023/outtemp [3]),
    .o(_al_u336_o));
  AL_MAP_LUT3 #(
    .EQN("(C@B@A)"),
    .INIT(8'h96))
    _al_u337 (
    .a(_al_u332_o),
    .b(_al_u336_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u337_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u338 (
    .a(\ADD02/ADD02/ADD01/p1_lutinv ),
    .b(_al_u337_o),
    .o(_al_u338_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~((D@C))*~(E)+~(A)*B*~((D@C))*~(E)+~(A)*~(B)*(D@C)*~(E)+A*~(B)*(D@C)*~(E)+~(A)*B*(D@C)*~(E)+A*B*(D@C)*~(E)+~(A)*~(B)*~((D@C))*E+A*~(B)*~((D@C))*E+~(A)*B*~((D@C))*E+A*~(B)*(D@C)*E+~(A)*B*(D@C)*E+A*B*(D@C)*E)"),
    .INIT(32'h7ee76ff6))
    _al_u339 (
    .a(_al_u144_o),
    .b(_al_u145_o),
    .c(_al_u169_o),
    .d(_al_u193_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u339_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u340 (
    .a(new_M2[2]),
    .b(_al_u240_o),
    .o(\ADD02/ADD01/ADD01/g2 ));
  AL_MAP_LUT5 #(
    .EQN("(~B*(A*~(C)*~(D)*~(E)+A*C*~(D)*E+~(A)*~(C)*D*E+~(A)*C*D*E))"),
    .INIT(32'h11200002))
    _al_u341 (
    .a(_al_u195_o),
    .b(_al_u339_o),
    .c(\ADD02/ADD01/ADD01/g2 ),
    .d(_al_u255_o),
    .e(\ADD02/ADD01/ADD01/p3_lutinv ),
    .o(_al_u341_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~(B*~(C*~A))))"),
    .INIT(32'hff8c0073))
    _al_u342 (
    .a(_al_u272_o),
    .b(_al_u269_o),
    .c(\exp_diff[4]_neg_lutinv ),
    .d(_al_u270_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u342_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(D*~(~C*~B)))"),
    .INIT(16'h02aa))
    _al_u343 (
    .a(_al_u242_o),
    .b(_al_u243_o),
    .c(_al_u244_o),
    .d(\exp_diff[4]_neg_lutinv ),
    .o(_al_u343_o));
  AL_MAP_LUT5 #(
    .EQN("(((~E*~B)@D)*~(C@A))"),
    .INIT(32'ha5008421))
    _al_u344 (
    .a(_al_u342_o),
    .b(_al_u343_o),
    .c(_al_u279_o),
    .d(_al_u251_o),
    .e(_al_u245_o),
    .o(\ADD02/ADD01/ADD02/n3 ));
  AL_MAP_LUT5 #(
    .EQN("(C*~(B*~(E*D*~A)))"),
    .INIT(32'h70303030))
    _al_u345 (
    .a(_al_u195_o),
    .b(_al_u241_o),
    .c(\ADD02/ADD01/ADD02/n3 ),
    .d(_al_u255_o),
    .e(\ADD02/ADD01/ADD01/p3_lutinv ),
    .o(_al_u345_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u346 (
    .a(_al_u285_o),
    .b(_al_u291_o),
    .o(\ADD02/ADD01/ADD02/p2_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u347 (
    .a(_al_u341_o),
    .b(_al_u345_o),
    .c(\ADD02/ADD01/ADD02/p2_lutinv ),
    .o(_al_u347_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*~A))"),
    .INIT(16'h8ccc))
    _al_u348 (
    .a(_al_u195_o),
    .b(_al_u241_o),
    .c(_al_u255_o),
    .d(\ADD02/ADD01/ADD01/p3_lutinv ),
    .o(_al_u348_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~((~A*~(C*B)))*~(D)+E*(~A*~(C*B))*~(D)+~(E)*(~A*~(C*B))*D+E*(~A*~(C*B))*D)"),
    .INIT(32'h15ff1500))
    _al_u349 (
    .a(\ADD02/ADD01/ADD02/g1 ),
    .b(\ADD02/ADD01/ADD02/p1_lutinv ),
    .c(\ADD02/ADD01/ADD02/g0 ),
    .d(\ADD02/ADD01/ADD02/p2_lutinv ),
    .e(_al_u285_o),
    .o(_al_u349_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(B*~(D*C*~A)))"),
    .INIT(32'h73338ccc))
    _al_u350 (
    .a(_al_u348_o),
    .b(_al_u349_o),
    .c(\ADD02/ADD01/ADD02/p2_lutinv ),
    .d(\ADD02/ADD01/ADD02/n3 ),
    .e(_al_u268_o),
    .o(_al_u350_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@(~B*~(C*~(~D*~A))))"),
    .INIT(32'h0313fcec))
    _al_u351 (
    .a(_al_u257_o),
    .b(_al_u292_o),
    .c(_al_u294_o),
    .d(\ADD02/ADD01/ADD02/g0 ),
    .e(\ADD02/ADD02/ADD01/p0_lutinv ),
    .o(_al_u351_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*~A)"),
    .INIT(32'h00000040))
    _al_u352 (
    .a(_al_u328_o),
    .b(_al_u338_o),
    .c(_al_u347_o),
    .d(_al_u350_o),
    .e(_al_u351_o),
    .o(_al_u352_o));
  AL_MAP_LUT5 #(
    .EQN("((C@B)*~((D@A))*~(E)+~((C@B))*(D@A)*~(E)+(C@B)*(D@A)*~(E)+~((C@B))*~((D@A))*E+(C@B)*~((D@A))*E+~((C@B))*(D@A)*E)"),
    .INIT(32'hebd77dbe))
    _al_u353 (
    .a(_al_u318_o),
    .b(_al_u332_o),
    .c(_al_u336_o),
    .d(_al_u322_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u353_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u354 (
    .a(_al_u353_o),
    .b(\ADD02/ADD02/ADD01/p1_lutinv ),
    .c(\ADD02/ADD02/ADD01/p0_lutinv ),
    .o(_al_u354_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(~B*~(D*~(~E*~A))))"),
    .INIT(32'hf0c0e0c0))
    _al_u355 (
    .a(_al_u257_o),
    .b(_al_u292_o),
    .c(_al_u354_o),
    .d(_al_u294_o),
    .e(\ADD02/ADD01/ADD02/g0 ),
    .o(_al_u355_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hdfdcd3d0))
    _al_u356 (
    .a(_al_u71_o),
    .b(exp_diff[2]),
    .c(exp_diff[3]),
    .d(_al_u108_o),
    .e(_al_u92_o),
    .o(_al_u356_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(~C*~A))"),
    .INIT(8'hc8))
    _al_u357 (
    .a(_al_u140_o),
    .b(\exp_diff[4]_neg_lutinv ),
    .c(_al_u116_o),
    .o(u194_sel_is_0_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((B*~A))*~(C)+D*(B*~A)*~(C)+~(D)*(B*~A)*C+D*(B*~A)*C)"),
    .INIT(16'hb0bf))
    _al_u358 (
    .a(_al_u356_o),
    .b(u194_sel_is_0_o),
    .c(_al_u78_o),
    .d(n1[12]),
    .o(_al_u358_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hdfd3dcd0))
    _al_u359 (
    .a(_al_u134_o),
    .b(exp_diff[2]),
    .c(exp_diff[3]),
    .d(_al_u137_o),
    .e(_al_u120_o),
    .o(_al_u359_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*~A))"),
    .INIT(16'h0bbb))
    _al_u360 (
    .a(_al_u359_o),
    .b(_al_u300_o),
    .c(_al_u78_o),
    .d(n2[12]),
    .o(_al_u360_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@B@A)"),
    .INIT(8'h69))
    _al_u361 (
    .a(_al_u358_o),
    .b(_al_u360_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD02/ADD02/p0_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hdfdcd3d0))
    _al_u362 (
    .a(n63_lutinv),
    .b(exp_diff[2]),
    .c(exp_diff[3]),
    .d(_al_u233_o),
    .e(_al_u231_o),
    .o(_al_u362_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*~A))"),
    .INIT(16'hb0bb))
    _al_u363 (
    .a(_al_u362_o),
    .b(_al_u297_o),
    .c(_al_u78_o),
    .d(n1[14]),
    .o(_al_u363_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h0213))
    _al_u364 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u216_o),
    .d(_al_u209_o),
    .o(_al_u364_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(~C*B))"),
    .INIT(8'h51))
    _al_u365 (
    .a(_al_u364_o),
    .b(_al_u215_o),
    .c(_al_u103_o),
    .o(_al_u365_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u366 (
    .a(_al_u78_o),
    .b(n2[14]),
    .o(_al_u366_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@A@(~D*~(C*~B)))"),
    .INIT(32'haa65559a))
    _al_u367 (
    .a(_al_u363_o),
    .b(_al_u365_o),
    .c(_al_u300_o),
    .d(_al_u366_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD02/ADD02/p2_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hb9fda8ec))
    _al_u368 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u163_o),
    .d(_al_u166_o),
    .e(_al_u148_o),
    .o(_al_u368_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((B*~A))*~(C)+D*(B*~A)*~(C)+~(D)*(B*~A)*C+D*(B*~A)*C)"),
    .INIT(16'hb0bf))
    _al_u369 (
    .a(_al_u368_o),
    .b(u194_sel_is_0_o),
    .c(_al_u78_o),
    .d(n1[13]),
    .o(_al_u369_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*~(B)*C*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+A*B*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'hbf9dae8c))
    _al_u370 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u180_o),
    .d(_al_u183_o),
    .e(_al_u190_o),
    .o(_al_u370_o));
  AL_MAP_LUT4 #(
    .EQN("~((B*~A)*~(D)*~(C)+(B*~A)*D*~(C)+~((B*~A))*D*C+(B*~A)*D*C)"),
    .INIT(16'h0bfb))
    _al_u371 (
    .a(_al_u370_o),
    .b(u194_sel_is_0_o),
    .c(_al_u78_o),
    .d(n2[13]),
    .o(_al_u371_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@B@A)"),
    .INIT(8'h69))
    _al_u372 (
    .a(_al_u369_o),
    .b(_al_u371_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD02/ADD02/p1_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u373 (
    .a(\ADD02/ADD02/ADD02/p0_lutinv ),
    .b(\ADD02/ADD02/ADD02/p2_lutinv ),
    .c(\ADD02/ADD02/ADD02/p1_lutinv ),
    .o(\ADD02/ADD02/ADD02/n10 ));
  AL_MAP_LUT4 #(
    .EQN("(~B*(D*~(C)*~(A)+D*C*~(A)+~(D)*C*A+D*C*A))"),
    .INIT(16'h3120))
    _al_u374 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u203_o),
    .d(_al_u197_o),
    .o(_al_u374_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*~C))"),
    .INIT(16'h2022))
    _al_u375 (
    .a(_al_u300_o),
    .b(_al_u374_o),
    .c(n198_lutinv),
    .d(exp_diff[3]),
    .o(_al_u375_o));
  AL_MAP_LUT4 #(
    .EQN("(C@(~A*~(D*B)))"),
    .INIT(16'he1a5))
    _al_u376 (
    .a(_al_u375_o),
    .b(_al_u78_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .d(n2[15]),
    .o(new_M2[15]));
  AL_MAP_LUT5 #(
    .EQN("(~(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*~(A)*~(C)+~(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*A*~(C)+~(~(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B))*A*C+~(E*~(D)*~(B)+E*D*~(B)+~(E)*D*B+E*D*B)*A*C)"),
    .INIT(32'ha0aca3af))
    _al_u377 (
    .a(n198_lutinv),
    .b(exp_diff[2]),
    .c(exp_diff[3]),
    .d(_al_u223_o),
    .e(_al_u226_o),
    .o(_al_u377_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*A))"),
    .INIT(16'h7077))
    _al_u378 (
    .a(_al_u297_o),
    .b(_al_u377_o),
    .c(_al_u78_o),
    .d(n1[15]),
    .o(_al_u378_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u379 (
    .a(new_M2[15]),
    .b(_al_u378_o),
    .o(\ADD02/ADD02/ADD02/p3_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u380 (
    .a(\ADD02/ADD02/ADD02/n10 ),
    .b(\ADD02/ADD02/ADD02/p3_lutinv ),
    .o(_al_u380_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*B*C*D*~(E)+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E+A*B*C*D*E)"),
    .INIT(32'hfce88ecf))
    _al_u381 (
    .a(_al_u318_o),
    .b(_al_u332_o),
    .c(_al_u336_o),
    .d(_al_u322_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u381_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(~D*~A)))"),
    .INIT(16'hc0d0))
    _al_u382 (
    .a(\ADD02/ADD02/ADD01/n1 ),
    .b(_al_u353_o),
    .c(_al_u381_o),
    .d(\ADD02/ADD02/ADD01/g1 ),
    .o(_al_u382_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u383 (
    .a(_al_u358_o),
    .b(_al_u360_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD02/ADD02/g0 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~((D@C))+~(A)*B*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C))"),
    .INIT(16'hd44d))
    _al_u384 (
    .a(\ADD02/ADD02/ADD02/g0 ),
    .b(_al_u369_o),
    .c(_al_u371_o),
    .d(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u384_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(~C*~(B*~A)))"),
    .INIT(16'hf40b))
    _al_u385 (
    .a(_al_u365_o),
    .b(_al_u300_o),
    .c(_al_u366_o),
    .d(\M04/M01/M01/invSL_lutinv ),
    .o(new_M2[14]));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+~(A)*B*C*D*E)"),
    .INIT(32'h40dcc4fd))
    _al_u386 (
    .a(_al_u384_o),
    .b(new_M2[15]),
    .c(new_M2[14]),
    .d(_al_u378_o),
    .e(_al_u363_o),
    .o(_al_u386_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u387 (
    .a(_al_u140_o),
    .b(exp_diff[3]),
    .c(\exp_diff[4]_neg_lutinv ),
    .o(_al_u387_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(B*A))"),
    .INIT(16'h0777))
    _al_u388 (
    .a(_al_u387_o),
    .b(_al_u319_o),
    .c(_al_u78_o),
    .d(n2[18]),
    .o(_al_u388_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u389 (
    .a(_al_u388_o),
    .b(\M04/M01/M01/invSL_lutinv ),
    .o(new_M2[18]));
  AL_MAP_LUT4 #(
    .EQN("(~C*(~D*~(A)*~(B)+~D*A*~(B)+~(~D)*A*B+~D*A*B))"),
    .INIT(16'h080b))
    _al_u390 (
    .a(n63_lutinv),
    .b(exp_diff[2]),
    .c(exp_diff[3]),
    .d(_al_u231_o),
    .o(_al_u390_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*A))"),
    .INIT(16'h7077))
    _al_u391 (
    .a(_al_u390_o),
    .b(_al_u297_o),
    .c(_al_u78_o),
    .d(n1[18]),
    .o(_al_u391_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u392 (
    .a(new_M2[18]),
    .b(_al_u391_o),
    .o(\ADD02/ADD03/ADD01/p2_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u393 (
    .a(_al_u301_o),
    .b(exp_diff[3]),
    .o(_al_u393_o));
  AL_MAP_LUT5 #(
    .EQN("(D@(~(E*C)*~(B*A)))"),
    .INIT(32'hf8078877))
    _al_u394 (
    .a(_al_u393_o),
    .b(_al_u300_o),
    .c(_al_u78_o),
    .d(\M04/M01/M01/invSL_lutinv ),
    .e(n2[17]),
    .o(new_M2[17]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~C)*~(B*A))"),
    .INIT(16'h7077))
    _al_u395 (
    .a(_al_u297_o),
    .b(_al_u167_o),
    .c(_al_u78_o),
    .d(n1[17]),
    .o(_al_u395_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u396 (
    .a(new_M2[17]),
    .b(_al_u395_o),
    .o(\ADD02/ADD03/ADD01/p1_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~(E*~D)*~(~C*~B*A))"),
    .INIT(32'hfd00fdfd))
    _al_u397 (
    .a(_al_u297_o),
    .b(_al_u330_o),
    .c(exp_diff[3]),
    .d(_al_u78_o),
    .e(n1[19]),
    .o(_al_u397_o));
  AL_MAP_LUT5 #(
    .EQN("(D@(~(E*C)*~(B*A)))"),
    .INIT(32'hf8078877))
    _al_u398 (
    .a(_al_u300_o),
    .b(_al_u205_o),
    .c(_al_u78_o),
    .d(\M04/M01/M01/invSL_lutinv ),
    .e(n2[19]),
    .o(new_M2[19]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u399 (
    .a(_al_u397_o),
    .b(new_M2[19]),
    .o(\ADD02/ADD03/ADD01/p3_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("~(E*~((~C*B*A))*~(D)+E*(~C*B*A)*~(D)+~(E)*(~C*B*A)*D+E*(~C*B*A)*D)"),
    .INIT(32'hf700f7ff))
    _al_u400 (
    .a(u194_sel_is_0_o),
    .b(_al_u310_o),
    .c(exp_diff[3]),
    .d(_al_u78_o),
    .e(n1[16]),
    .o(_al_u400_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*C)*~(~B*A))"),
    .INIT(16'h0ddd))
    _al_u401 (
    .a(_al_u387_o),
    .b(_al_u138_o),
    .c(_al_u78_o),
    .d(n2[16]),
    .o(_al_u401_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@B@A)"),
    .INIT(8'h69))
    _al_u402 (
    .a(_al_u400_o),
    .b(_al_u401_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD03/ADD01/p0_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u403 (
    .a(\ADD02/ADD03/ADD01/p2_lutinv ),
    .b(\ADD02/ADD03/ADD01/p1_lutinv ),
    .c(\ADD02/ADD03/ADD01/p3_lutinv ),
    .d(\ADD02/ADD03/ADD01/p0_lutinv ),
    .o(_al_u403_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~D*~(B*~(C*~A))))"),
    .INIT(32'hff8c0000))
    _al_u404 (
    .a(_al_u355_o),
    .b(_al_u380_o),
    .c(_al_u382_o),
    .d(_al_u386_o),
    .e(_al_u403_o),
    .o(_al_u404_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u405 (
    .a(_al_u400_o),
    .b(_al_u401_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD03/ADD01/g0 ));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+~(A)*B*C)"),
    .INIT(8'h71))
    _al_u406 (
    .a(\ADD02/ADD03/ADD01/g0 ),
    .b(new_M2[17]),
    .c(_al_u395_o),
    .o(_al_u406_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*B*C)"),
    .INIT(8'h4d))
    _al_u407 (
    .a(_al_u406_o),
    .b(new_M2[18]),
    .c(_al_u391_o),
    .o(_al_u407_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C)"),
    .INIT(8'hb2))
    _al_u408 (
    .a(_al_u407_o),
    .b(_al_u397_o),
    .c(new_M2[19]),
    .o(_al_u408_o));
  AL_MAP_LUT4 #(
    .EQN("~(D*~((B*A))*~(C)+D*(B*A)*~(C)+~(D)*(B*A)*C+D*(B*A)*C)"),
    .INIT(16'h707f))
    _al_u409 (
    .a(u194_sel_is_0_o),
    .b(n5_lutinv),
    .c(_al_u78_o),
    .d(n1[22]),
    .o(_al_u409_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D)*~(~C*B*A))"),
    .INIT(32'h00f7f7f7))
    _al_u410 (
    .a(_al_u300_o),
    .b(_al_u215_o),
    .c(_al_u171_o),
    .d(_al_u78_o),
    .e(n2[22]),
    .o(_al_u410_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@B@A)"),
    .INIT(8'h69))
    _al_u411 (
    .a(_al_u409_o),
    .b(_al_u410_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD03/ADD02/p2_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~(E*~D)*~(~C*B*A))"),
    .INIT(32'hf700f7f7))
    _al_u412 (
    .a(_al_u297_o),
    .b(_al_u166_o),
    .c(_al_u171_o),
    .d(_al_u78_o),
    .e(n1[21]),
    .o(_al_u412_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D)*~(C*~B*A))"),
    .INIT(32'h00dfdfdf))
    _al_u413 (
    .a(_al_u300_o),
    .b(_al_u171_o),
    .c(_al_u180_o),
    .d(_al_u78_o),
    .e(n2[21]),
    .o(_al_u413_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@B@A)"),
    .INIT(8'h69))
    _al_u414 (
    .a(_al_u412_o),
    .b(_al_u413_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD03/ADD02/p1_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~(E*~D)*~(~C*B*A))"),
    .INIT(32'hf700f7f7))
    _al_u415 (
    .a(_al_u297_o),
    .b(_al_u71_o),
    .c(_al_u171_o),
    .d(_al_u78_o),
    .e(n1[20]),
    .o(_al_u415_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*D)*~(~C*B*A))"),
    .INIT(32'h00f7f7f7))
    _al_u416 (
    .a(_al_u300_o),
    .b(_al_u134_o),
    .c(_al_u171_o),
    .d(_al_u78_o),
    .e(n2[20]),
    .o(_al_u416_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u417 (
    .a(_al_u415_o),
    .b(_al_u416_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD03/ADD02/g0 ));
  AL_MAP_LUT4 #(
    .EQN("(A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+~(A)*~(B)*~(C)*D+A*~(B)*~(C)*D+~(A)*B*~(C)*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'hc7f8))
    _al_u418 (
    .a(_al_u387_o),
    .b(n198_lutinv),
    .c(_al_u66_o),
    .d(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD03/ADD02/p3_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u419 (
    .a(\ADD02/ADD03/ADD02/p2_lutinv ),
    .b(\ADD02/ADD03/ADD02/p1_lutinv ),
    .c(\ADD02/ADD03/ADD02/g0 ),
    .d(\ADD02/ADD03/ADD02/p3_lutinv ),
    .o(\ADD02/ADD03/ADD02/n18 ));
  AL_MAP_LUT3 #(
    .EQN("(~A*(C@B))"),
    .INIT(8'h14))
    _al_u420 (
    .a(_al_u412_o),
    .b(_al_u413_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD03/ADD02/g1 ));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~((D@C))+~(A)*~(B)*(D@C)+A*~(B)*(D@C)+A*B*(D@C))"),
    .INIT(16'h2bb2))
    _al_u421 (
    .a(\ADD02/ADD03/ADD02/g1 ),
    .b(_al_u409_o),
    .c(_al_u410_o),
    .d(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD03/ADD02/n6_lutinv ));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*~(E@(B*A)))"),
    .INIT(32'h00080007))
    _al_u422 (
    .a(_al_u387_o),
    .b(n198_lutinv),
    .c(_al_u78_o),
    .d(_al_u66_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD03/ADD02/g3 ));
  AL_MAP_LUT5 #(
    .EQN("(~E*~C*~A*~(D*B))"),
    .INIT(32'h00000105))
    _al_u423 (
    .a(\ADD02/ADD03/ADD02/n18 ),
    .b(\ADD02/ADD03/ADD02/n6_lutinv ),
    .c(\ADD02/ADD03/ADD02/g3 ),
    .d(\ADD02/ADD03/ADD02/p3_lutinv ),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u423_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@B@A)"),
    .INIT(8'h69))
    _al_u424 (
    .a(_al_u415_o),
    .b(_al_u416_o),
    .c(\M04/M01/M01/invSL_lutinv ),
    .o(\ADD02/ADD03/ADD02/p0_lutinv ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u425 (
    .a(\ADD02/ADD03/ADD02/p1_lutinv ),
    .b(\ADD02/ADD03/ADD02/p0_lutinv ),
    .o(\ADD02/ADD03/ADD02/n3 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u426 (
    .a(\ADD02/ADD03/ADD02/n3 ),
    .b(\ADD02/ADD03/ADD02/p2_lutinv ),
    .c(\ADD02/ADD03/ADD02/p3_lutinv ),
    .o(\ADD02/ADD03/ADD02/n20 ));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*~A)))"),
    .INIT(16'h10f0))
    _al_u427 (
    .a(_al_u404_o),
    .b(_al_u408_o),
    .c(_al_u423_o),
    .d(\ADD02/ADD03/ADD02/n20 ),
    .o(_al_u427_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@(B*~A))"),
    .INIT(8'h4b))
    _al_u428 (
    .a(_al_u355_o),
    .b(_al_u382_o),
    .c(\ADD02/ADD02/ADD02/p0_lutinv ),
    .o(_al_u428_o));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*~A))"),
    .INIT(8'hb4))
    _al_u429 (
    .a(_al_u352_o),
    .b(_al_u427_o),
    .c(_al_u428_o),
    .o(M_result2[12]));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*A)"),
    .INIT(8'h02))
    _al_u430 (
    .a(_al_u347_o),
    .b(_al_u350_o),
    .c(_al_u351_o),
    .o(_al_u430_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u431 (
    .a(\ADD02/ADD02/ADD01/g1 ),
    .b(\ADD02/ADD02/ADD01/g2 ),
    .o(_al_u431_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u432 (
    .a(_al_u431_o),
    .b(\ADD02/ADD02/ADD01/n1 ),
    .o(_al_u432_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@(~E*~(B*~(C*~A))))"),
    .INIT(32'h00ff738c))
    _al_u433 (
    .a(_al_u296_o),
    .b(_al_u432_o),
    .c(\ADD02/ADD02/ADD01/n3 ),
    .d(_al_u337_o),
    .e(_al_u323_o),
    .o(_al_u433_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~B*~(C*~(~D*~A))))"),
    .INIT(32'hfcec0000))
    _al_u434 (
    .a(_al_u257_o),
    .b(_al_u292_o),
    .c(_al_u294_o),
    .d(\ADD02/ADD01/ADD02/g0 ),
    .e(\ADD02/ADD02/ADD01/p0_lutinv ),
    .o(_al_u434_o));
  AL_MAP_LUT3 #(
    .EQN("~(B@(~C*~A))"),
    .INIT(8'h36))
    _al_u435 (
    .a(_al_u434_o),
    .b(\ADD02/ADD02/ADD01/p1_lutinv ),
    .c(\ADD02/ADD02/ADD01/g0 ),
    .o(_al_u435_o));
  AL_MAP_LUT5 #(
    .EQN("(C@(A*~(~E*~D*B)))"),
    .INIT(32'h5a5a5ad2))
    _al_u436 (
    .a(_al_u427_o),
    .b(_al_u430_o),
    .c(_al_u433_o),
    .d(_al_u328_o),
    .e(_al_u435_o),
    .o(M_result2[11]));
  AL_MAP_LUT4 #(
    .EQN("(C@(A*~(~D*B)))"),
    .INIT(16'h5ad2))
    _al_u437 (
    .a(_al_u427_o),
    .b(_al_u430_o),
    .c(_al_u328_o),
    .d(_al_u435_o),
    .o(M_result2[10]));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~C*~B*A))"),
    .INIT(16'hfd00))
    _al_u438 (
    .a(_al_u347_o),
    .b(_al_u350_o),
    .c(_al_u351_o),
    .d(_al_u423_o),
    .o(_al_u438_o));
  AL_MAP_LUT5 #(
    .EQN("(C@(A*~(E*~(~D*~B))))"),
    .INIT(32'hf0d25a5a))
    _al_u439 (
    .a(_al_u438_o),
    .b(_al_u404_o),
    .c(_al_u435_o),
    .d(_al_u408_o),
    .e(\ADD02/ADD03/ADD02/n20 ),
    .o(M_result2[9]));
  AL_MAP_LUT3 #(
    .EQN("(C*~(~B*A))"),
    .INIT(8'hd0))
    _al_u440 (
    .a(_al_u347_o),
    .b(_al_u350_o),
    .c(_al_u423_o),
    .o(_al_u440_o));
  AL_MAP_LUT5 #(
    .EQN("(D@(A*~(E*~(~C*~B))))"),
    .INIT(32'hfd0255aa))
    _al_u441 (
    .a(_al_u440_o),
    .b(_al_u404_o),
    .c(_al_u408_o),
    .d(_al_u351_o),
    .e(\ADD02/ADD03/ADD02/n20 ),
    .o(M_result2[8]));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u442 (
    .a(\ADD02/ADD01/ADD02/g1 ),
    .b(\ADD02/ADD01/ADD02/p1_lutinv ),
    .c(\ADD02/ADD01/ADD02/g0 ),
    .o(_al_u442_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@(B*~A))"),
    .INIT(8'h4b))
    _al_u443 (
    .a(_al_u345_o),
    .b(_al_u442_o),
    .c(\ADD02/ADD01/ADD02/p2_lutinv ),
    .o(_al_u443_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~(D*C*~A))"),
    .INIT(16'h8ccc))
    _al_u444 (
    .a(_al_u443_o),
    .b(_al_u423_o),
    .c(_al_u341_o),
    .d(_al_u345_o),
    .o(_al_u444_o));
  AL_MAP_LUT5 #(
    .EQN("(C@(B*~(E*~(~D*~A))))"),
    .INIT(32'hf0b43c3c))
    _al_u445 (
    .a(_al_u404_o),
    .b(_al_u444_o),
    .c(_al_u350_o),
    .d(_al_u408_o),
    .e(\ADD02/ADD03/ADD02/n20 ),
    .o(M_result2[7]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u446 (
    .a(_al_u423_o),
    .b(_al_u341_o),
    .c(_al_u345_o),
    .o(_al_u446_o));
  AL_MAP_LUT5 #(
    .EQN("(D@(B*~(E*~(~C*~A))))"),
    .INIT(32'hfb0433cc))
    _al_u447 (
    .a(_al_u404_o),
    .b(_al_u446_o),
    .c(_al_u408_o),
    .d(_al_u443_o),
    .e(\ADD02/ADD03/ADD02/n20 ),
    .o(M_result2[6]));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u448 (
    .a(_al_u423_o),
    .b(_al_u341_o),
    .c(\ADD02/ADD01/ADD02/p0_lutinv ),
    .o(_al_u448_o));
  AL_MAP_LUT3 #(
    .EQN("(B@(~C*~A))"),
    .INIT(8'hc9))
    _al_u449 (
    .a(_al_u257_o),
    .b(\ADD02/ADD01/ADD02/p1_lutinv ),
    .c(\ADD02/ADD01/ADD02/g0 ),
    .o(_al_u449_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@(B*~(E*~(~C*~A))))"),
    .INIT(32'h04fbcc33))
    _al_u450 (
    .a(_al_u404_o),
    .b(_al_u448_o),
    .c(_al_u408_o),
    .d(_al_u449_o),
    .e(\ADD02/ADD03/ADD02/n20 ),
    .o(M_result2[5]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u451 (
    .a(_al_u423_o),
    .b(_al_u341_o),
    .o(_al_u451_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u452 (
    .a(_al_u348_o),
    .b(\ADD02/ADD01/ADD02/p0_lutinv ),
    .o(_al_u452_o));
  AL_MAP_LUT5 #(
    .EQN("(D@(B*~(E*~(~C*~A))))"),
    .INIT(32'hfb0433cc))
    _al_u453 (
    .a(_al_u404_o),
    .b(_al_u451_o),
    .c(_al_u408_o),
    .d(_al_u452_o),
    .e(\ADD02/ADD03/ADD02/n20 ),
    .o(M_result2[4]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u454 (
    .a(_al_u195_o),
    .b(_al_u255_o),
    .o(_al_u454_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u455 (
    .a(_al_u454_o),
    .b(_al_u339_o),
    .o(_al_u455_o));
  AL_MAP_LUT5 #(
    .EQN("(D*~C*~(E*~(~B*~A)))"),
    .INIT(32'h01000f00))
    _al_u456 (
    .a(_al_u404_o),
    .b(_al_u408_o),
    .c(_al_u455_o),
    .d(_al_u423_o),
    .e(\ADD02/ADD03/ADD02/n20 ),
    .o(_al_u456_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(~B*~(C*~A)))"),
    .INIT(16'hdc23))
    _al_u457 (
    .a(_al_u195_o),
    .b(\ADD02/ADD01/ADD01/g2 ),
    .c(_al_u255_o),
    .d(\ADD02/ADD01/ADD01/p3_lutinv ),
    .o(_al_u457_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u458 (
    .a(_al_u456_o),
    .b(_al_u457_o),
    .o(M_result2[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u459 (
    .a(_al_u423_o),
    .b(_al_u339_o),
    .o(_al_u459_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(B*~(D*~(~C*~A))))"),
    .INIT(32'hfb3304cc))
    _al_u460 (
    .a(_al_u404_o),
    .b(_al_u459_o),
    .c(_al_u408_o),
    .d(\ADD02/ADD03/ADD02/n20 ),
    .e(_al_u454_o),
    .o(M_result2[2]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u461 (
    .a(_al_u423_o),
    .b(M_result[0]),
    .o(_al_u461_o));
  AL_MAP_LUT5 #(
    .EQN("(D@C@(~B*(E@A)))"),
    .INIT(32'h1ee12dd2))
    _al_u462 (
    .a(_al_u144_o),
    .b(_al_u145_o),
    .c(_al_u169_o),
    .d(_al_u193_o),
    .e(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u462_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(B*~(D*~(~C*~A))))"),
    .INIT(32'hfb3304cc))
    _al_u463 (
    .a(_al_u404_o),
    .b(_al_u461_o),
    .c(_al_u408_o),
    .d(\ADD02/ADD03/ADD02/n20 ),
    .e(_al_u462_o),
    .o(M_result2[1]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u464 (
    .a(_al_u328_o),
    .b(_al_u347_o),
    .c(_al_u350_o),
    .d(_al_u351_o),
    .o(_al_u464_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@(~C*~(D*~(B*~A))))"),
    .INIT(32'h040ffbf0))
    _al_u465 (
    .a(_al_u355_o),
    .b(_al_u382_o),
    .c(\ADD02/ADD02/ADD02/g0 ),
    .d(\ADD02/ADD02/ADD02/p0_lutinv ),
    .e(\ADD02/ADD02/ADD02/p1_lutinv ),
    .o(_al_u465_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(B*~(D*~C*A)))"),
    .INIT(32'h3b33c4cc))
    _al_u466 (
    .a(_al_u464_o),
    .b(_al_u427_o),
    .c(_al_u428_o),
    .d(_al_u338_o),
    .e(_al_u465_o),
    .o(M_result2[13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u467 (
    .a(_al_u347_o),
    .b(\ADD02/ADD02/ADD01/p2_lutinv ),
    .o(_al_u467_o));
  AL_MAP_LUT5 #(
    .EQN("(~((B*~A))*~(C)*~(D)*~(E)+~((B*~A))*C*~(D)*~(E)+(B*~A)*C*~(D)*~(E)+~((B*~A))*~(C)*D*~(E)+(B*~A)*~(C)*D*~(E)+~((B*~A))*C*D*~(E)+(B*~A)*C*D*~(E)+~((B*~A))*~(C)*~(D)*E+(B*~A)*~(C)*~(D)*E+~((B*~A))*C*~(D)*E+(B*~A)*~(C)*D*E+(B*~A)*C*D*E)"),
    .INIT(32'h44bffffb))
    _al_u468 (
    .a(_al_u355_o),
    .b(_al_u382_o),
    .c(\ADD02/ADD02/ADD02/g0 ),
    .d(\ADD02/ADD02/ADD02/p0_lutinv ),
    .e(\ADD02/ADD02/ADD02/p1_lutinv ),
    .o(_al_u468_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    _al_u469 (
    .a(_al_u467_o),
    .b(_al_u338_o),
    .c(_al_u468_o),
    .d(_al_u350_o),
    .e(_al_u351_o),
    .o(_al_u469_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@(C*~(~E*~(B*~A))))"),
    .INIT(32'hf00f40bf))
    _al_u470 (
    .a(_al_u355_o),
    .b(_al_u382_o),
    .c(_al_u384_o),
    .d(\ADD02/ADD02/ADD02/p2_lutinv ),
    .e(_al_u468_o),
    .o(_al_u470_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*B*C)"),
    .INIT(8'h4d))
    _al_u471 (
    .a(_al_u384_o),
    .b(new_M2[14]),
    .c(_al_u363_o),
    .o(_al_u471_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@(~C*~(D*~(B*~A))))"),
    .INIT(32'h040ffbf0))
    _al_u472 (
    .a(_al_u355_o),
    .b(_al_u382_o),
    .c(_al_u471_o),
    .d(\ADD02/ADD02/ADD02/n10 ),
    .e(\ADD02/ADD02/ADD02/p3_lutinv ),
    .o(_al_u472_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(B*~(~C*A)))"),
    .INIT(16'h3bc4))
    _al_u473 (
    .a(_al_u469_o),
    .b(_al_u427_o),
    .c(_al_u470_o),
    .d(_al_u472_o),
    .o(M_result2[15]));
  AL_MAP_LUT5 #(
    .EQN("(D@(B*~(~E*C*A)))"),
    .INIT(32'h33ccb34c))
    _al_u474 (
    .a(_al_u464_o),
    .b(_al_u427_o),
    .c(_al_u338_o),
    .d(_al_u470_o),
    .e(_al_u468_o),
    .o(M_result2[14]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~A*~(D*B))"),
    .INIT(16'h0105))
    _al_u475 (
    .a(\ADD02/ADD03/ADD02/n18 ),
    .b(\ADD02/ADD03/ADD02/n6_lutinv ),
    .c(\ADD02/ADD03/ADD02/g3 ),
    .d(\ADD02/ADD03/ADD02/p3_lutinv ),
    .o(_al_u475_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~(~B*~A)))"),
    .INIT(16'h10f0))
    _al_u476 (
    .a(_al_u404_o),
    .b(_al_u408_o),
    .c(_al_u475_o),
    .d(\ADD02/ADD03/ADD02/n20 ),
    .o(_al_u476_o));
  AL_MAP_LUT3 #(
    .EQN("~(~B*~(C)*~(A)+~B*C*~(A)+~(~B)*C*A+~B*C*A)"),
    .INIT(8'h4e))
    _al_u477 (
    .a(_al_u476_o),
    .b(n1[31]),
    .c(n2[31]),
    .o(result[31]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u478 (
    .a(_al_u470_o),
    .b(_al_u472_o),
    .o(_al_u478_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~(B*~(C*~A)))"),
    .INIT(16'h0073))
    _al_u479 (
    .a(_al_u355_o),
    .b(_al_u380_o),
    .c(_al_u382_o),
    .d(_al_u386_o),
    .o(_al_u479_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@D@(C*~(B*A)))"),
    .INIT(32'h8f70708f))
    _al_u480 (
    .a(_al_u469_o),
    .b(_al_u478_o),
    .c(_al_u427_o),
    .d(_al_u479_o),
    .e(\ADD02/ADD03/ADD01/p0_lutinv ),
    .o(M_result2[16]));
  AL_MAP_LUT4 #(
    .EQN("~(B@(~C*~(D*~A)))"),
    .INIT(16'h393c))
    _al_u481 (
    .a(_al_u479_o),
    .b(\ADD02/ADD03/ADD01/p1_lutinv ),
    .c(\ADD02/ADD03/ADD01/g0 ),
    .d(\ADD02/ADD03/ADD01/p0_lutinv ),
    .o(_al_u481_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(~D*~(B*~(C*~A))))"),
    .INIT(32'hff8c0073))
    _al_u482 (
    .a(_al_u355_o),
    .b(_al_u380_o),
    .c(_al_u382_o),
    .d(_al_u386_o),
    .e(\ADD02/ADD03/ADD01/p0_lutinv ),
    .o(_al_u482_o));
  AL_MAP_LUT5 #(
    .EQN("(D@(C*~(E*B*A)))"),
    .INIT(32'h8f700ff0))
    _al_u483 (
    .a(_al_u469_o),
    .b(_al_u478_o),
    .c(_al_u427_o),
    .d(_al_u481_o),
    .e(_al_u482_o),
    .o(M_result2[17]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u484 (
    .a(\ADD02/ADD03/ADD01/p1_lutinv ),
    .b(\ADD02/ADD03/ADD01/p0_lutinv ),
    .o(\ADD02/ADD03/ADD01/n3 ));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u485 (
    .a(\ADD02/ADD03/ADD01/n3 ),
    .b(\ADD02/ADD03/ADD01/p2_lutinv ),
    .o(_al_u485_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~(~D*~(B*~(C*~A))))"),
    .INIT(32'hff8c0000))
    _al_u486 (
    .a(_al_u355_o),
    .b(_al_u380_o),
    .c(_al_u382_o),
    .d(_al_u386_o),
    .e(\ADD02/ADD03/ADD01/n3 ),
    .o(_al_u486_o));
  AL_MAP_LUT4 #(
    .EQN("~(D@(~B*~(C*A)))"),
    .INIT(16'h13ec))
    _al_u487 (
    .a(_al_u486_o),
    .b(_al_u407_o),
    .c(\ADD02/ADD03/ADD01/p2_lutinv ),
    .d(\ADD02/ADD03/ADD01/p3_lutinv ),
    .o(_al_u487_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(C*~(D*B*A)))"),
    .INIT(32'h8f0f70f0))
    _al_u488 (
    .a(_al_u469_o),
    .b(_al_u478_o),
    .c(_al_u427_o),
    .d(_al_u485_o),
    .e(_al_u487_o),
    .o(M_result2[19]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u489 (
    .a(\ADD02/ADD03/ADD01/p1_lutinv ),
    .b(\ADD02/ADD03/ADD01/p0_lutinv ),
    .o(_al_u489_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@(B*~A))"),
    .INIT(8'h4b))
    _al_u490 (
    .a(_al_u486_o),
    .b(_al_u406_o),
    .c(\ADD02/ADD03/ADD01/p2_lutinv ),
    .o(_al_u490_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(C*~(D*B*A)))"),
    .INIT(32'h8f0f70f0))
    _al_u491 (
    .a(_al_u469_o),
    .b(_al_u478_o),
    .c(_al_u427_o),
    .d(_al_u489_o),
    .e(_al_u490_o),
    .o(M_result2[18]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u492 (
    .a(\ADD02/ADD03/ADD01/p2_lutinv ),
    .b(\ADD02/ADD03/ADD01/p3_lutinv ),
    .o(\ADD02/ADD03/ADD01/n14 ));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u493 (
    .a(\ADD02/ADD03/ADD01/n14 ),
    .b(\ADD02/ADD03/ADD01/p1_lutinv ),
    .c(\ADD02/ADD03/ADD01/p0_lutinv ),
    .o(_al_u493_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@(~B*~A))"),
    .INIT(8'h1e))
    _al_u494 (
    .a(_al_u404_o),
    .b(_al_u408_o),
    .c(\ADD02/ADD03/ADD02/p0_lutinv ),
    .o(_al_u494_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(D*~(C*B*A)))"),
    .INIT(32'h80ff7f00))
    _al_u495 (
    .a(_al_u493_o),
    .b(_al_u469_o),
    .c(_al_u478_o),
    .d(_al_u427_o),
    .e(_al_u494_o),
    .o(M_result2[20]));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*B*A)"),
    .INIT(32'h00000080))
    _al_u496 (
    .a(_al_u469_o),
    .b(_al_u489_o),
    .c(\ADD02/ADD03/ADD01/n14 ),
    .d(_al_u470_o),
    .e(_al_u472_o),
    .o(_al_u496_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~(~B*~A)))"),
    .INIT(16'h010f))
    _al_u497 (
    .a(_al_u404_o),
    .b(_al_u408_o),
    .c(\ADD02/ADD03/ADD02/g0 ),
    .d(\ADD02/ADD03/ADD02/p0_lutinv ),
    .o(_al_u497_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@D@(B*~(~C*A)))"),
    .INIT(32'h3bc4c43b))
    _al_u498 (
    .a(_al_u496_o),
    .b(_al_u427_o),
    .c(_al_u494_o),
    .d(_al_u497_o),
    .e(\ADD02/ADD03/ADD02/p1_lutinv ),
    .o(M_result2[21]));
  AL_MAP_LUT5 #(
    .EQN("(E@(~B*~(D*C*~A)))"),
    .INIT(32'hdccc2333))
    _al_u499 (
    .a(_al_u497_o),
    .b(\ADD02/ADD03/ADD02/n6_lutinv ),
    .c(\ADD02/ADD03/ADD02/p2_lutinv ),
    .d(\ADD02/ADD03/ADD02/p1_lutinv ),
    .e(\ADD02/ADD03/ADD02/p3_lutinv ),
    .o(_al_u499_o));
  AL_MAP_LUT5 #(
    .EQN("(~((~B*~A))*~(C)*~(D)*~(E)+~((~B*~A))*C*~(D)*~(E)+(~B*~A)*C*~(D)*~(E)+~((~B*~A))*~(C)*D*~(E)+(~B*~A)*~(C)*D*~(E)+~((~B*~A))*C*D*~(E)+~((~B*~A))*~(C)*~(D)*E+(~B*~A)*~(C)*~(D)*E+(~B*~A)*C*~(D)*E+~((~B*~A))*~(C)*D*E+(~B*~A)*~(C)*D*E+(~B*~A)*C*D*E)"),
    .INIT(32'h1f1feffe))
    _al_u500 (
    .a(_al_u404_o),
    .b(_al_u408_o),
    .c(\ADD02/ADD03/ADD02/p1_lutinv ),
    .d(\ADD02/ADD03/ADD02/g0 ),
    .e(\ADD02/ADD03/ADD02/p0_lutinv ),
    .o(_al_u500_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u501 (
    .a(\ADD02/ADD03/ADD02/g1 ),
    .b(\ADD02/ADD03/ADD02/p1_lutinv ),
    .c(\ADD02/ADD03/ADD02/g0 ),
    .o(_al_u501_o));
  AL_MAP_LUT5 #(
    .EQN("~(E@(C*~(D*~(~B*~A))))"),
    .INIT(32'h10f0ef0f))
    _al_u502 (
    .a(_al_u404_o),
    .b(_al_u408_o),
    .c(_al_u501_o),
    .d(\ADD02/ADD03/ADD02/n3 ),
    .e(\ADD02/ADD03/ADD02/p2_lutinv ),
    .o(_al_u502_o));
  AL_MAP_LUT5 #(
    .EQN("(~(B)*~(C)*~((~E*~D*A))+B*C*~((~E*~D*A))+~(B)*~(C)*(~E*~D*A)+~(B)*C*(~E*~D*A)+B*C*(~E*~D*A))"),
    .INIT(32'hc3c3c3e3))
    _al_u503 (
    .a(_al_u496_o),
    .b(_al_u499_o),
    .c(_al_u427_o),
    .d(_al_u500_o),
    .e(_al_u502_o),
    .o(M_result2[23]));
  AL_MAP_LUT4 #(
    .EQN("(D@(B*~(~C*A)))"),
    .INIT(16'h3bc4))
    _al_u504 (
    .a(_al_u496_o),
    .b(_al_u427_o),
    .c(_al_u500_o),
    .d(_al_u502_o),
    .o(M_result2[22]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u505 (
    .a(_al_u476_o),
    .b(\M04/M01/M01/invSL_lutinv ),
    .o(_al_u505_o));
  AL_MAP_LUT4 #(
    .EQN("((D*B)*~(A)*~(C)+(D*B)*A*~(C)+~((D*B))*A*C+(D*B)*A*C)"),
    .INIT(16'haca0))
    _al_u506 (
    .a(\NM/n4 [0]),
    .b(M_result2[23]),
    .c(_al_u505_o),
    .d(M_result[0]),
    .o(result[0]));
  AL_MAP_LUT5 #(
    .EQN("(~(B)*~(C)*~((~D*A))*~(E)+B*~(C)*~((~D*A))*~(E)+B*C*~((~D*A))*~(E)+~(B)*~(C)*(~D*A)*~(E)+B*~(C)*(~D*A)*~(E)+~(B)*C*(~D*A)*~(E)+B*C*(~D*A)*~(E)+~(B)*~(C)*~((~D*A))*E+~(B)*C*~((~D*A))*E+B*C*~((~D*A))*E+~(B)*~(C)*(~D*A)*E+B*C*(~D*A)*E)"),
    .INIT(32'hf3d3cfef))
    _al_u507 (
    .a(_al_u496_o),
    .b(_al_u499_o),
    .c(_al_u427_o),
    .d(_al_u500_o),
    .e(_al_u502_o),
    .o(_al_u507_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'h4c5f))
    _al_u508 (
    .a(M_result2[23]),
    .b(_al_u507_o),
    .c(M_result2[1]),
    .d(M_result[0]),
    .o(_al_u508_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'ha3))
    _al_u509 (
    .a(\NM/n4 [1]),
    .b(_al_u508_o),
    .c(_al_u505_o),
    .o(result[1]));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C)"),
    .INIT(8'hbd))
    _al_u510 (
    .a(_al_u499_o),
    .b(_al_u427_o),
    .c(_al_u502_o),
    .o(_al_u510_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u511 (
    .a(M_result2[21]),
    .b(_al_u510_o),
    .o(_al_u511_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u512 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[2]),
    .d(M_result[0]),
    .o(_al_u512_o));
  AL_MAP_LUT5 #(
    .EQN("(~(B*~(E*~C))*~(A)*~(D)+~(B*~(E*~C))*A*~(D)+~(~(B*~(E*~C)))*A*D+~(B*~(E*~C))*A*D)"),
    .INIT(32'haa3faa33))
    _al_u513 (
    .a(\NM/n4 [2]),
    .b(_al_u512_o),
    .c(_al_u507_o),
    .d(_al_u505_o),
    .e(M_result2[1]),
    .o(result[2]));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u514 (
    .a(M_result2[21]),
    .b(_al_u510_o),
    .o(_al_u514_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u515 (
    .a(_al_u514_o),
    .b(M_result2[20]),
    .o(_al_u515_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u516 (
    .a(_al_u515_o),
    .b(_al_u511_o),
    .c(M_result2[1]),
    .d(M_result[0]),
    .o(_al_u516_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*~B)*~(C*A))"),
    .INIT(16'h4c5f))
    _al_u517 (
    .a(M_result2[23]),
    .b(_al_u507_o),
    .c(M_result2[3]),
    .d(M_result2[2]),
    .o(_al_u517_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(A)*~(D)+~(C*B)*A*~(D)+~(~(C*B))*A*D+~(C*B)*A*D)"),
    .INIT(16'haa3f))
    _al_u518 (
    .a(\NM/n4 [3]),
    .b(_al_u516_o),
    .c(_al_u517_o),
    .d(_al_u505_o),
    .o(result[3]));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*B)*~(E*A))"),
    .INIT(32'h0105030f))
    _al_u519 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(_al_u505_o),
    .d(M_result2[4]),
    .e(M_result2[2]),
    .o(_al_u519_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~(E*D*B*A))"),
    .INIT(32'h70f0f0f0))
    _al_u520 (
    .a(_al_u469_o),
    .b(_al_u478_o),
    .c(_al_u427_o),
    .d(_al_u489_o),
    .e(\ADD02/ADD03/ADD01/n14 ),
    .o(_al_u520_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u521 (
    .a(_al_u497_o),
    .b(\ADD02/ADD03/ADD02/p1_lutinv ),
    .o(_al_u521_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(~(B)*~(C)*~(D)+B*C*D))"),
    .INIT(16'h4001))
    _al_u522 (
    .a(_al_u510_o),
    .b(_al_u520_o),
    .c(_al_u521_o),
    .d(_al_u494_o),
    .o(_al_u522_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u523 (
    .a(_al_u522_o),
    .b(M_result2[19]),
    .o(_al_u523_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*~C)*~(E*B))"),
    .INIT(32'h2022a0aa))
    _al_u524 (
    .a(_al_u519_o),
    .b(_al_u523_o),
    .c(_al_u507_o),
    .d(M_result2[3]),
    .e(M_result[0]),
    .o(_al_u524_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~(E*C)*B)*~(D*~A))"),
    .INIT(32'ha2f32233))
    _al_u525 (
    .a(\NM/n4 [4]),
    .b(_al_u524_o),
    .c(_al_u515_o),
    .d(_al_u505_o),
    .e(M_result2[1]),
    .o(result[4]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u526 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[3]),
    .d(M_result2[5]),
    .o(_al_u526_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u527 (
    .a(_al_u526_o),
    .b(_al_u507_o),
    .c(M_result2[4]),
    .o(_al_u527_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u528 (
    .a(_al_u515_o),
    .b(_al_u523_o),
    .c(M_result2[2]),
    .d(M_result2[1]),
    .o(_al_u528_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C+~(A)*B*C)"),
    .INIT(8'h7e))
    _al_u529 (
    .a(_al_u427_o),
    .b(_al_u487_o),
    .c(_al_u494_o),
    .o(_al_u529_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u530 (
    .a(M_result2[21]),
    .b(_al_u510_o),
    .c(_al_u529_o),
    .d(M_result2[18]),
    .o(_al_u530_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u531 (
    .a(_al_u527_o),
    .b(_al_u528_o),
    .c(_al_u530_o),
    .d(M_result[0]),
    .o(_al_u531_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'ha3))
    _al_u532 (
    .a(\NM/n4 [5]),
    .b(_al_u531_o),
    .c(_al_u505_o),
    .o(result[5]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u533 (
    .a(M_result2[23]),
    .b(M_result2[6]),
    .o(_al_u533_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(D*~C)*~(E*A))"),
    .INIT(32'h10113033))
    _al_u534 (
    .a(_al_u511_o),
    .b(_al_u533_o),
    .c(_al_u507_o),
    .d(M_result2[5]),
    .e(M_result2[4]),
    .o(_al_u534_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C+~(A)*B*C)"),
    .INIT(8'h7e))
    _al_u535 (
    .a(_al_u427_o),
    .b(_al_u490_o),
    .c(_al_u487_o),
    .o(_al_u535_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u536 (
    .a(_al_u522_o),
    .b(_al_u535_o),
    .c(M_result2[17]),
    .o(_al_u536_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(E*C)*~(D*A))"),
    .INIT(32'h040c44cc))
    _al_u537 (
    .a(_al_u515_o),
    .b(_al_u534_o),
    .c(_al_u536_o),
    .d(M_result2[3]),
    .e(M_result[0]),
    .o(_al_u537_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u538 (
    .a(_al_u523_o),
    .b(_al_u530_o),
    .c(M_result2[2]),
    .d(M_result2[1]),
    .o(_al_u538_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(A)*~(D)+~(C*B)*A*~(D)+~(~(C*B))*A*D+~(C*B)*A*D)"),
    .INIT(16'haa3f))
    _al_u539 (
    .a(\NM/n4 [6]),
    .b(_al_u537_o),
    .c(_al_u538_o),
    .d(_al_u505_o),
    .o(result[6]));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u540 (
    .a(_al_u514_o),
    .b(_al_u529_o),
    .o(_al_u540_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*(~(B)*~(C)*~(D)+B*C*D))"),
    .INIT(16'h4001))
    _al_u541 (
    .a(M_result2[17]),
    .b(_al_u490_o),
    .c(_al_u487_o),
    .d(_al_u427_o),
    .o(_al_u541_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*A)"),
    .INIT(32'h00020000))
    _al_u542 (
    .a(_al_u541_o),
    .b(M_result2[21]),
    .c(_al_u510_o),
    .d(M_result2[20]),
    .e(M_result2[16]),
    .o(_al_u542_o));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u543 (
    .a(M_result2[18]),
    .b(M_result2[2]),
    .o(_al_u543_o));
  AL_MAP_LUT5 #(
    .EQN("(~(E*B)*~(D*C*A))"),
    .INIT(32'h13335fff))
    _al_u544 (
    .a(_al_u540_o),
    .b(_al_u542_o),
    .c(_al_u543_o),
    .d(M_result2[17]),
    .e(M_result2[1]),
    .o(_al_u544_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C+~(A)*B*C)"),
    .INIT(8'h7e))
    _al_u545 (
    .a(_al_u520_o),
    .b(_al_u521_o),
    .c(_al_u494_o),
    .o(_al_u545_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u546 (
    .a(_al_u545_o),
    .b(_al_u541_o),
    .c(_al_u510_o),
    .d(M_result2[16]),
    .o(_al_u546_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u547 (
    .a(_al_u546_o),
    .b(M_result2[15]),
    .c(M_result[0]),
    .o(_al_u547_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u548 (
    .a(_al_u544_o),
    .b(_al_u547_o),
    .c(_al_u530_o),
    .d(M_result2[3]),
    .o(_al_u548_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u549 (
    .a(M_result2[23]),
    .b(M_result2[8]),
    .o(_al_u549_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(D*B)*~(E*A))"),
    .INIT(32'h0105030f))
    _al_u550 (
    .a(_al_u515_o),
    .b(_al_u511_o),
    .c(_al_u549_o),
    .d(M_result2[6]),
    .e(M_result2[5]),
    .o(_al_u550_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u551 (
    .a(_al_u523_o),
    .b(_al_u507_o),
    .c(M_result2[7]),
    .d(M_result2[4]),
    .o(_al_u551_o));
  AL_MAP_LUT5 #(
    .EQN("(~(D*C*B)*~(A)*~(E)+~(D*C*B)*A*~(E)+~(~(D*C*B))*A*E+~(D*C*B)*A*E)"),
    .INIT(32'haaaa3fff))
    _al_u552 (
    .a(\NM/n4 [8]),
    .b(_al_u548_o),
    .c(_al_u550_o),
    .d(_al_u551_o),
    .e(_al_u505_o),
    .o(result[8]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*A)"),
    .INIT(16'h0200))
    _al_u553 (
    .a(_al_u522_o),
    .b(_al_u535_o),
    .c(M_result2[17]),
    .d(M_result2[16]),
    .o(_al_u553_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u554 (
    .a(_al_u515_o),
    .b(_al_u553_o),
    .c(M_result2[4]),
    .d(M_result[0]),
    .o(_al_u554_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u555 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[7]),
    .d(M_result2[5]),
    .o(_al_u555_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u556 (
    .a(_al_u554_o),
    .b(_al_u555_o),
    .c(_al_u507_o),
    .d(M_result2[6]),
    .o(_al_u556_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u557 (
    .a(_al_u514_o),
    .b(M_result2[20]),
    .c(M_result2[19]),
    .o(_al_u557_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u558 (
    .a(_al_u557_o),
    .b(_al_u536_o),
    .c(M_result2[3]),
    .d(M_result2[1]),
    .o(_al_u558_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u559 (
    .a(_al_u514_o),
    .b(_al_u529_o),
    .c(M_result2[18]),
    .o(_al_u559_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u560 (
    .a(_al_u556_o),
    .b(_al_u558_o),
    .c(_al_u559_o),
    .d(M_result2[2]),
    .o(_al_u560_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'ha3))
    _al_u561 (
    .a(\NM/n4 [7]),
    .b(_al_u560_o),
    .c(_al_u505_o),
    .o(result[7]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u562 (
    .a(_al_u515_o),
    .b(_al_u507_o),
    .c(M_result2[8]),
    .d(M_result2[6]),
    .o(_al_u562_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u563 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[9]),
    .d(M_result2[7]),
    .o(_al_u563_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u564 (
    .a(_al_u562_o),
    .b(_al_u563_o),
    .c(_al_u536_o),
    .d(M_result2[3]),
    .o(_al_u564_o));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u565 (
    .a(_al_u479_o),
    .b(\ADD02/ADD03/ADD01/p0_lutinv ),
    .o(_al_u565_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C+A*B*C)"),
    .INIT(8'hbd))
    _al_u566 (
    .a(_al_u565_o),
    .b(_al_u481_o),
    .c(_al_u490_o),
    .o(_al_u566_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u567 (
    .a(_al_u566_o),
    .b(M_result2[16]),
    .o(_al_u567_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u568 (
    .a(_al_u540_o),
    .b(_al_u567_o),
    .c(M_result2[15]),
    .o(_al_u568_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u569 (
    .a(_al_u523_o),
    .b(_al_u542_o),
    .c(M_result2[5]),
    .d(M_result2[2]),
    .o(_al_u569_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(D*C)*~(E*A))"),
    .INIT(32'h04440ccc))
    _al_u570 (
    .a(_al_u568_o),
    .b(_al_u569_o),
    .c(_al_u530_o),
    .d(M_result2[4]),
    .e(M_result2[1]),
    .o(_al_u570_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u571 (
    .a(_al_u546_o),
    .b(M_result2[15]),
    .o(_al_u571_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u572 (
    .a(_al_u571_o),
    .b(M_result2[14]),
    .o(_al_u572_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u573 (
    .a(_al_u564_o),
    .b(_al_u570_o),
    .c(_al_u572_o),
    .d(M_result[0]),
    .o(_al_u573_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'ha3))
    _al_u574 (
    .a(\NM/n4 [9]),
    .b(_al_u573_o),
    .c(_al_u505_o),
    .o(result[9]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u575 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[11]),
    .d(M_result2[9]),
    .o(_al_u575_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(D*~C)*~(E*A))"),
    .INIT(32'h4044c0cc))
    _al_u576 (
    .a(_al_u515_o),
    .b(_al_u575_o),
    .c(_al_u507_o),
    .d(M_result2[10]),
    .e(M_result2[8]),
    .o(_al_u576_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u577 (
    .a(M_result2[21]),
    .b(_al_u510_o),
    .c(_al_u529_o),
    .d(M_result2[18]),
    .o(_al_u577_o));
  AL_MAP_LUT5 #(
    .EQN("(~((C*~(B*A)))*~(D)*~(E)+(C*~(B*A))*~(D)*~(E)+~((C*~(B*A)))*D*~(E)+(C*~(B*A))*~(D)*E+~((C*~(B*A)))*D*E+(C*~(B*A))*D*E)"),
    .INIT(32'hff708fff))
    _al_u578 (
    .a(_al_u469_o),
    .b(_al_u478_o),
    .c(_al_u427_o),
    .d(_al_u481_o),
    .e(_al_u482_o),
    .o(_al_u578_o));
  AL_MAP_LUT4 #(
    .EQN("((B*~A)*~(C)*~(D)+~((B*~A))*C*~(D)+(B*~A)*C*~(D)+~((B*~A))*~(C)*D+(B*~A)*~(C)*D+~((B*~A))*C*D)"),
    .INIT(16'hbff4))
    _al_u579 (
    .a(_al_u469_o),
    .b(_al_u427_o),
    .c(_al_u470_o),
    .d(_al_u472_o),
    .o(_al_u579_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u580 (
    .a(_al_u578_o),
    .b(_al_u579_o),
    .o(_al_u580_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u581 (
    .a(_al_u577_o),
    .b(_al_u580_o),
    .c(M_result2[13]),
    .o(_al_u581_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u582 (
    .a(_al_u576_o),
    .b(_al_u581_o),
    .c(_al_u536_o),
    .d(M_result2[5]),
    .e(M_result2[1]),
    .o(_al_u582_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u583 (
    .a(_al_u559_o),
    .b(_al_u557_o),
    .c(M_result2[7]),
    .d(M_result2[6]),
    .o(_al_u583_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u584 (
    .a(_al_u582_o),
    .b(_al_u583_o),
    .c(_al_u553_o),
    .d(M_result2[4]),
    .o(_al_u584_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u585 (
    .a(_al_u540_o),
    .b(_al_u567_o),
    .c(M_result2[15]),
    .d(M_result2[14]),
    .o(_al_u585_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C+~(A)*B*C)"),
    .INIT(8'h7e))
    _al_u586 (
    .a(_al_u427_o),
    .b(_al_u465_o),
    .c(_al_u470_o),
    .o(_al_u586_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u587 (
    .a(_al_u578_o),
    .b(M_result2[15]),
    .c(_al_u586_o),
    .o(_al_u587_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u588 (
    .a(_al_u577_o),
    .b(_al_u587_o),
    .c(M_result2[12]),
    .o(_al_u588_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u589 (
    .a(_al_u585_o),
    .b(_al_u588_o),
    .c(M_result2[2]),
    .d(M_result[0]),
    .o(_al_u589_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u590 (
    .a(_al_u584_o),
    .b(_al_u589_o),
    .c(_al_u568_o),
    .d(M_result2[3]),
    .o(_al_u590_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(A)*~(C)+~B*A*~(C)+~(~B)*A*C+~B*A*C)"),
    .INIT(8'ha3))
    _al_u591 (
    .a(\NM/n4 [11]),
    .b(_al_u590_o),
    .c(_al_u505_o),
    .o(result[11]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u592 (
    .a(_al_u542_o),
    .b(_al_u530_o),
    .c(M_result2[3]),
    .d(M_result2[5]),
    .o(_al_u592_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(D*C)*~(E*A))"),
    .INIT(32'h04440ccc))
    _al_u593 (
    .a(_al_u568_o),
    .b(_al_u592_o),
    .c(_al_u523_o),
    .d(M_result2[6]),
    .e(M_result2[2]),
    .o(_al_u593_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u594 (
    .a(_al_u515_o),
    .b(_al_u536_o),
    .c(M_result2[7]),
    .d(M_result2[4]),
    .o(_al_u594_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~(C*B)*~(E*A))"),
    .INIT(32'h0015003f))
    _al_u595 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[10]),
    .d(_al_u505_o),
    .e(M_result2[8]),
    .o(_al_u595_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u596 (
    .a(_al_u594_o),
    .b(_al_u595_o),
    .c(_al_u507_o),
    .d(M_result2[9]),
    .o(_al_u596_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u597 (
    .a(_al_u593_o),
    .b(_al_u596_o),
    .c(_al_u581_o),
    .d(M_result[0]),
    .o(_al_u597_o));
  AL_MAP_LUT5 #(
    .EQN("(~(~(E*C)*B)*~(D*~A))"),
    .INIT(32'ha2f32233))
    _al_u598 (
    .a(\NM/n4 [10]),
    .b(_al_u597_o),
    .c(_al_u572_o),
    .d(_al_u505_o),
    .e(M_result2[1]),
    .o(result[10]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u599 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[12]),
    .d(M_result2[10]),
    .o(_al_u599_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(D*~C)*~(E*A))"),
    .INIT(32'h4044c0cc))
    _al_u600 (
    .a(_al_u515_o),
    .b(_al_u599_o),
    .c(_al_u507_o),
    .d(M_result2[11]),
    .e(M_result2[9]),
    .o(_al_u600_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u601 (
    .a(_al_u600_o),
    .b(_al_u585_o),
    .c(_al_u536_o),
    .d(M_result2[3]),
    .e(M_result2[6]),
    .o(_al_u601_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u602 (
    .a(_al_u559_o),
    .b(_al_u557_o),
    .c(M_result2[8]),
    .d(M_result2[7]),
    .o(_al_u602_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u603 (
    .a(_al_u601_o),
    .b(_al_u602_o),
    .c(_al_u553_o),
    .d(M_result2[5]),
    .o(_al_u603_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u604 (
    .a(_al_u588_o),
    .b(_al_u581_o),
    .c(M_result2[2]),
    .d(M_result2[1]),
    .o(_al_u604_o));
  AL_MAP_LUT3 #(
    .EQN("(~(A)*~(B)*~(C)+A*~(B)*~(C)+~(A)*B*~(C)+A*~(B)*C+~(A)*B*C+A*B*C)"),
    .INIT(8'he7))
    _al_u605 (
    .a(_al_u427_o),
    .b(_al_u472_o),
    .c(_al_u482_o),
    .o(_al_u605_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u606 (
    .a(_al_u586_o),
    .b(_al_u605_o),
    .c(M_result2[12]),
    .d(M_result2[11]),
    .o(_al_u606_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u607 (
    .a(_al_u545_o),
    .b(_al_u541_o),
    .c(_al_u606_o),
    .d(_al_u510_o),
    .o(_al_u607_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u608 (
    .a(_al_u604_o),
    .b(_al_u568_o),
    .c(_al_u607_o),
    .d(M_result2[4]),
    .e(M_result[0]),
    .o(_al_u608_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(A)*~(D)+~(C*B)*A*~(D)+~(~(C*B))*A*D+~(C*B)*A*D)"),
    .INIT(16'haa3f))
    _al_u609 (
    .a(\NM/n4 [12]),
    .b(_al_u603_o),
    .c(_al_u608_o),
    .d(_al_u505_o),
    .o(result[12]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u610 (
    .a(_al_u515_o),
    .b(_al_u507_o),
    .c(M_result2[13]),
    .d(M_result2[11]),
    .o(_al_u610_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(D*B)*~(C*A))"),
    .INIT(32'h0000135f))
    _al_u611 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[12]),
    .d(M_result2[14]),
    .e(_al_u505_o),
    .o(_al_u611_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u612 (
    .a(_al_u610_o),
    .b(_al_u611_o),
    .c(_al_u536_o),
    .d(M_result2[8]),
    .o(_al_u612_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u613 (
    .a(_al_u612_o),
    .b(_al_u568_o),
    .c(_al_u530_o),
    .d(M_result2[9]),
    .e(M_result2[6]),
    .o(_al_u613_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u614 (
    .a(_al_u523_o),
    .b(_al_u542_o),
    .c(M_result2[10]),
    .d(M_result2[7]),
    .o(_al_u614_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    _al_u615 (
    .a(_al_u586_o),
    .b(_al_u605_o),
    .c(M_result2[12]),
    .d(M_result2[11]),
    .e(M_result2[10]),
    .o(_al_u615_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u616 (
    .a(_al_u522_o),
    .b(_al_u615_o),
    .c(_al_u541_o),
    .o(_al_u616_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    _al_u617 (
    .a(_al_u541_o),
    .b(_al_u606_o),
    .c(M_result2[21]),
    .d(_al_u510_o),
    .e(M_result2[20]),
    .o(_al_u617_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u618 (
    .a(_al_u614_o),
    .b(_al_u616_o),
    .c(_al_u617_o),
    .d(M_result2[2]),
    .e(M_result2[1]),
    .o(_al_u618_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u619 (
    .a(_al_u613_o),
    .b(_al_u618_o),
    .c(_al_u572_o),
    .d(M_result2[5]),
    .o(_al_u619_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u620 (
    .a(_al_u588_o),
    .b(_al_u581_o),
    .c(M_result2[3]),
    .d(M_result2[4]),
    .o(_al_u620_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~A*(C*~(D)*~(E)+~(C)*D*E))"),
    .INIT(32'h01000010))
    _al_u621 (
    .a(M_result2[19]),
    .b(M_result2[16]),
    .c(_al_u565_o),
    .d(_al_u481_o),
    .e(_al_u490_o),
    .o(_al_u621_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+~(A)*~(B)*C+A*~(B)*C+~(A)*B*C)"),
    .INIT(8'h7e))
    _al_u622 (
    .a(_al_u427_o),
    .b(_al_u433_o),
    .c(_al_u328_o),
    .o(_al_u622_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    _al_u623 (
    .a(M_result2[15]),
    .b(_al_u586_o),
    .c(M_result2[12]),
    .d(_al_u622_o),
    .e(M_result2[9]),
    .o(_al_u623_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*C*B*~A)"),
    .INIT(16'h0040))
    _al_u624 (
    .a(_al_u545_o),
    .b(_al_u621_o),
    .c(_al_u623_o),
    .d(_al_u510_o),
    .o(_al_u624_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u625 (
    .a(_al_u619_o),
    .b(_al_u620_o),
    .c(_al_u624_o),
    .d(M_result[0]),
    .o(_al_u625_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u626 (
    .a(\NM/n4 [14]),
    .b(_al_u625_o),
    .c(_al_u505_o),
    .o(result[14]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u627 (
    .a(_al_u536_o),
    .b(_al_u507_o),
    .c(M_result2[12]),
    .d(M_result2[7]),
    .o(_al_u627_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*B)*~(D*A))"),
    .INIT(32'h0000153f))
    _al_u628 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[13]),
    .d(M_result2[11]),
    .e(_al_u505_o),
    .o(_al_u628_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u629 (
    .a(_al_u627_o),
    .b(_al_u515_o),
    .c(_al_u628_o),
    .d(M_result2[10]),
    .o(_al_u629_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u630 (
    .a(_al_u629_o),
    .b(_al_u568_o),
    .c(_al_u616_o),
    .d(M_result2[5]),
    .e(M_result[0]),
    .o(_al_u630_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u631 (
    .a(_al_u630_o),
    .b(_al_u588_o),
    .c(_al_u581_o),
    .d(M_result2[3]),
    .e(M_result2[2]),
    .o(_al_u631_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u632 (
    .a(_al_u523_o),
    .b(_al_u542_o),
    .c(M_result2[9]),
    .d(M_result2[6]),
    .o(_al_u632_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u633 (
    .a(_al_u617_o),
    .b(_al_u530_o),
    .c(M_result2[8]),
    .d(M_result2[1]),
    .o(_al_u633_o));
  AL_MAP_LUT4 #(
    .EQN("(C*B*~(D*A))"),
    .INIT(16'h40c0))
    _al_u634 (
    .a(_al_u572_o),
    .b(_al_u632_o),
    .c(_al_u633_o),
    .d(M_result2[4]),
    .o(_al_u634_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u635 (
    .a(\NM/n4 [13]),
    .b(_al_u631_o),
    .c(_al_u634_o),
    .d(_al_u505_o),
    .o(result[13]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u636 (
    .a(_al_u536_o),
    .b(M_result2[9]),
    .o(_al_u636_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u637 (
    .a(_al_u636_o),
    .b(_al_u515_o),
    .c(M_result2[12]),
    .o(_al_u637_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u638 (
    .a(_al_u428_o),
    .b(_al_u465_o),
    .o(_al_u638_o));
  AL_MAP_LUT4 #(
    .EQN("~(~D*~(B)*~((C*~A))+~D*B*~((C*~A))+~(~D)*B*(C*~A)+~D*B*(C*~A))"),
    .INIT(16'hbf10))
    _al_u639 (
    .a(_al_u352_o),
    .b(_al_u638_o),
    .c(_al_u427_o),
    .d(_al_u468_o),
    .o(_al_u639_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u64 (
    .a(n1[26]),
    .b(n1[25]),
    .c(n1[24]),
    .d(n1[23]),
    .o(_al_u64_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*~B*~A)"),
    .INIT(32'h00010000))
    _al_u640 (
    .a(_al_u579_o),
    .b(_al_u639_o),
    .c(_al_u622_o),
    .d(M_result2[9]),
    .e(M_result2[8]),
    .o(_al_u640_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*~C*B*A)"),
    .INIT(32'h00000008))
    _al_u641 (
    .a(_al_u621_o),
    .b(_al_u640_o),
    .c(M_result2[21]),
    .d(_al_u510_o),
    .e(M_result2[20]),
    .o(_al_u641_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u642 (
    .a(_al_u637_o),
    .b(_al_u624_o),
    .c(_al_u641_o),
    .d(M_result2[1]),
    .e(M_result[0]),
    .o(_al_u642_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u643 (
    .a(_al_u642_o),
    .b(_al_u588_o),
    .c(_al_u581_o),
    .d(M_result2[5]),
    .e(M_result2[4]),
    .o(_al_u643_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u644 (
    .a(_al_u542_o),
    .b(M_result2[8]),
    .o(_al_u644_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~(D*C)*~(E*A))"),
    .INIT(32'h01110333))
    _al_u645 (
    .a(_al_u568_o),
    .b(_al_u644_o),
    .c(_al_u530_o),
    .d(M_result2[10]),
    .e(M_result2[7]),
    .o(_al_u645_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*B)*~(D*A))"),
    .INIT(32'h0000153f))
    _al_u646 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[15]),
    .d(M_result2[13]),
    .e(_al_u505_o),
    .o(_al_u646_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*~C)*~(E*B))"),
    .INIT(32'h2022a0aa))
    _al_u647 (
    .a(_al_u646_o),
    .b(_al_u523_o),
    .c(_al_u507_o),
    .d(M_result2[14]),
    .e(M_result2[11]),
    .o(_al_u647_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u648 (
    .a(_al_u647_o),
    .b(_al_u616_o),
    .c(_al_u617_o),
    .d(M_result2[3]),
    .e(M_result2[2]),
    .o(_al_u648_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u649 (
    .a(_al_u645_o),
    .b(_al_u648_o),
    .c(_al_u572_o),
    .d(M_result2[6]),
    .o(_al_u649_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u65 (
    .a(n1[28]),
    .b(n1[27]),
    .o(_al_u65_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u650 (
    .a(\NM/n4 [15]),
    .b(_al_u643_o),
    .c(_al_u649_o),
    .d(_al_u505_o),
    .o(result[15]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u651 (
    .a(_al_u515_o),
    .b(_al_u536_o),
    .c(M_result2[13]),
    .d(M_result2[10]),
    .o(_al_u651_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u652 (
    .a(M_result2[23]),
    .b(M_result2[16]),
    .o(_al_u652_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u653 (
    .a(_al_u511_o),
    .b(_al_u652_o),
    .c(M_result2[14]),
    .d(_al_u505_o),
    .o(_al_u653_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u654 (
    .a(_al_u651_o),
    .b(_al_u653_o),
    .c(_al_u507_o),
    .d(M_result2[15]),
    .o(_al_u654_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u655 (
    .a(_al_u530_o),
    .b(M_result2[11]),
    .o(_al_u655_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*A*~(D*B))"),
    .INIT(16'h020a))
    _al_u656 (
    .a(_al_u654_o),
    .b(_al_u568_o),
    .c(_al_u655_o),
    .d(M_result2[8]),
    .o(_al_u656_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u657 (
    .a(_al_u586_o),
    .b(M_result2[12]),
    .o(_al_u657_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u658 (
    .a(_al_u622_o),
    .b(M_result2[9]),
    .o(_al_u658_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*A)"),
    .INIT(16'h0800))
    _al_u659 (
    .a(_al_u657_o),
    .b(_al_u658_o),
    .c(M_result2[8]),
    .d(M_result2[7]),
    .o(_al_u659_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*A)"),
    .INIT(16'h0008))
    _al_u66 (
    .a(_al_u64_o),
    .b(_al_u65_o),
    .c(n1[30]),
    .d(n1[29]),
    .o(_al_u66_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u660 (
    .a(_al_u571_o),
    .b(_al_u659_o),
    .o(_al_u660_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u661 (
    .a(_al_u572_o),
    .b(_al_u660_o),
    .c(M_result2[7]),
    .d(M_result[0]),
    .o(_al_u661_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u662 (
    .a(_al_u523_o),
    .b(_al_u617_o),
    .c(M_result2[12]),
    .d(M_result2[4]),
    .o(_al_u662_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u663 (
    .a(_al_u616_o),
    .b(_al_u542_o),
    .c(M_result2[3]),
    .d(M_result2[9]),
    .o(_al_u663_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u664 (
    .a(_al_u656_o),
    .b(_al_u661_o),
    .c(_al_u662_o),
    .d(_al_u663_o),
    .o(_al_u664_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u665 (
    .a(_al_u624_o),
    .b(M_result2[2]),
    .o(_al_u665_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u666 (
    .a(_al_u665_o),
    .b(_al_u588_o),
    .c(M_result2[5]),
    .o(_al_u666_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u667 (
    .a(_al_u546_o),
    .b(_al_u640_o),
    .o(_al_u667_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u668 (
    .a(_al_u666_o),
    .b(_al_u667_o),
    .c(_al_u581_o),
    .d(M_result2[6]),
    .e(M_result2[1]),
    .o(_al_u668_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u669 (
    .a(\NM/n4 [16]),
    .b(_al_u664_o),
    .c(_al_u668_o),
    .d(_al_u505_o),
    .o(result[16]));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u67 (
    .a(n1[23]),
    .b(n2[23]),
    .o(_al_u67_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u670 (
    .a(_al_u588_o),
    .b(_al_u581_o),
    .c(M_result2[7]),
    .d(M_result2[6]),
    .o(_al_u670_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u671 (
    .a(_al_u670_o),
    .b(_al_u667_o),
    .c(_al_u624_o),
    .d(M_result2[3]),
    .e(M_result2[2]),
    .o(_al_u671_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u672 (
    .a(_al_u616_o),
    .b(_al_u542_o),
    .c(M_result2[10]),
    .d(M_result2[4]),
    .o(_al_u672_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(D*C)*~(E*A))"),
    .INIT(32'h04440ccc))
    _al_u673 (
    .a(_al_u568_o),
    .b(_al_u672_o),
    .c(_al_u530_o),
    .d(M_result2[12]),
    .e(M_result2[9]),
    .o(_al_u673_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u674 (
    .a(_al_u515_o),
    .b(_al_u507_o),
    .c(M_result2[16]),
    .d(M_result2[14]),
    .o(_al_u674_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*B)*~(D*A))"),
    .INIT(32'h0000153f))
    _al_u675 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[17]),
    .d(M_result2[15]),
    .e(_al_u505_o),
    .o(_al_u675_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u676 (
    .a(_al_u674_o),
    .b(_al_u675_o),
    .c(_al_u536_o),
    .d(M_result2[11]),
    .o(_al_u676_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u677 (
    .a(_al_u523_o),
    .b(_al_u617_o),
    .c(M_result2[13]),
    .d(M_result2[5]),
    .o(_al_u677_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u678 (
    .a(_al_u671_o),
    .b(_al_u673_o),
    .c(_al_u676_o),
    .d(_al_u677_o),
    .o(_al_u678_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u679 (
    .a(M_result2[8]),
    .b(M_result2[7]),
    .o(_al_u679_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C)*~(B)+~A*C*~(B)+~(~A)*C*B+~A*C*B)"),
    .INIT(8'hd1))
    _al_u68 (
    .a(_al_u66_o),
    .b(_al_u67_o),
    .c(n1[22]),
    .o(n87_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u680 (
    .a(_al_u657_o),
    .b(_al_u658_o),
    .c(_al_u679_o),
    .d(M_result2[6]),
    .o(_al_u680_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~D*C*~B*A)"),
    .INIT(32'h00000020))
    _al_u681 (
    .a(_al_u680_o),
    .b(_al_u545_o),
    .c(_al_u621_o),
    .d(_al_u510_o),
    .e(M_result2[15]),
    .o(_al_u681_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u682 (
    .a(_al_u660_o),
    .b(_al_u681_o),
    .c(M_result2[1]),
    .d(M_result[0]),
    .o(_al_u682_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u683 (
    .a(_al_u682_o),
    .b(_al_u572_o),
    .c(M_result2[8]),
    .o(_al_u683_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u684 (
    .a(\NM/n4 [17]),
    .b(_al_u678_o),
    .c(_al_u683_o),
    .d(_al_u505_o),
    .o(result[17]));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u685 (
    .a(_al_u536_o),
    .b(M_result2[13]),
    .o(_al_u685_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u686 (
    .a(_al_u685_o),
    .b(_al_u515_o),
    .c(M_result2[16]),
    .o(_al_u686_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*B)*~(D*A))"),
    .INIT(32'h0000153f))
    _al_u687 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[19]),
    .d(M_result2[17]),
    .e(_al_u505_o),
    .o(_al_u687_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*~C))"),
    .INIT(16'h8088))
    _al_u688 (
    .a(_al_u686_o),
    .b(_al_u687_o),
    .c(_al_u507_o),
    .d(M_result2[18]),
    .o(_al_u688_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u689 (
    .a(_al_u624_o),
    .b(M_result2[5]),
    .o(_al_u689_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u69 (
    .a(_al_u67_o),
    .b(n1[21]),
    .c(n1[20]),
    .o(n89_lutinv));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(D*C)*~(E*B))"),
    .INIT(32'h01110555))
    _al_u690 (
    .a(_al_u689_o),
    .b(_al_u667_o),
    .c(_al_u581_o),
    .d(M_result2[9]),
    .e(M_result2[4]),
    .o(_al_u690_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*~A*~(E@(D*~C)))"),
    .INIT(32'h01001011))
    _al_u691 (
    .a(_al_u579_o),
    .b(M_result2[13]),
    .c(_al_u352_o),
    .d(_al_u427_o),
    .e(_al_u428_o),
    .o(_al_u691_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u692 (
    .a(M_result2[9]),
    .b(M_result2[8]),
    .c(M_result2[7]),
    .d(M_result2[6]),
    .o(_al_u692_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*B*A)"),
    .INIT(32'h00800000))
    _al_u693 (
    .a(_al_u546_o),
    .b(_al_u691_o),
    .c(_al_u692_o),
    .d(_al_u622_o),
    .e(M_result2[5]),
    .o(_al_u693_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u694 (
    .a(_al_u693_o),
    .b(_al_u588_o),
    .c(M_result2[8]),
    .d(M_result2[1]),
    .o(_al_u694_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u695 (
    .a(_al_u616_o),
    .b(_al_u617_o),
    .c(M_result2[7]),
    .d(M_result2[6]),
    .o(_al_u695_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u696 (
    .a(_al_u688_o),
    .b(_al_u690_o),
    .c(_al_u694_o),
    .d(_al_u695_o),
    .o(_al_u696_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u697 (
    .a(_al_u660_o),
    .b(_al_u681_o),
    .c(M_result2[3]),
    .d(M_result2[2]),
    .o(_al_u697_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u698 (
    .a(_al_u523_o),
    .b(_al_u530_o),
    .c(M_result2[15]),
    .d(M_result2[14]),
    .o(_al_u698_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(D*C)*~(E*A))"),
    .INIT(32'h04440ccc))
    _al_u699 (
    .a(_al_u568_o),
    .b(_al_u698_o),
    .c(_al_u542_o),
    .d(M_result2[12]),
    .e(M_result2[11]),
    .o(_al_u699_o));
  AL_MAP_LUT4 #(
    .EQN("(C@A@(D*~B))"),
    .INIT(16'h695a))
    _al_u70 (
    .a(n1[24]),
    .b(n1[23]),
    .c(n2[24]),
    .d(n2[23]),
    .o(_al_u70_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u700 (
    .a(_al_u697_o),
    .b(_al_u699_o),
    .c(_al_u572_o),
    .d(M_result2[10]),
    .o(_al_u700_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u701 (
    .a(\NM/n4 [19]),
    .b(_al_u696_o),
    .c(_al_u700_o),
    .d(_al_u505_o),
    .o(result[19]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u702 (
    .a(_al_u568_o),
    .b(_al_u542_o),
    .c(M_result2[11]),
    .d(M_result2[10]),
    .o(_al_u702_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u703 (
    .a(_al_u693_o),
    .b(_al_u588_o),
    .c(M_result2[7]),
    .d(M_result[0]),
    .o(_al_u703_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*B)*~(D*A))"),
    .INIT(32'h0000153f))
    _al_u704 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[18]),
    .d(M_result2[16]),
    .e(_al_u505_o),
    .o(_al_u704_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*~B))"),
    .INIT(8'h8a))
    _al_u705 (
    .a(_al_u704_o),
    .b(_al_u507_o),
    .c(M_result2[17]),
    .o(_al_u705_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u706 (
    .a(_al_u515_o),
    .b(_al_u536_o),
    .c(M_result2[15]),
    .d(M_result2[12]),
    .o(_al_u706_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u707 (
    .a(_al_u702_o),
    .b(_al_u703_o),
    .c(_al_u705_o),
    .d(_al_u706_o),
    .o(_al_u707_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u708 (
    .a(_al_u624_o),
    .b(M_result2[4]),
    .o(_al_u708_o));
  AL_MAP_LUT3 #(
    .EQN("(~A*~(C*B))"),
    .INIT(8'h15))
    _al_u709 (
    .a(_al_u708_o),
    .b(_al_u667_o),
    .c(M_result2[3]),
    .o(_al_u709_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'hacca))
    _al_u71 (
    .a(n87_lutinv),
    .b(n89_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u71_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(D*A)))"),
    .INIT(16'he0c0))
    _al_u710 (
    .a(_al_u571_o),
    .b(_al_u523_o),
    .c(M_result2[14]),
    .d(M_result2[9]),
    .o(_al_u710_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*B*A*~(E*D))"),
    .INIT(32'h00080808))
    _al_u711 (
    .a(_al_u707_o),
    .b(_al_u709_o),
    .c(_al_u710_o),
    .d(_al_u581_o),
    .e(M_result2[8]),
    .o(_al_u711_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u712 (
    .a(_al_u616_o),
    .b(_al_u617_o),
    .c(M_result2[6]),
    .d(M_result2[5]),
    .o(_al_u712_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u713 (
    .a(_al_u712_o),
    .b(_al_u530_o),
    .c(M_result2[13]),
    .o(_al_u713_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u714 (
    .a(_al_u713_o),
    .b(_al_u660_o),
    .c(_al_u681_o),
    .d(M_result2[2]),
    .e(M_result2[1]),
    .o(_al_u714_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u715 (
    .a(\NM/n4 [18]),
    .b(_al_u711_o),
    .c(_al_u714_o),
    .d(_al_u505_o),
    .o(result[18]));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u716 (
    .a(_al_u536_o),
    .b(_al_u507_o),
    .c(M_result2[19]),
    .d(M_result2[14]),
    .o(_al_u716_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(C*B)*~(D*A))"),
    .INIT(32'h0000153f))
    _al_u717 (
    .a(_al_u511_o),
    .b(M_result2[23]),
    .c(M_result2[20]),
    .d(M_result2[18]),
    .e(_al_u505_o),
    .o(_al_u717_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u718 (
    .a(_al_u716_o),
    .b(_al_u515_o),
    .c(_al_u717_o),
    .d(M_result2[17]),
    .o(_al_u718_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u719 (
    .a(_al_u718_o),
    .b(_al_u624_o),
    .c(M_result2[6]),
    .o(_al_u719_o));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(C)*~((D*~B))+A*~(C)*~((D*~B))+A*C*~((D*~B))+A*~(C)*(D*~B))"),
    .INIT(16'h8eaf))
    _al_u72 (
    .a(n1[24]),
    .b(n1[23]),
    .c(n2[24]),
    .d(n2[23]),
    .o(\ADD01/ADD01/c1_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u720 (
    .a(_al_u545_o),
    .b(_al_u510_o),
    .c(_al_u535_o),
    .d(_al_u587_o),
    .o(_al_u720_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u721 (
    .a(_al_u692_o),
    .b(_al_u622_o),
    .o(_al_u721_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u722 (
    .a(_al_u721_o),
    .b(M_result2[12]),
    .o(_al_u722_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u723 (
    .a(M_result2[5]),
    .b(M_result2[4]),
    .o(_al_u723_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u724 (
    .a(_al_u720_o),
    .b(_al_u722_o),
    .c(_al_u723_o),
    .d(M_result2[3]),
    .o(_al_u724_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u725 (
    .a(_al_u724_o),
    .b(_al_u523_o),
    .c(M_result2[16]),
    .d(M_result[0]),
    .o(_al_u725_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E*C)*~(D*B))"),
    .INIT(32'h020a22aa))
    _al_u726 (
    .a(_al_u725_o),
    .b(_al_u568_o),
    .c(_al_u542_o),
    .d(M_result2[12]),
    .e(M_result2[13]),
    .o(_al_u726_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u727 (
    .a(_al_u667_o),
    .b(_al_u588_o),
    .c(M_result2[9]),
    .d(M_result2[5]),
    .o(_al_u727_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u728 (
    .a(_al_u693_o),
    .b(_al_u581_o),
    .c(M_result2[10]),
    .d(M_result2[2]),
    .o(_al_u728_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u729 (
    .a(_al_u719_o),
    .b(_al_u726_o),
    .c(_al_u727_o),
    .d(_al_u728_o),
    .o(_al_u729_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+~(A)*~(B)*C*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+A*B*~(C)*D*~(E)+~(A)*B*C*D*~(E)+A*B*C*D*~(E)+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*B*C*D*E)"),
    .INIT(32'h80ecc8fe))
    _al_u73 (
    .a(\ADD01/ADD01/c1_lutinv ),
    .b(n1[26]),
    .c(n1[25]),
    .d(n2[26]),
    .e(n2[25]),
    .o(\ADD01/ctemp_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u730 (
    .a(_al_u572_o),
    .b(_al_u681_o),
    .c(M_result2[11]),
    .d(M_result2[3]),
    .o(_al_u730_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u731 (
    .a(_al_u616_o),
    .b(_al_u530_o),
    .c(M_result2[15]),
    .d(M_result2[7]),
    .o(_al_u731_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u732 (
    .a(_al_u731_o),
    .b(_al_u617_o),
    .c(M_result2[8]),
    .o(_al_u732_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u733 (
    .a(_al_u730_o),
    .b(_al_u732_o),
    .c(_al_u660_o),
    .d(M_result2[4]),
    .o(_al_u733_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u734 (
    .a(\NM/n4 [20]),
    .b(_al_u729_o),
    .c(_al_u733_o),
    .d(_al_u505_o),
    .o(result[20]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u735 (
    .a(_al_u523_o),
    .b(_al_u616_o),
    .c(M_result2[17]),
    .d(M_result2[8]),
    .o(_al_u735_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u736 (
    .a(_al_u735_o),
    .b(_al_u724_o),
    .c(_al_u617_o),
    .d(M_result2[9]),
    .e(M_result2[1]),
    .o(_al_u736_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*~B)*~(D*A))"),
    .INIT(16'h45cf))
    _al_u737 (
    .a(_al_u536_o),
    .b(_al_u507_o),
    .c(M_result2[20]),
    .d(M_result2[15]),
    .o(_al_u737_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(A*~(~B*~(D*~C))))"),
    .INIT(32'h00007577))
    _al_u738 (
    .a(M_result2[21]),
    .b(M_result2[23]),
    .c(_al_u510_o),
    .d(M_result2[19]),
    .e(_al_u505_o),
    .o(_al_u738_o));
  AL_MAP_LUT4 #(
    .EQN("(C*A*~(D*B))"),
    .INIT(16'h20a0))
    _al_u739 (
    .a(_al_u737_o),
    .b(_al_u515_o),
    .c(_al_u738_o),
    .d(M_result2[18]),
    .o(_al_u739_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u74 (
    .a(n1[28]),
    .b(n2[28]),
    .o(\ADD01/ADD02/g1 ));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u740 (
    .a(_al_u736_o),
    .b(_al_u739_o),
    .c(_al_u693_o),
    .d(M_result2[3]),
    .o(_al_u740_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~B*~(C*A)))"),
    .INIT(16'hec00))
    _al_u741 (
    .a(_al_u571_o),
    .b(_al_u542_o),
    .c(M_result2[12]),
    .d(M_result2[14]),
    .o(_al_u741_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u742 (
    .a(_al_u588_o),
    .b(_al_u581_o),
    .c(M_result2[11]),
    .d(M_result2[10]),
    .o(_al_u742_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u743 (
    .a(_al_u667_o),
    .b(_al_u624_o),
    .c(M_result2[7]),
    .d(M_result2[6]),
    .o(_al_u743_o));
  AL_MAP_LUT4 #(
    .EQN("(D*C*~B*A)"),
    .INIT(16'h2000))
    _al_u744 (
    .a(_al_u740_o),
    .b(_al_u741_o),
    .c(_al_u742_o),
    .d(_al_u743_o),
    .o(_al_u744_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~A*(D@C))"),
    .INIT(16'h0110))
    _al_u745 (
    .a(M_result2[5]),
    .b(M_result2[4]),
    .c(_al_u456_o),
    .d(_al_u457_o),
    .o(_al_u745_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'h00080000))
    _al_u746 (
    .a(_al_u692_o),
    .b(_al_u745_o),
    .c(M_result2[12]),
    .d(_al_u622_o),
    .e(M_result2[2]),
    .o(_al_u746_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u747 (
    .a(_al_u720_o),
    .b(_al_u746_o),
    .o(_al_u747_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u748 (
    .a(_al_u530_o),
    .b(M_result2[16]),
    .o(_al_u748_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~(E*B)*~(D*A))"),
    .INIT(32'h0103050f))
    _al_u749 (
    .a(_al_u568_o),
    .b(_al_u747_o),
    .c(_al_u748_o),
    .d(M_result2[13]),
    .e(M_result[0]),
    .o(_al_u749_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+~(A)*~(B)*~(C)*D*~(E)+A*~(B)*~(C)*D*~(E)+~(A)*B*~(C)*D*~(E)+~(A)*~(B)*C*D*~(E)+A*~(B)*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*~(B)*C*~(D)*E+~(A)*~(B)*~(C)*D*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+~(A)*~(B)*C*D*E+A*~(B)*C*D*E+~(A)*B*C*D*E)"),
    .INIT(32'h7f133701))
    _al_u75 (
    .a(\ADD01/ADD02/g1 ),
    .b(n1[30]),
    .c(n1[29]),
    .d(n2[30]),
    .e(n2[29]),
    .o(_al_u75_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C*B))"),
    .INIT(8'h2a))
    _al_u750 (
    .a(_al_u749_o),
    .b(_al_u660_o),
    .c(M_result2[5]),
    .o(_al_u750_o));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D*C))"),
    .INIT(16'h0888))
    _al_u751 (
    .a(_al_u744_o),
    .b(_al_u750_o),
    .c(_al_u681_o),
    .d(M_result2[4]),
    .o(_al_u751_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*~A))"),
    .INIT(8'h23))
    _al_u752 (
    .a(\NM/n4 [21]),
    .b(_al_u751_o),
    .c(_al_u505_o),
    .o(result[21]));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u753 (
    .a(_al_u660_o),
    .b(_al_u681_o),
    .c(M_result2[6]),
    .d(M_result2[5]),
    .o(_al_u753_o));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*C*~(D)+~(A)*B*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'he2e0))
    _al_u754 (
    .a(M_result2[21]),
    .b(M_result2[23]),
    .c(M_result2[22]),
    .d(M_result2[20]),
    .o(_al_u754_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~B*~(C*A))"),
    .INIT(16'h0013))
    _al_u755 (
    .a(_al_u515_o),
    .b(_al_u754_o),
    .c(M_result2[19]),
    .d(_al_u505_o),
    .o(_al_u755_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*A)"),
    .INIT(8'h20))
    _al_u756 (
    .a(_al_u522_o),
    .b(_al_u535_o),
    .c(M_result2[16]),
    .o(_al_u756_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D*C)*~(E*B))"),
    .INIT(32'h02220aaa))
    _al_u757 (
    .a(_al_u755_o),
    .b(_al_u616_o),
    .c(_al_u756_o),
    .d(M_result2[17]),
    .e(M_result2[9]),
    .o(_al_u757_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D*B)*~(C*A))"),
    .INIT(16'h135f))
    _al_u758 (
    .a(_al_u724_o),
    .b(_al_u747_o),
    .c(M_result2[2]),
    .d(M_result2[1]),
    .o(_al_u758_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u759 (
    .a(_al_u617_o),
    .b(_al_u542_o),
    .c(M_result2[15]),
    .d(M_result2[10]),
    .o(_al_u759_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u76 (
    .a(n1[28]),
    .b(n2[28]),
    .o(\ADD01/ADD02/p1_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(D*C*B*A)"),
    .INIT(16'h8000))
    _al_u760 (
    .a(_al_u753_o),
    .b(_al_u757_o),
    .c(_al_u758_o),
    .d(_al_u759_o),
    .o(_al_u760_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u761 (
    .a(_al_u578_o),
    .b(_al_u579_o),
    .c(_al_u639_o),
    .o(_al_u761_o));
  AL_MAP_LUT4 #(
    .EQN("(B*(~(A)*C*~(D)+A*~(C)*D))"),
    .INIT(16'h0840))
    _al_u762 (
    .a(_al_u427_o),
    .b(M_result2[1]),
    .c(_al_u449_o),
    .d(_al_u452_o),
    .o(_al_u762_o));
  AL_MAP_LUT5 #(
    .EQN("(~(B)*~((D*A))*~((E@C))+B*~((D*A))*~((E@C))+B*(D*A)*~((E@C))+~(B)*~((D*A))*(E@C)+~(B)*(D*A)*(E@C)+B*(D*A)*(E@C))"),
    .INIT(32'hdbf3bd3f))
    _al_u763 (
    .a(_al_u427_o),
    .b(_al_u457_o),
    .c(_al_u195_o),
    .d(_al_u339_o),
    .e(_al_u255_o),
    .o(_al_u763_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u764 (
    .a(_al_u762_o),
    .b(_al_u763_o),
    .o(_al_u764_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u765 (
    .a(_al_u577_o),
    .b(_al_u761_o),
    .c(_al_u721_o),
    .d(_al_u764_o),
    .e(M_result[0]),
    .o(_al_u765_o));
  AL_MAP_LUT3 #(
    .EQN("(~B*~(C*A))"),
    .INIT(8'h13))
    _al_u766 (
    .a(_al_u581_o),
    .b(_al_u765_o),
    .c(M_result2[12]),
    .o(_al_u766_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(~B*~(D*A)))"),
    .INIT(16'he0c0))
    _al_u767 (
    .a(_al_u540_o),
    .b(_al_u523_o),
    .c(M_result2[18]),
    .d(M_result2[17]),
    .o(_al_u767_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*A*~(D*C))"),
    .INIT(16'h0222))
    _al_u768 (
    .a(_al_u766_o),
    .b(_al_u767_o),
    .c(_al_u588_o),
    .d(M_result2[11]),
    .o(_al_u768_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(~A*~(C*B)))"),
    .INIT(16'hea00))
    _al_u769 (
    .a(_al_u568_o),
    .b(_al_u571_o),
    .c(M_result2[13]),
    .d(M_result2[14]),
    .o(_al_u769_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(E@C)*~(D@B))"),
    .INIT(32'h80200802))
    _al_u77 (
    .a(\ADD01/ADD02/p1_lutinv ),
    .b(n1[30]),
    .c(n1[29]),
    .d(n2[30]),
    .e(n2[29]),
    .o(\ADD01/ADD02/n17 ));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*A))"),
    .INIT(16'h153f))
    _al_u770 (
    .a(_al_u693_o),
    .b(_al_u624_o),
    .c(M_result2[8]),
    .d(M_result2[4]),
    .o(_al_u770_o));
  AL_MAP_LUT5 #(
    .EQN("(C*~B*A*~(E*D))"),
    .INIT(32'h00202020))
    _al_u771 (
    .a(_al_u768_o),
    .b(_al_u769_o),
    .c(_al_u770_o),
    .d(_al_u667_o),
    .e(M_result2[7]),
    .o(_al_u771_o));
  AL_MAP_LUT4 #(
    .EQN("(~(C*B)*~(D*~A))"),
    .INIT(16'h2a3f))
    _al_u772 (
    .a(\NM/n4 [22]),
    .b(_al_u760_o),
    .c(_al_u771_o),
    .d(_al_u505_o),
    .o(result[22]));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~B*~A)"),
    .INIT(16'h0001))
    _al_u773 (
    .a(_al_u578_o),
    .b(_al_u579_o),
    .c(_al_u639_o),
    .d(_al_u762_o),
    .o(_al_u773_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~(B@A))"),
    .INIT(8'h90))
    _al_u774 (
    .a(_al_u427_o),
    .b(_al_u454_o),
    .c(M_result[0]),
    .o(_al_u774_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*B*~(~A*~(E*C)))"),
    .INIT(32'h00c80088))
    _al_u775 (
    .a(_al_u764_o),
    .b(_al_u692_o),
    .c(_al_u745_o),
    .d(_al_u622_o),
    .e(_al_u774_o),
    .o(_al_u775_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u776 (
    .a(_al_u773_o),
    .b(_al_u577_o),
    .c(_al_u775_o),
    .o(_al_u776_o));
  AL_MAP_LUT3 #(
    .EQN("(C*~B*~A)"),
    .INIT(8'h10))
    _al_u777 (
    .a(_al_u578_o),
    .b(M_result2[15]),
    .c(M_result2[14]),
    .o(_al_u777_o));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(~B*~(~D*A)))"),
    .INIT(16'h0c0e))
    _al_u778 (
    .a(_al_u615_o),
    .b(_al_u777_o),
    .c(_al_u535_o),
    .d(M_result2[17]),
    .o(_al_u778_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(C*~B*(E@D)))"),
    .INIT(32'haa8a8aaa))
    _al_u779 (
    .a(_al_u507_o),
    .b(_al_u510_o),
    .c(M_result2[20]),
    .d(_al_u521_o),
    .e(_al_u499_o),
    .o(_al_u779_o));
  AL_MAP_LUT5 #(
    .EQN("(B*~(C*(A*~(D)*~(E)+~(A)*D*~(E)+A*D*~(E)+A*D*E)))"),
    .INIT(32'h4ccc0c4c))
    _al_u78 (
    .a(\ADD01/ctemp_lutinv ),
    .b(_al_u75_o),
    .c(\ADD01/ADD02/n17 ),
    .d(n1[27]),
    .e(n2[27]),
    .o(_al_u78_o));
  AL_MAP_LUT5 #(
    .EQN("(D*~B*~A*~(E*C))"),
    .INIT(32'h01001100))
    _al_u780 (
    .a(_al_u641_o),
    .b(_al_u776_o),
    .c(_al_u778_o),
    .d(_al_u779_o),
    .e(_al_u522_o),
    .o(_al_u780_o));
  AL_MAP_LUT5 #(
    .EQN("(~C*~A*~(B*~(~E*~D)))"),
    .INIT(32'h01010105))
    _al_u781 (
    .a(_al_u542_o),
    .b(_al_u720_o),
    .c(_al_u530_o),
    .d(_al_u746_o),
    .e(M_result2[12]),
    .o(_al_u781_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u782 (
    .a(_al_u78_o),
    .b(n1[23]),
    .c(n2[23]),
    .o(E[0]));
  AL_MAP_LUT5 #(
    .EQN("~(E@(~D*~C*B*A))"),
    .INIT(32'h0008fff7))
    _al_u783 (
    .a(_al_u780_o),
    .b(_al_u781_o),
    .c(_al_u681_o),
    .d(_al_u505_o),
    .e(E[0]),
    .o(\ADD03/ADD01/p0_neg ));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u784 (
    .a(_al_u505_o),
    .b(E[0]),
    .o(_al_u784_o));
  AL_MAP_LUT4 #(
    .EQN("(C*~(D*~B*A))"),
    .INIT(16'hd0f0))
    _al_u785 (
    .a(_al_u781_o),
    .b(_al_u681_o),
    .c(_al_u784_o),
    .d(_al_u780_o),
    .o(_al_u785_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*~(~A*~(D*~C)))"),
    .INIT(16'h2322))
    _al_u786 (
    .a(_al_u545_o),
    .b(_al_u510_o),
    .c(_al_u535_o),
    .d(_al_u578_o),
    .o(_al_u786_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u787 (
    .a(_al_u786_o),
    .b(_al_u577_o),
    .c(_al_u580_o),
    .d(_al_u639_o),
    .o(_al_u787_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*B*~A)"),
    .INIT(16'h0400))
    _al_u788 (
    .a(M_result2[21]),
    .b(_al_u692_o),
    .c(_al_u622_o),
    .d(M_result2[5]),
    .o(_al_u788_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*D*~C*B*A)"),
    .INIT(32'h00000800))
    _al_u789 (
    .a(_al_u567_o),
    .b(_al_u788_o),
    .c(_al_u510_o),
    .d(_al_u691_o),
    .e(_al_u529_o),
    .o(_al_u789_o));
  AL_MAP_LUT3 #(
    .EQN("~(C@B@A)"),
    .INIT(8'h69))
    _al_u79 (
    .a(\ADD01/ADD01/c1_lutinv ),
    .b(n1[25]),
    .c(n2[25]),
    .o(_al_u79_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(E*~D*~C*B))"),
    .INIT(32'h55515555))
    _al_u790 (
    .a(_al_u640_o),
    .b(_al_u657_o),
    .c(M_result2[15]),
    .d(_al_u622_o),
    .e(M_result2[9]),
    .o(_al_u790_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*B*~(~A*~(E*C)))"),
    .INIT(32'h00c80088))
    _al_u791 (
    .a(_al_u764_o),
    .b(_al_u692_o),
    .c(_al_u745_o),
    .d(_al_u622_o),
    .e(_al_u774_o),
    .o(_al_u791_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u792 (
    .a(_al_u577_o),
    .b(_al_u791_o),
    .c(_al_u761_o),
    .o(_al_u792_o));
  AL_MAP_LUT5 #(
    .EQN("(~B*A*~(C*~(~E*D)))"),
    .INIT(32'h02022202))
    _al_u793 (
    .a(_al_u787_o),
    .b(_al_u789_o),
    .c(_al_u546_o),
    .d(_al_u790_o),
    .e(_al_u792_o),
    .o(_al_u793_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u794 (
    .a(_al_u78_o),
    .b(n1[24]),
    .c(n2[24]),
    .o(E[1]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'h78))
    _al_u795 (
    .a(_al_u505_o),
    .b(E[0]),
    .c(E[1]),
    .o(_al_u795_o));
  AL_MAP_LUT4 #(
    .EQN("(C@A@(~D*~B))"),
    .INIT(16'h5a69))
    _al_u796 (
    .a(_al_u785_o),
    .b(_al_u793_o),
    .c(_al_u795_o),
    .d(_al_u505_o),
    .o(result[24]));
  AL_MAP_LUT5 #(
    .EQN("(~B*~A*(C*~(D)*~(E)+~(C)*D*E))"),
    .INIT(32'h01000010))
    _al_u797 (
    .a(M_result2[21]),
    .b(_al_u529_o),
    .c(_al_u565_o),
    .d(_al_u481_o),
    .e(_al_u490_o),
    .o(_al_u797_o));
  AL_MAP_LUT5 #(
    .EQN("(~A*~(~D*B*~(E*~C)))"),
    .INIT(32'h55155511))
    _al_u798 (
    .a(_al_u617_o),
    .b(_al_u797_o),
    .c(_al_u615_o),
    .d(_al_u510_o),
    .e(_al_u790_o),
    .o(_al_u798_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*C*~B*A)"),
    .INIT(32'h00200000))
    _al_u799 (
    .a(_al_u692_o),
    .b(M_result2[12]),
    .c(_al_u723_o),
    .d(_al_u622_o),
    .e(_al_u763_o),
    .o(_al_u799_o));
  AL_MAP_LUT3 #(
    .EQN("(A*~(C@B))"),
    .INIT(8'h82))
    _al_u80 (
    .a(_al_u67_o),
    .b(n1[24]),
    .c(n2[24]),
    .o(\ADD01/ADD01/n3 ));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*~A)"),
    .INIT(32'h00040000))
    _al_u800 (
    .a(_al_u545_o),
    .b(_al_u587_o),
    .c(_al_u510_o),
    .d(_al_u535_o),
    .e(_al_u799_o),
    .o(_al_u800_o));
  AL_MAP_LUT4 #(
    .EQN("(~A*~(D*C*B))"),
    .INIT(16'h1555))
    _al_u801 (
    .a(_al_u800_o),
    .b(_al_u577_o),
    .c(_al_u775_o),
    .d(_al_u761_o),
    .o(_al_u801_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u802 (
    .a(_al_u505_o),
    .b(E[0]),
    .c(E[1]),
    .o(_al_u802_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u803 (
    .a(_al_u78_o),
    .b(n1[25]),
    .c(n2[25]),
    .o(E[2]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u804 (
    .a(_al_u802_o),
    .b(E[2]),
    .o(_al_u804_o));
  AL_MAP_LUT4 #(
    .EQN("(~(~C*B)*~(D*A))"),
    .INIT(16'h51f3))
    _al_u805 (
    .a(_al_u720_o),
    .b(_al_u522_o),
    .c(_al_u621_o),
    .d(_al_u799_o),
    .o(_al_u805_o));
  AL_MAP_LUT5 #(
    .EQN("~(C@(~D*~(E*B*A)))"),
    .INIT(32'h0f780ff0))
    _al_u806 (
    .a(_al_u798_o),
    .b(_al_u801_o),
    .c(_al_u804_o),
    .d(_al_u505_o),
    .e(_al_u805_o),
    .o(_al_u806_o));
  AL_MAP_LUT5 #(
    .EQN("(A@(~(B)*~((~D*~C))*~(E)+~(B)*~((~D*~C))*E+B*~((~D*~C))*E+~(B)*(~D*~C)*E))"),
    .INIT(32'h5559999a))
    _al_u807 (
    .a(_al_u806_o),
    .b(_al_u785_o),
    .c(_al_u793_o),
    .d(_al_u505_o),
    .e(E[1]),
    .o(result[25]));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~((~C*~B))*~(D)+~(A)*~((~C*~B))*D+A*~((~C*~B))*D+~(A)*(~C*~B)*D)"),
    .INIT(16'hfd54))
    _al_u808 (
    .a(_al_u785_o),
    .b(_al_u793_o),
    .c(_al_u505_o),
    .d(E[1]),
    .o(_al_u808_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u809 (
    .a(_al_u790_o),
    .b(_al_u545_o),
    .c(_al_u510_o),
    .o(_al_u809_o));
  AL_MAP_LUT3 #(
    .EQN("(B@(~C*A))"),
    .INIT(8'hc6))
    _al_u81 (
    .a(_al_u78_o),
    .b(_al_u79_o),
    .c(\ADD01/ADD01/n3 ),
    .o(exp_diff[2]));
  AL_MAP_LUT4 #(
    .EQN("(D*~C*~B*~A)"),
    .INIT(16'h0100))
    _al_u810 (
    .a(M_result2[21]),
    .b(_al_u510_o),
    .c(_al_u529_o),
    .d(_al_u615_o),
    .o(_al_u810_o));
  AL_MAP_LUT3 #(
    .EQN("(~C*~B*~A)"),
    .INIT(8'h01))
    _al_u811 (
    .a(_al_u809_o),
    .b(_al_u607_o),
    .c(_al_u810_o),
    .o(_al_u811_o));
  AL_MAP_LUT4 #(
    .EQN("(D*~(C*B*A))"),
    .INIT(16'h7f00))
    _al_u812 (
    .a(_al_u577_o),
    .b(_al_u775_o),
    .c(_al_u761_o),
    .d(_al_u805_o),
    .o(_al_u812_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*A)"),
    .INIT(8'h80))
    _al_u813 (
    .a(_al_u811_o),
    .b(_al_u812_o),
    .c(_al_u804_o),
    .o(_al_u813_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*~(B*A))"),
    .INIT(16'h0007))
    _al_u814 (
    .a(_al_u811_o),
    .b(_al_u812_o),
    .c(_al_u505_o),
    .d(E[2]),
    .o(_al_u814_o));
  AL_MAP_LUT5 #(
    .EQN("(E*~D*~C*B*A)"),
    .INIT(32'h00080000))
    _al_u815 (
    .a(_al_u541_o),
    .b(_al_u657_o),
    .c(M_result2[15]),
    .d(M_result2[16]),
    .e(M_result2[11]),
    .o(_al_u815_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*B*~(~C*~A))"),
    .INIT(16'h00c8))
    _al_u816 (
    .a(_al_u815_o),
    .b(_al_u797_o),
    .c(_al_u615_o),
    .d(_al_u510_o),
    .o(_al_u816_o));
  AL_MAP_LUT3 #(
    .EQN("(C*B*~A)"),
    .INIT(8'h40))
    _al_u817 (
    .a(_al_u790_o),
    .b(_al_u522_o),
    .c(_al_u621_o),
    .o(_al_u817_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*~C*B*~A)"),
    .INIT(16'h0004))
    _al_u818 (
    .a(_al_u545_o),
    .b(_al_u621_o),
    .c(_al_u510_o),
    .d(_al_u691_o),
    .o(_al_u818_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u819 (
    .a(_al_u78_o),
    .b(n1[26]),
    .c(n2[26]),
    .o(E[3]));
  AL_MAP_LUT5 #(
    .EQN("(D@B@(A*~(C)*~(E)+~(A)*C*~(E)+A*C*~(E)+A*C*E))"),
    .INIT(32'h936cc936))
    _al_u82 (
    .a(\ADD01/ADD01/c1_lutinv ),
    .b(n1[26]),
    .c(n1[25]),
    .d(n2[26]),
    .e(n2[25]),
    .o(\C023/outtemp [3]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'h78))
    _al_u820 (
    .a(_al_u802_o),
    .b(E[2]),
    .c(E[3]),
    .o(_al_u820_o));
  AL_MAP_LUT5 #(
    .EQN("~(D@(~E*~(~C*~B*~A)))"),
    .INIT(32'h00fffe01))
    _al_u821 (
    .a(_al_u816_o),
    .b(_al_u817_o),
    .c(_al_u818_o),
    .d(_al_u820_o),
    .e(_al_u505_o),
    .o(_al_u821_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(~C*~(~B*~A)))"),
    .INIT(16'hf10e))
    _al_u822 (
    .a(_al_u808_o),
    .b(_al_u813_o),
    .c(_al_u814_o),
    .d(_al_u821_o),
    .o(result[26]));
  AL_MAP_LUT4 #(
    .EQN("(~C*~(D*~B*A))"),
    .INIT(16'h0d0f))
    _al_u823 (
    .a(_al_u805_o),
    .b(_al_u792_o),
    .c(_al_u505_o),
    .d(_al_u798_o),
    .o(_al_u823_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*A)"),
    .INIT(4'h2))
    _al_u824 (
    .a(_al_u818_o),
    .b(_al_u505_o),
    .o(_al_u824_o));
  AL_MAP_LUT5 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)*~(E)+A*~(B)*~(C)*~(D)*~(E)+~(A)*B*~(C)*~(D)*~(E)+A*B*~(C)*~(D)*~(E)+A*~(B)*C*~(D)*~(E)+~(A)*B*C*~(D)*~(E)+A*B*C*~(D)*~(E)+~(A)*B*~(C)*D*~(E)+A*B*~(C)*D*~(E)+A*B*C*D*~(E)+~(A)*~(B)*~(C)*~(D)*E+A*~(B)*~(C)*~(D)*E+~(A)*B*~(C)*~(D)*E+A*B*~(C)*~(D)*E+A*~(B)*C*~(D)*E+~(A)*B*C*~(D)*E+A*B*C*~(D)*E+A*~(B)*~(C)*D*E+~(A)*B*~(C)*D*E+A*B*~(C)*D*E+A*~(B)*C*D*E+A*B*C*D*E)"),
    .INIT(32'haeef8cef))
    _al_u825 (
    .a(_al_u823_o),
    .b(_al_u824_o),
    .c(_al_u804_o),
    .d(_al_u820_o),
    .e(_al_u812_o),
    .o(_al_u825_o));
  AL_MAP_LUT4 #(
    .EQN("(~D*A*~(~C*~B))"),
    .INIT(16'h00a8))
    _al_u826 (
    .a(_al_u546_o),
    .b(_al_u659_o),
    .c(_al_u680_o),
    .d(M_result2[15]),
    .o(_al_u826_o));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u827 (
    .a(_al_u505_o),
    .b(E[0]),
    .c(E[1]),
    .d(E[2]),
    .e(E[3]),
    .o(_al_u827_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u828 (
    .a(_al_u78_o),
    .b(n1[27]),
    .c(n2[27]),
    .o(E[4]));
  AL_MAP_LUT2 #(
    .EQN("(B@A)"),
    .INIT(4'h6))
    _al_u829 (
    .a(_al_u827_o),
    .b(E[4]),
    .o(_al_u829_o));
  AL_MAP_LUT4 #(
    .EQN("(~(D@B)*~(C@A))"),
    .INIT(16'h8421))
    _al_u83 (
    .a(n1[25]),
    .b(n1[24]),
    .c(n2[25]),
    .d(n2[24]),
    .o(\ADD01/ADD01/n7 ));
  AL_MAP_LUT5 #(
    .EQN("~(C@(~D*~(E*~B*~A)))"),
    .INIT(32'h0fe10ff0))
    _al_u830 (
    .a(_al_u826_o),
    .b(_al_u789_o),
    .c(_al_u829_o),
    .d(_al_u505_o),
    .e(_al_u801_o),
    .o(_al_u830_o));
  AL_MAP_LUT5 #(
    .EQN("~(C@(B*~(E*D*A)))"),
    .INIT(32'h4bc3c3c3))
    _al_u831 (
    .a(_al_u808_o),
    .b(_al_u825_o),
    .c(_al_u830_o),
    .d(_al_u806_o),
    .e(_al_u821_o),
    .o(result[27]));
  AL_MAP_LUT5 #(
    .EQN("(A*~(D@(~E*~(C*B))))"),
    .INIT(32'h00aa2a80))
    _al_u832 (
    .a(_al_u821_o),
    .b(_al_u811_o),
    .c(_al_u812_o),
    .d(_al_u804_o),
    .e(_al_u505_o),
    .o(_al_u832_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u833 (
    .a(_al_u505_o),
    .b(_al_u793_o),
    .o(_al_u833_o));
  AL_MAP_LUT5 #(
    .EQN("(A*~(B*(~(C)*~(D)*~(E)+~(C)*~(D)*E+C*~(D)*E+~(C)*D*E)))"),
    .INIT(32'ha222aaa2))
    _al_u834 (
    .a(_al_u825_o),
    .b(_al_u832_o),
    .c(_al_u833_o),
    .d(_al_u785_o),
    .e(_al_u795_o),
    .o(_al_u834_o));
  AL_MAP_LUT5 #(
    .EQN("(~E*~(~D*~C*B*~A))"),
    .INIT(32'h0000fffb))
    _al_u835 (
    .a(_al_u660_o),
    .b(_al_u801_o),
    .c(_al_u693_o),
    .d(_al_u681_o),
    .e(_al_u505_o),
    .o(_al_u835_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u836 (
    .a(_al_u78_o),
    .b(n1[28]),
    .c(n2[28]),
    .o(E[5]));
  AL_MAP_LUT3 #(
    .EQN("(C@(B*A))"),
    .INIT(8'h78))
    _al_u837 (
    .a(_al_u827_o),
    .b(E[4]),
    .c(E[5]),
    .o(_al_u837_o));
  AL_MAP_LUT4 #(
    .EQN("(D@(A*~(B)*~(C)+~(A)*B*~(C)+A*B*~(C)+A*B*C))"),
    .INIT(16'h718e))
    _al_u838 (
    .a(_al_u834_o),
    .b(_al_u835_o),
    .c(_al_u829_o),
    .d(_al_u837_o),
    .o(result[28]));
  AL_MAP_LUT5 #(
    .EQN("(C*~(B*~(E*D*A)))"),
    .INIT(32'hb0303030))
    _al_u839 (
    .a(_al_u808_o),
    .b(_al_u825_o),
    .c(_al_u830_o),
    .d(_al_u806_o),
    .e(_al_u821_o),
    .o(_al_u839_o));
  AL_MAP_LUT4 #(
    .EQN("~(B@(A*~(D*C)))"),
    .INIT(16'h3999))
    _al_u84 (
    .a(_al_u78_o),
    .b(\C023/outtemp [3]),
    .c(\ADD01/ADD01/n7 ),
    .d(_al_u67_o),
    .o(exp_diff[3]));
  AL_MAP_LUT2 #(
    .EQN("(B*~A)"),
    .INIT(4'h4))
    _al_u840 (
    .a(_al_u835_o),
    .b(_al_u829_o),
    .o(_al_u840_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u841 (
    .a(_al_u78_o),
    .b(n1[29]),
    .c(n2[29]),
    .o(E[6]));
  AL_MAP_LUT5 #(
    .EQN("(E*D*C*B*A)"),
    .INIT(32'h80000000))
    _al_u842 (
    .a(_al_u802_o),
    .b(E[2]),
    .c(E[3]),
    .d(E[4]),
    .e(E[5]),
    .o(_al_u842_o));
  AL_MAP_LUT2 #(
    .EQN("(B*A)"),
    .INIT(4'h8))
    _al_u843 (
    .a(E[6]),
    .b(_al_u842_o),
    .o(_al_u843_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u844 (
    .a(E[5]),
    .b(E[6]),
    .o(_al_u844_o));
  AL_MAP_LUT2 #(
    .EQN("(~B*~A)"),
    .INIT(4'h1))
    _al_u845 (
    .a(n1[30]),
    .b(n2[30]),
    .o(_al_u845_o));
  AL_MAP_LUT5 #(
    .EQN("(E@(~C*~(D*~B*~A)))"),
    .INIT(32'hf1f00e0f))
    _al_u846 (
    .a(_al_u839_o),
    .b(_al_u840_o),
    .c(_al_u843_o),
    .d(_al_u844_o),
    .e(_al_u845_o),
    .o(result[30]));
  AL_MAP_LUT5 #(
    .EQN("~(E@(~C*~(D)*~((~B*~A))+~C*D*~((~B*~A))+~(~C)*D*(~B*~A)+~C*D*(~B*~A)))"),
    .INIT(32'h1f0ee0f1))
    _al_u847 (
    .a(_al_u839_o),
    .b(_al_u840_o),
    .c(_al_u842_o),
    .d(_al_u837_o),
    .e(E[6]),
    .o(result[29]));
  AL_MAP_LUT4 #(
    .EQN("(B*A*~(D@C))"),
    .INIT(16'h8008))
    _al_u85 (
    .a(\ADD01/ADD01/n7 ),
    .b(_al_u67_o),
    .c(n1[26]),
    .d(n2[26]),
    .o(\ADD01/ADD01/n20 ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(C)*~((~D*B))+~(A)*C*~((~D*B))+A*C*~((~D*B))+~(A)*C*(~D*B))"),
    .INIT(16'hf571))
    _al_u86 (
    .a(n1[28]),
    .b(n1[27]),
    .c(n2[28]),
    .d(n2[27]),
    .o(_al_u86_o));
  AL_MAP_LUT4 #(
    .EQN("(B*~A*~(~D*C))"),
    .INIT(16'h4404))
    _al_u87 (
    .a(\ADD01/ADD01/n20 ),
    .b(_al_u75_o),
    .c(\ADD01/ADD02/n17 ),
    .d(_al_u86_o),
    .o(_al_u87_o));
  AL_MAP_LUT2 #(
    .EQN("~(B@A)"),
    .INIT(4'h9))
    _al_u88 (
    .a(n1[27]),
    .b(n2[27]),
    .o(\ADD01/ADD02/p0_lutinv ));
  AL_MAP_LUT4 #(
    .EQN("(~(A)*~(B)*~(C)*~(D)+A*B*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*~(B)*C*D+~(A)*B*C*D+A*B*C*D)"),
    .INIT(16'he699))
    _al_u89 (
    .a(_al_u87_o),
    .b(\ADD01/ctemp_lutinv ),
    .c(\ADD01/ADD02/n17 ),
    .d(\ADD01/ADD02/p0_lutinv ),
    .o(\exp_diff[4]_neg_lutinv ));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u90 (
    .a(_al_u67_o),
    .b(n1[17]),
    .c(n1[16]),
    .o(n93_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u91 (
    .a(_al_u67_o),
    .b(n1[19]),
    .c(n1[18]),
    .o(n91_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(B*~(A)*~((D@C))+B*A*~((D@C))+~(B)*A*(D@C)+B*A*(D@C))"),
    .INIT(16'h3553))
    _al_u92 (
    .a(n93_lutinv),
    .b(n91_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u92_o));
  AL_MAP_LUT5 #(
    .EQN("(~D*~C*(~E*~(A)*~(B)+~E*A*~(B)+~(~E)*A*B+~E*A*B))"),
    .INIT(32'h0008000b))
    _al_u93 (
    .a(_al_u71_o),
    .b(exp_diff[2]),
    .c(exp_diff[3]),
    .d(\exp_diff[4]_neg_lutinv ),
    .e(_al_u92_o),
    .o(_al_u93_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u94 (
    .a(_al_u67_o),
    .b(n1[7]),
    .c(n1[6]),
    .o(n103_lutinv));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u95 (
    .a(_al_u67_o),
    .b(n1[5]),
    .c(n1[4]),
    .o(n105_lutinv));
  AL_MAP_LUT4 #(
    .EQN("~(A*~(B)*~((D@C))+A*B*~((D@C))+~(A)*B*(D@C)+A*B*(D@C))"),
    .INIT(16'h5335))
    _al_u96 (
    .a(n103_lutinv),
    .b(n105_lutinv),
    .c(_al_u70_o),
    .d(_al_u67_o),
    .o(_al_u96_o));
  AL_MAP_LUT3 #(
    .EQN("(B*~(C)*~(A)+B*C*~(A)+~(B)*C*A+B*C*A)"),
    .INIT(8'he4))
    _al_u97 (
    .a(_al_u67_o),
    .b(n1[3]),
    .c(n1[2]),
    .o(n107_lutinv));
  AL_MAP_LUT4 #(
    .EQN("(A*~(B)*~(C)*~(D)+~(A)*~(B)*C*~(D)+A*~(B)*C*~(D)+A*B*C*~(D)+A*~(B)*~(C)*D+~(A)*B*~(C)*D+A*B*~(C)*D+~(A)*~(B)*C*D+A*~(B)*C*D+A*B*C*D)"),
    .INIT(16'hbeb2))
    _al_u98 (
    .a(n107_lutinv),
    .b(_al_u70_o),
    .c(_al_u67_o),
    .d(n1[1]),
    .o(_al_u98_o));
  AL_MAP_LUT4 #(
    .EQN("(~B*(~D*~(C)*~(A)+~D*C*~(A)+~(~D)*C*A+~D*C*A))"),
    .INIT(16'h2031))
    _al_u99 (
    .a(exp_diff[2]),
    .b(exp_diff[3]),
    .c(_al_u96_o),
    .d(_al_u98_o),
    .o(_al_u99_o));

endmodule 

