



`timescale 1ps/1ps
module TEST_TOP1(
    input wire i_clk,
    input wire[31:0] a,
    input wire[31:0] b,
    output reg[31:0] c,

        //串口接口
    input wire i_rx2,
    output wire o_tx2
);




endmodule