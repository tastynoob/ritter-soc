// Verilog netlist created by TD v5.0.38657
// Sun Feb 27 22:05:53 2022

`timescale 1ns / 1ps
module BRAM_ITCM  // bram_itcm.v(14)
  (
  addra,
  clka,
  dia,
  wea,
  doa
  );

  input [13:0] addra;  // bram_itcm.v(29)
  input clka;  // bram_itcm.v(31)
  input [31:0] dia;  // bram_itcm.v(28)
  input [3:0] wea;  // bram_itcm.v(30)
  output [31:0] doa;  // bram_itcm.v(26)

  parameter ADDR_WIDTH_A = 14;
  parameter ADDR_WIDTH_B = 14;
  parameter DATA_DEPTH_A = 16384;
  parameter DATA_DEPTH_B = 16384;
  parameter DATA_WIDTH_A = 32;
  parameter DATA_WIDTH_B = 32;
  parameter REGMODE_A = "NOREG";
  parameter WRITEMODE_A = "NORMAL";
  wire [0:0] addra_piped;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i0_008;
  wire inst_doa_i0_009;
  wire inst_doa_i0_010;
  wire inst_doa_i0_011;
  wire inst_doa_i0_012;
  wire inst_doa_i0_013;
  wire inst_doa_i0_014;
  wire inst_doa_i0_015;
  wire inst_doa_i0_016;
  wire inst_doa_i0_017;
  wire inst_doa_i0_018;
  wire inst_doa_i0_019;
  wire inst_doa_i0_020;
  wire inst_doa_i0_021;
  wire inst_doa_i0_022;
  wire inst_doa_i0_023;
  wire inst_doa_i0_024;
  wire inst_doa_i0_025;
  wire inst_doa_i0_026;
  wire inst_doa_i0_027;
  wire inst_doa_i0_028;
  wire inst_doa_i0_029;
  wire inst_doa_i0_030;
  wire inst_doa_i0_031;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i1_008;
  wire inst_doa_i1_009;
  wire inst_doa_i1_010;
  wire inst_doa_i1_011;
  wire inst_doa_i1_012;
  wire inst_doa_i1_013;
  wire inst_doa_i1_014;
  wire inst_doa_i1_015;
  wire inst_doa_i1_016;
  wire inst_doa_i1_017;
  wire inst_doa_i1_018;
  wire inst_doa_i1_019;
  wire inst_doa_i1_020;
  wire inst_doa_i1_021;
  wire inst_doa_i1_022;
  wire inst_doa_i1_023;
  wire inst_doa_i1_024;
  wire inst_doa_i1_025;
  wire inst_doa_i1_026;
  wire inst_doa_i1_027;
  wire inst_doa_i1_028;
  wire inst_doa_i1_029;
  wire inst_doa_i1_030;
  wire inst_doa_i1_031;

  AL_DFF_X addra_pipe (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[13]),
    .en(1'b1),
    .sr(1'b0),
    .ss(1'b0),
    .q(addra_piped));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'h5000011F08000000801B81E00000001FFFE01E4FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h00000407E000008080808080808000000000000000000000001F80003C445500),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n63,open_n64,addra[13]}),
    .dia({open_n68,open_n69,open_n70,open_n71,open_n72,open_n73,open_n74,dia[0],open_n75}),
    .wea(wea[0]),
    .doa({open_n90,open_n91,open_n92,open_n93,open_n94,open_n95,open_n96,open_n97,inst_doa_i0_000}));
  // address_offset=0;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1A(256'h4000003248000005001B06600000001FFFFFE04FFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1B(256'h00000405E0000080808080808080000000000000000000001F80000005E01001),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n123,open_n124,addra[13]}),
    .dia({open_n128,open_n129,open_n130,open_n131,open_n132,open_n133,open_n134,dia[1],open_n135}),
    .wea(wea[0]),
    .doa({open_n150,open_n151,open_n152,open_n153,open_n154,open_n155,open_n156,open_n157,inst_doa_i0_001}));
  // address_offset=0;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000880000C00C00060000800040060804110000060041011104107302C0A0155),
    .INIT_01(256'h80200108000C0003000029061008000300121830300118000066000020424000),
    .INIT_02(256'h142208440C10200801090820000010820090900080044480040044C080404100),
    .INIT_03(256'h000380040C60B200401918C600003860012100A0010800001000000000001102),
    .INIT_04(256'h04000000002C00000000400000820003000030118C0000380053231806000060),
    .INIT_05(256'h0100000000C080CCC198638C71C4803028430200004D240880C000C000000502),
    .INIT_06(256'h080403058602187260030218101A0209801811120140C0404006000100044870),
    .INIT_07(256'h3060C3030CDE02131A061830C100C36064C0C0660B00C360C4C0401248C10066),
    .INIT_08(256'h3060318008818060C18300003000A240810400C0C60630C00030000586280020),
    .INIT_09(256'h000080005800C03254080330B071818082000CC008006180C30C006303060227),
    .INIT_0A(256'h2C18C6199802410300C00D8124E00014231C0160048200012008021600001020),
    .INIT_0B(256'h04080601000C6018003018C40000404519000590208000000419400C00240300),
    .INIT_0C(256'h8000040C1400000220010042103000198180000000440000C021003118000060),
    .INIT_0D(256'h0824803000000000C0000402300C6018018182000A0000000000000048000801),
    .INIT_0E(256'h0200C08700218604C081AA00000006007000A000810000002060100630014000),
    .INIT_0F(256'h809902903460460C001600011406080990B04A019201003831C10E0006008800),
    .INIT_10(256'h0240000200000400000000184000008000000C04C81C04C81013210132080990),
    .INIT_11(256'h202020040201000803000004810200240D068004000800080008080000080800),
    .INIT_12(256'h0400305200000810404000100000208640081040841002410010408202010100),
    .INIT_13(256'h0040190068000A00000000000000800040000000001080100020111082040006),
    .INIT_14(256'h8010420000144044900220000028001000051200A81000000540000001008902),
    .INIT_15(256'h0000200008001808842204001800000181000200002408200800020000044044),
    .INIT_16(256'h000000C20000080000001A200000020000008038064004000000000000040002),
    .INIT_17(256'h6040000120041206834002000400000204000004000810000100009000002000),
    .INIT_18(256'h2002900A240050C8012088104080120020820820201020040404008040200100),
    .INIT_19(256'h2408041000120000000000081440010000800000420800800608200010006004),
    .INIT_1A(256'h5400018E40000005000106600000001FFFFFFF8932194A529414130508640000),
    .INIT_1B(256'h00000001E00C000000000000000000004123000080000000000018002AD55155),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n183,open_n184,addra[13]}),
    .dia({open_n188,open_n189,open_n190,open_n191,open_n192,open_n193,open_n194,dia[2],open_n195}),
    .wea(wea[0]),
    .doa({open_n210,open_n211,open_n212,open_n213,open_n214,open_n215,open_n216,open_n217,inst_doa_i0_002}));
  // address_offset=0;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0008000000000000000000000000008001100000000000000000040020000000),
    .INIT_01(256'h8020010800000000000020001000000000000000000000000000000000420000),
    .INIT_02(256'h1022004000000008000808000000008000808000000004000000000080004100),
    .INIT_03(256'h0000000000208200000108400000000001010080000800000000000000001100),
    .INIT_04(256'h0000000000000000000000000082000000000010800000000010210000000000),
    .INIT_05(256'h0100000000000000000000000000000020000000000504000000000000000502),
    .INIT_06(256'h0000000000000000000000000000000800001112010000000000000100044800),
    .INIT_07(256'h00000000000000100A0000000000000004000000000000000000000248010000),
    .INIT_08(256'h0000000008800000000000000000A24081000000000000000000000400280020),
    .INIT_09(256'h0000800040000030140800008010000082000000080000000000000000000224),
    .INIT_0A(256'h0000000000000000000000000000000021000000048000010008001000000000),
    .INIT_0B(256'h0000000000002000001000000000004001000080200000000401000000040000),
    .INIT_0C(256'h0000000014000002000000000000000000000000000000000020000100000000),
    .INIT_0D(256'h08240000000000000000000200000000000000000A0000000000000040000000),
    .INIT_0E(256'h020000000000000400802800000000000000A000800000000000000000010000),
    .INIT_0F(256'h0000000004000000000000010000000000804A00020000200000000002008800),
    .INIT_10(256'h0040000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h2020200400010008010000008102002401020004000800000008080000080800),
    .INIT_12(256'h0400004000000800000000000000208440081040841002410010408202010100),
    .INIT_13(256'h0040010008000000000000000000000000000000001080000020111082040000),
    .INIT_14(256'h8010020000044044900200000008000000011200A81000000540000001008902),
    .INIT_15(256'h0000000000000808842204000000000001000000000400000000000000044040),
    .INIT_16(256'h000000000000000000000A200000020000008008004000000000000000000000),
    .INIT_17(256'h2040000020041200810002000400000204000004000810000100000000000000),
    .INIT_18(256'h0000000000001088012080104080120020820820201020040404008000200100),
    .INIT_19(256'h2008000000120000000000001040000000000000020000800008000010000004),
    .INIT_1A(256'h400001C160000005800C07FFFFFFFFE000000010000000000000000000240000),
    .INIT_1B(256'h00080001E000800000000000000000073800B981800000000000000230444410),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n243,open_n244,addra[13]}),
    .dia({open_n248,open_n249,open_n250,open_n251,open_n252,open_n253,open_n254,dia[3],open_n255}),
    .wea(wea[0]),
    .doa({open_n270,open_n271,open_n272,open_n273,open_n274,open_n275,open_n276,open_n277,inst_doa_i0_003}));
  // address_offset=0;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hEB6140A047E67D35BFDBBBF00A413404A2494A28B08AD455AA4569DE569EC3FF),
    .INIT_01(256'h4B0D029228E5DC4DE7659BA3E0740015FCF74F9F17E308048C3308885395B35F),
    .INIT_02(256'hE3DCA7B3C70F5EA364F2F75EA20D4F75E84F2E5D7A43E27AEBD03E7142393AA1),
    .INIT_03(256'hC1068E0B35CA1C41204E31ABC4C46C23029E735004F5F1552EC4D248BC012E49),
    .INIT_04(256'h620267FFE7E61FFEFFDFD9F8010CA489D8421A231A155C6C60E9C63443A82639),
    .INIT_05(256'hDC4956ABBA43CE767EEFA6F4D34DF0DFD8D13D0000D86179D84E006FC0000A30),
    .INIT_06(256'h981E81FCFB86CCDE29F9C60B30EF0FD6FBEE2A8568FC40CBF88329626A51B3DF),
    .INIT_07(256'h1D3E7D75F76BFF6D354BE81F436C7D383B70402399D87D387C43C47DB76271BB),
    .INIT_08(256'hDC3E1EF84624FB3E72F5EFBBD7265DB66AEDAE7A7BB39F787A5FF240FB1262C1),
    .INIT_09(256'h890841C12F8E7206C98551DF5FAEBEF82955477942562EEE7DF76E3DF99BC1D9),
    .INIT_0A(256'h722E738CCD06C885D165D7436DBC012B063643212331C0D0502145C34050F45C),
    .INIT_0B(256'h1193890AC2E5C98C08668E7A0961309F0AA22B6C044047E0094EA107806025A0),
    .INIT_0C(256'hA8682285A8DDDDDD5AB4B6F7BDE82BCEFCD03FFEE26A0A005480841E0FE50036),
    .INIT_0D(256'h4153411D89EEFD3E56142A111E37BD4E00C6DF78159F8FF9C0FFFF9D24027FBC),
    .INIT_0E(256'h8444688DD112CA99672CC508B987C28FDA4D4FFE0B5FFFCFBE37A80B98EA347F),
    .INIT_0F(256'h41A9F54A90D1CA5698739F047222541A9D1D90DED094828D5D735B5868222114),
    .INIT_10(256'hAE3EF8D9C79FFDDF6FFEEFEDDFFFAB8FE3EF7A0D4FA20D4FA8353A8353D41A9D),
    .INIT_11(256'hD55FDFBBFF7EFF77EEFFFD5D7EF9D7DBB67DEFE3DBF7BEFBE96557FEB55557EE),
    .INIT_12(256'h0BFF94BD80F9F76BDFFD7FFEB818DF7BBF77EFBF6BEFDDBEFFAFBF7DF9F4FEFF),
    .INIT_13(256'h1F3AEAE3B637FEFFFE6FFCDFBE7FDFFFF9BFF37FFF8F7DF6AADDCEEF7DEBFFE3),
    .INIT_14(256'h422A34A8FFF9242948455451FFF6AA68BFFE453F57CFDDFDEABBEDFFD6FB40F9),
    .INIT_15(256'h7FFFF7FFFDFFF7B77BDDEBFFCA5FFFF8C2ED7D013FFBB5EFFFAFFFD78119242A),
    .INIT_16(256'h7FF77F6EFFFD58DFF1E7F5DFBBFBD5DF6FFB71D73ABF7DF6BFDFFFFFFFFEFFFF),
    .INIT_17(256'hDF3FFF575AFBEDDB3EF7F1EDFBDFBFF52BFF5AABE964AF8D96FDD58E0FFFEEFB),
    .INIT_18(256'hD7BD75FCD9BFEF77EE5F7BEFBF7EEDF7DF7DF7DF9F4FDFFAABFBF77FEFDFEEFD),
    .INIT_19(256'hDFF7FDB6FFECED79EF6D9EFF4F3FCEFFF7B8FFFFC1F7E77F7A97D67FEFEFBF0B),
    .INIT_1A(256'h410001AF30000000001A08600000000000000005EB35AD6B5B7B7ADEBB5B4BE6),
    .INIT_1B(256'h00000001FFF18000000000000000000702983C44000000002060678032AC1515),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n303,open_n304,addra[13]}),
    .dia({open_n308,open_n309,open_n310,open_n311,open_n312,open_n313,open_n314,dia[4],open_n315}),
    .wea(wea[0]),
    .doa({open_n330,open_n331,open_n332,open_n333,open_n334,open_n335,open_n336,open_n337,inst_doa_i0_004}));
  // address_offset=0;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h159E8061382D826A40245C0FF41244FB4193124953741C9951699621A9611400),
    .INIT_01(256'hB47A756D538A22A2188A245C1C88000A0308B060680075514244F777BC625CE4),
    .INIT_02(256'h1C23184C1830A14EA30D08A5E49A308A14B0D0C284CC15841424C182A4C27554),
    .INIT_03(256'h0A4951F58834E39AC0314A5438289254FD61A5A0030A38E0518C249543FC51C6),
    .INIT_04(256'h94015D63C039759CEE807147F2D349D222956554A40AA0929D1629480C52C8C5),
    .INIT_05(256'hA9B6291D4D82318981104108208382202526C2000227978BA6B89F903FFFD5CB),
    .INIT_06(256'h0711460F04019022560201740B1008690410555A9B00B0210754929594A7FCEE),
    .INIT_07(256'hA2C1828A089410120A941060809082C6448C82C4062082C680B02C4248858244),
    .INIT_08(256'h23C0610599C90441890A1F55A448A24EBD1E508484646086F5AC2497042C943A),
    .INIT_09(256'hAA32AA3E506884B9162A2E20A0514106D68AB8875DB451108208984202243A26),
    .INIT_0A(256'h8C50843332F135022E9B288C9243FED42948245AD7C60D65A04EAA1CB6AD5920),
    .INIT_0B(256'hE66C575555183A3156993084169E416F555594B2A880081FF6B140F87FB54256),
    .INIT_0C(256'h5817C51A57222222A54949CE727016110125E6D819D4687EAB3D02A1F0544FC9),
    .INIT_0D(256'hCE2C80227B8588C0A9F15402E14842B13F291087EA6F1B38179DA7035819B851),
    .INIT_0E(256'hB3CD81626E61156F8CD13E01D6DF957165B2BA98E5AAA781E04050346715CA18),
    .INIT_0F(256'h8C560AB567E3652800D420F9D46D28C562E64FF12BED0172A28884A797E6DF3D),
    .INIT_10(256'h5BDF7FE60601162693FD3F936FFF56FA9C11CC62B05C62B0518AC518AC28C562),
    .INIT_11(256'hAAE7FF654A9F3EC91B7FFAB791463BFD49D6991C25F8492DFF9ABFFD4AFABFD9),
    .INIT_12(256'hFCFC2BD200C008BA32D2805947E728FE7EC9144F9D1FB3DF27D448BE468F11FF),
    .INIT_13(256'hEFE4155049DF4FF715BB3B76DFF4FEF2D6ECEDD8507092595522B110821CBE04),
    .INIT_14(256'hBFF5CF7F0A16DBDEB7FEEBFE142F57B74285BACEADF4227B5544D37E2984BF46),
    .INIT_15(256'hFBB9BFADCFEF184884221CFC15E02F813F12820018245D115A5007287EE6DBDD),
    .INIT_16(256'h9FE9FC9B7FFABFA24E1A9A2844F6AA269BF6C82C85489669462E2EF7FFB7F76B),
    .INIT_17(256'h68DFFEADE77D1EA4EB4C8E12FC2244FADFFEA57D1F9B747E6BFB2BF00C08B134),
    .INIT_18(256'hAF6ADA8B7E4C5FCFD9E8ADF44FFD9EFBE8BE8BE468F23FF55CFFECA953E7D923),
    .INIT_19(256'hB60A16797893CAF0DE5B331AB4C83F180AEF0304422900A69568A06014D146F7),
    .INIT_1A(256'h100000AD40000001000F8D60000000000000001A958A5294A6464791A4E55558),
    .INIT_1B(256'h00080001FFFC800000000000000000067920467E800000004000007FA2914501),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n363,open_n364,addra[13]}),
    .dia({open_n368,open_n369,open_n370,open_n371,open_n372,open_n373,open_n374,dia[5],open_n375}),
    .wea(wea[0]),
    .doa({open_n390,open_n391,open_n392,open_n393,open_n394,open_n395,open_n396,open_n397,inst_doa_i0_005}));
  // address_offset=0;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h108880011801824A402404000410408041101040400408001020062029210400),
    .INIT_01(256'h84625569120822A20002241C1008000A00083060600010004044000020424880),
    .INIT_02(256'h1C23184C1830A14C830D08A14492308A14B0D082848C15841424C182A4C24544),
    .INIT_03(256'h0A0950048820E21A40314A5428289254016100A0030A08A05108208440001186),
    .INIT_04(256'h9401100000194000000020040092481222002554A400A092801629480C5200C4),
    .INIT_05(256'h212609044180218981104108208002202406020000051602048080900000054A),
    .INIT_06(256'h0701460304011020400201700B10002904105112810080200704801104244820),
    .INIT_07(256'h22C18282089400120A94106080808240448082C4060082408080200248850244),
    .INIT_08(256'h23C0610499C90441890A10442048A240951250848444208685A0049704281428),
    .INIT_09(256'h2222AA00504084B8142A2E20A05141049682B88619A041108208004202243226),
    .INIT_0A(256'h0C1084111080050202800880004000142948244A14860905200AAA14A2A10920),
    .INIT_0B(256'h062C161505182031001130840080404051440492A88008000491400800154240),
    .INIT_0C(256'h1010040815222222214949084210001101058000000400408821022130104048),
    .INIT_0D(256'h8C248020500100C08800040221484211012900800A2000001200000248098041),
    .INIT_0E(256'h320980222061140480812A00040014502000A000A4800000004050046001CA00),
    .INIT_0F(256'h845002916420240800042001040C084500E24A210A290070A08884A006049821),
    .INIT_10(256'h51C1072600000220900110122000547000000422801C2280108A0108A0084500),
    .INIT_11(256'h2AA0204400810088110002A2810628244982101C24084104169AA8014AAAA811),
    .INIT_12(256'h94002342000008902002800140002084408810409410224100504082060B0100),
    .INIT_13(256'hE0C4111049C80100019003204180200006400C80007082095522311082140004),
    .INIT_14(256'hBDD5CB570006DBD6B7BAABAE000955974001BAC0A8302202154412002904BF06),
    .INIT_15(256'h80000800020008488422140011A000012512820000044810005000280006DBD5),
    .INIT_16(256'h800880910002A72000000A2044042A2090048828844082094020000000010000),
    .INIT_17(256'h20C000A8A5041224C1080E120420400AD400A554169B507269022A7000001104),
    .INIT_18(256'h28428A032640108811A08410408112082082082060B020055404088010201102),
    .INIT_19(256'h200802490012020010122000B0C0310008400000020800808508200010104084),
    .INIT_1A(256'h5100014938000005800887E00000000000000018108842108404050104A41010),
    .INIT_1B(256'h00080405FFFD8080808080808080000438003DEF800000000080800024DB5541),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n423,open_n424,addra[13]}),
    .dia({open_n428,open_n429,open_n430,open_n431,open_n432,open_n433,open_n434,dia[6],open_n435}),
    .wea(wea[0]),
    .doa({open_n450,open_n451,open_n452,open_n453,open_n454,open_n455,open_n456,open_n457,inst_doa_i0_006}));
  // address_offset=0;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hCF41152A8E92E911E99B802000B9ED00146D6AAAF4007E770077C3741F1988C3),
    .INIT_01(256'h090C0AE7A0AC515F26545FE74272AAA750B7DD3AB5749A02A46F00800AAD8774),
    .INIT_02(256'hAD59DA9DAEB5AA96375755EA0B5D755EA1357573AF5D29AF5D7AD2E82BD4A0EA),
    .INIT_03(256'h55A7A200B1C170200ABA718E875678E9006AF40AA950335CB4F58368940184D6),
    .INIT_04(256'h8954776764CEDDB3700A5A200404DAA7556AB2A718A15C7902C74E3296AD156A),
    .INIT_05(256'h044956AA10EB88ECE9DD77CEFBEDE5B29ED328AAA4D8682889CA60C240002060),
    .INIT_06(256'h5CDC27AFD7463AF86807A89A8699AEC1D59D22A5EC06CCD3E8AE612A6A1101F1),
    .INIT_07(256'h7574EB2FAEDF56EBB05F5D3AE852EB6872E2EB775BB5EB68E0CAD77523D044F7),
    .INIT_08(256'h74E8F79A41239AE6D7972C98779A0997604486D3DE9EB2C96A39B223D6800B04),
    .INIT_09(256'h558A0080B9F5D646C11377F232E1979B3136AFCDE21CE5A2DB5D28EB1346448B),
    .INIT_0A(256'h60BCE719990EC22B80E183136DE800005EB11BE4092A78160AB03E666952F66B),
    .INIT_0B(256'h0A0620200841C5DAA96759E8A9208A9B78A86055472A9440019A0A0D0062B709),
    .INIT_0C(256'hA6A8102D0059994C4212042104854BBB85CABD6324208D81C0402B741A653060),
    .INIT_0D(256'h54432A781D48B22AC21AA0A4343D651A0197D968003F6C4D6AFDFF59A2A459A1),
    .INIT_0E(256'h6422149F8085C680C52384523803CE0FB0480CC31B8EBFEB316C854EB068947C),
    .INIT_0F(256'h13B9400288C5CE812D4ED30248B6813B907600A5841654D975D71E58602A2124),
    .INIT_10(256'hA62490C0AFABBD904C0805D8145629846182009DCA009DCA0277202773013B90),
    .INIT_11(256'hC55A04308FE48127F6A16D4C74D5F4016CE1BFE35E859FDA496150B6B551510C),
    .INIT_12(256'h0A1DB014D5F2A50F1C150352A0089F128177EFB27BE0DC208E6D3A49F9A8FE29),
    .INIT_13(256'h008CB85960302212442AC000024C0EB160081039DC092F34DFC9CAAA594B1A96),
    .INIT_14(256'h6C4A1C80B933BD336989C401726157A0274CA8CD0020ED0D3A122C84AC2F3624),
    .INIT_15(256'h2CDFA3A4386345D352C548C2D877485D82AF70AC655891E3240AE8008013BD31),
    .INIT_16(256'h68446EC0B25D48D890C5015C48F97D5B26E82D72AE2B4DB286DB29B8220EF2F8),
    .INIT_17(256'h92AC5B534C8A41B6704E208F60CCF6D5285358AA0964A905962D94855D56E4CB),
    .INIT_18(256'hCB80012D481CC7406C905E692706C074D00524D1508884BAA960B631FCD52442),
    .INIT_19(256'hCA32624477009E5B8CE31295488DCE4040205358B0E3AA5726078CEFCE8BE702),
    .INIT_1A(256'h0540010C00000000000B00600000000000000000607084210870721C3949D9D3),
    .INIT_1B(256'h00000001E00C000000000000000000033EDF467E000000000000000002F10154),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n483,open_n484,addra[13]}),
    .dia({open_n488,open_n489,open_n490,open_n491,open_n492,open_n493,open_n494,dia[7],open_n495}),
    .wea(wea[0]),
    .doa({open_n510,open_n511,open_n512,open_n513,open_n514,open_n515,open_n516,open_n517,inst_doa_i0_007}));
  // address_offset=0;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h6B6066A6C31631918CC92B800A6D9F00A26DEFBE8C0AF77728D7C8CC529EE0FF),
    .INIT_01(256'h428D8A96ACD151548665C0E183373310CCC1C60C867B02AE219808805FB5B622),
    .INIT_02(256'h8310C60280CC18A378C2C6581B6D8C65810C2C79637308638B1B300D5B31BAAA),
    .INIT_03(256'hF5A6240B77CB08652C4631A98756648A0298BD5CC4C55606AC57DB6A8402A871),
    .INIT_04(256'h0A62E6F4B58096586A948EA0052CB6ACDD6A8AA31B150E6520E8C63741AD371B),
    .INIT_05(256'hDE4992CBB833CC0230660670C30DFCCE5AD831CCD1D8682D890F602300002A24),
    .INIT_06(256'h98FEA0CC0196A00301CCCE833486CF9062E60AA16CE30A1DD8A94D6A6B58B3CB),
    .INIT_07(256'h4D18000CC02198A03029860C331F301900303100783130180E0CD581B5224D01),
    .INIT_08(256'hCC1C8C4A66364A923454ABBBCFB715254AE5AB3139998E295A4F7B48010362C4),
    .INIT_09(256'hDDC55441A4BD3346E150D0CB4986324B29654329E2498E6838F36B9898D94510),
    .INIT_0A(256'h72252944410ECAC4902417436D98042B16B65B842B3932DA5C3155214952F4D3),
    .INIT_0B(256'h191329AAEAE7CDC6A966C7030921B09F80A84B2D46734700090631030068B0A8),
    .INIT_0C(256'h27803A8128CCCCD15AA6B6F7BDEE23864C5A36FBA06A1F0110C2C54C060FA014),
    .INIT_0D(256'h71534D0D8DF82812141A8AD00C93150600521F58101FEFBFA0DACCE5A70600B8),
    .INIT_0E(256'h0C74689C0192409017264568A007E089C2094FD9130FFFB40099AE0980E23557),
    .INIT_0F(256'h43A1654A98D1D896E17859067A30943A190C109E5406E2854D37391008102080),
    .INIT_10(256'hA4269859F116DDDB69F6ADE4D7EBA905A2A4521D0B221D0B2874328743943A19),
    .INIT_11(256'hD153DF997E2638566C37DD594EB8C45B3220EE41D2F7B29AE94053EEB15057E6),
    .INIT_12(256'h018A841DE6F9B04CDA3516A0A800D21BBE544913626F95A636ABA71D9174C6F2),
    .INIT_13(256'h090AE283902326914005185E3C11807D61031204478165B4AACCC00D65A2E161),
    .INIT_14(256'h002020081AB80000000410103576AA488E2E0023044AC56C421B647BC42900C8),
    .INIT_15(256'h1B12B43BC59E6133738DC1FF424FF2B8402565CB2111B7E67FA7F25180180002),
    .INIT_16(256'h4B316F2EBB1D588641A2F450181BD451653811C730A16D12B15190A9ADD2F6CA),
    .INIT_17(256'hD20ED35648DA4199106620C969DCA4C52AD35AAAA944A805861D958F80B6E6C2),
    .INIT_18(256'hD72171B4D98DE361EC101AE9031EC434D03501D11548963A28687633C5C50A41),
    .INIT_19(256'h57A6BD36AEE8FD76600C847D4C1B4EFAE5A8E5B0E8F7E75F7813D66A8BE2110B),
    .INIT_1A(256'h140001F910000005000986600000001FFFE01E65EB75AD6B5BFBFAFEFB58ABE2),
    .INIT_1B(256'h00000405FFF98000000000000000000747FFFB9180000000001F8000032CC500),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_008 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n543,open_n544,addra[13]}),
    .dia({open_n548,open_n549,open_n550,open_n551,open_n552,open_n553,open_n554,dia[8],open_n555}),
    .wea(wea[1]),
    .doa({open_n570,open_n571,open_n572,open_n573,open_n574,open_n575,open_n576,open_n577,inst_doa_i0_008}));
  // address_offset=0;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h5AE33826E0F20FB6949F2B3E802F8F6900EDFFFE8F507F7F41FFD04492012F00),
    .INIT_01(256'h4BCD8EB3BCF29FEC137EDBB86B703C003CFF61C3C9E3C6EAB588B22581BC8F7E),
    .INIT_02(256'h68DDE1B96323C6F37E3637C6BBEDA30C6B6323FF1B78EA1BE8FB8F330F8FBEEF),
    .INIT_03(256'h1FAE71A074CB046C102073886596609C54067B0F02311E0FA2FFE36EA25BCE78),
    .INIT_04(256'h0981EF775232BFFFFFF78E46B42DF2AC3FEFC367380D7E6111C00670002D3502),
    .INIT_05(256'h344DB2EFB40FDC300C619E53CF3C8501DAD84C0F01D8782F8D2BB3143DB2A024),
    .INIT_06(256'h7DFFEC3E187663CD06943FE0FDA03FA21CC1AC29CC0B25F7D9A83A7ACB598141),
    .INIT_07(256'h43860CFC330066A0F4F861C30C9B0C84980B0D19983F0C853213DE7D211E6C98),
    .INIT_08(256'h02858236E072308C0E285AB8479341175062970B00284117DB0C3B6818D32B8C),
    .INIT_09(256'h778B3C6C833B0F46E955F80507024C3729F5E013E0FF820D0C003B846C00B488),
    .INIT_0A(256'hE02210A021AED6004A106403EF8556800E74331E9868DA90C073D4C865D6FFCD),
    .INIT_0B(256'h8BB5B8200D14D7E0F96FC018192C809FE6ED1003C83C0E7E81000090AAF9F00C),
    .INIT_0C(256'h4254D89209DFFFFD4ABE1DEF76E007A03227FFF909101FE62A5201C26197E989),
    .INIT_0D(256'h73DA30000260FA7F2AC851000200890066387F89A09FFFFFF9DFFFEDA00E6E3A),
    .INIT_0E(256'hED7F41FC0C80314805321480201FE821CC905FDF38EDF97EE680C028421415A9),
    .INIT_0F(256'h03A7800393C3F90418F981D2F871003A700214B41C3E00C1030F383491BF25D6),
    .INIT_10(256'hA69DF778068A9C95EA6EC7E0DD567DBDC6BCC01D2C001D2C0074A0074A003A70),
    .INIT_11(256'hC54604721E3C47F47E636F7E44944481B03C8CF91781F3BFDD6771B6A745D11C),
    .INIT_12(256'hAA1F411878D8B40CCC355673C52697720DF4EB8E32637C0C472922393D2046AD),
    .INIT_13(256'h2909C0DC81B5FB7FE6FFFAFF7FFF8FF575FF75FFE6886FBCEA8DC8894D2A3BD8),
    .INIT_14(256'h570F99F3AEBBACAB68F90DE35D75FF45EBAEA0AB146ACD6DEA1B7CD6A42F22FC),
    .INIT_15(256'h12F3D46BAD0C719063018195E19572AE2C2D60F00518266B442AD014DE1135B9),
    .INIT_16(256'h53773F01E94FFF5E6BB6B452391BD455ED3B0780F821EF1EB1511009875EF042),
    .INIT_17(256'h929A9B7F08A240D81E662CC9C9F8AAF4BA9B50A21DE2E925F23697E00DF4E7AF),
    .INIT_18(256'hC3AC0EFD0899EE61B4153FC90E1B44EF9509239150E89298A8C8DA43D788FE57),
    .INIT_19(256'h1FF7FFB2FBAC48A4BB0FFDCFCEBEFE1BF7C28F7798E1E357F843806ECAEB8152),
    .INIT_1A(256'h051001D310000000800581E00000001FFFFFE04166738CE33971765C3F5BEBFC),
    .INIT_1B(256'h00000001E005800000000000000000003800C391000000001F800000009C0504),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n603,open_n604,addra[13]}),
    .dia({open_n608,open_n609,open_n610,open_n611,open_n612,open_n613,open_n614,dia[9],open_n615}),
    .wea(wea[1]),
    .doa({open_n630,open_n631,open_n632,open_n633,open_n634,open_n635,open_n636,open_n637,inst_doa_i0_009}));
  // address_offset=0;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h5BE301B6F3D23F9A9CBBBA4A516F9F5F1AEDEFFE9FB1F7FFC4FFF0CF939FC7F0),
    .INIT_01(256'h2F8D9EF3BCB1D3F48777C0B9EF73C0D4F88967CFCFFF67AEEF11866B93BD9F7C),
    .INIT_02(256'hE3C1C7B3F3EF1FF7FAF2F05E5F6F6F75E52F6F637F73E87F0BFB3F3F5F3FBEEE),
    .INIT_03(256'h3DF66B93F3CB4C7C8346F7B9F71F6599F01E7B0034F4BFDFAEF7236EDA7680F5),
    .INIT_04(256'h281AFFF7F3E1FFFFFFE71E0D9E7DFFFCDDEE8BEF78DDFF65D6C4DEF0E1EF3F1F),
    .INIT_05(256'hF469D7D0073FFF333E079E23CF3FEC07DAD8FCF039D87B7DDD1FF428D49E6234),
    .INIT_06(256'hF89FB0FC79F727CD0BACFFA3F4C7FFC47FC7EAE5FCD70FD7FCA9EBEAFB5A35CF),
    .INIT_07(256'h4D9F3CBCF321F1ECF1F9E78F3C7B3C981B333F19FCF73C98321FF7FDB71E5E19),
    .INIT_08(256'hCD9A8C7BF67A799E3478F5FBCFFF4DAD7E8FFB3D31E9CB3D2F03FBF878C36FCD),
    .INIT_09(256'hFFC975EA87FD374EE1F3FC4E0E887C7F3D75C138B3FD8E7B34F3BD9CF4F1FC40),
    .INIT_0A(256'h616739E647BFF234F139C323FD9E27C996F0DF97D87DFF90C373F5E14BF3FEDF),
    .INIT_0B(256'hA88691BA6BC3D7C7B9EEC538C9669C9FA6AFE34DD900E09651C68DE3CC7ABC9D),
    .INIT_0C(256'h7E7D98C3C9DFFFFD5BFEF7FFFFE1ABE6767A7FFBAED11FA93F5237CE87EFFA12),
    .INIT_0D(256'hF3DB038C4FF9FFBB318F60390EA31D66A85C7FAF849FFFFBF1FFE7B7A0CC6EE2),
    .INIT_0E(256'hDC771ABCF68A69E9372E441CBDF7E9B7C5CE1FDF1F6FFFFEE61E8189CBB8BFFF),
    .INIT_0F(256'h27E7F94AC9CBD9E19BF9E7CAF931E27E7E4FB0DE5C961A850D3FF85DE03B21D6),
    .INIT_10(256'hE61DF144CFDE9FD56E6EF7E5FD57B9DDCDBA413F2FC13F2FC4FCFC4FCFE27E7E),
    .INIT_11(256'hDFCE04321F7CC7746EE36F7D6EBD4F81B2FCFCF9DB87B2FBD9E7F1B7BFD7D10D),
    .INIT_12(256'h62BFCC3C81FDF78FDCFD3D0D9CBD97738F76EBAE3263DC1CC72BB7793D7866AD),
    .INIT_13(256'hA8AFE63D903FFFFFE67AE1A5677FAF7DBBFFFFD3E4AB7FF4FADFEAE210514459),
    .INIT_14(256'h7F6F38BCBCBBB72B6BF51E797973130B6FAE2089162FDDEDEABBEDFF84AF4059),
    .INIT_15(256'h9BE7DFF10F9777F2084038D7E7C14FFE7AFF5C05BFF8566F2CF28FFACBB1BE3B),
    .INIT_16(256'h737FBF20E14FFCDDEBCE31DFFBFBFDFF6FFB7FC379BFFDF6EFDFFFEFBFD3FA8E),
    .INIT_17(256'hD23A1BD35DA240D97E7F20FDCBDCFAFD2A1BFABAA9F7E917BE3CB7A66FF4FFAB),
    .INIT_18(256'hDFAD7FFDDB9DEE7164157FC93E1641EF95492799156C829AEBC0F243EF98EED6),
    .INIT_19(256'h5FF7FFF6FFECFDD2FB1DDDFF4E3FDE7BFFE96B57F9F3F77F78E7CF7FEFFF9FB3),
    .INIT_1A(256'h144001F210000000801101E00000001FFFFFFF97EBF7AD6F7BFBFAFEFFDBFBFE),
    .INIT_1B(256'h00080001E00180000000000000000000000043910000000000001C00032E9040),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n663,open_n664,addra[13]}),
    .dia({open_n668,open_n669,open_n670,open_n671,open_n672,open_n673,open_n674,dia[10],open_n675}),
    .wea(wea[1]),
    .doa({open_n690,open_n691,open_n692,open_n693,open_n694,open_n695,open_n696,open_n697,inst_doa_i0_010}));
  // address_offset=0;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h80003E000025002D034405B9C010003800000040010008004000800193200400),
    .INIT_01(256'h7052646043422E2860011F000003FF0C06760040481C80005A886E9780200C21),
    .INIT_02(256'h001D20001020C10004000780A090E0700A60001C04801304E004800004820055),
    .INIT_03(256'hC20014F08000001B1C00000008E802063CC0004FC20140204000F88025314E88),
    .INIT_04(256'hD1E118080C136202004F61F4720041102000454401008082A008000300420084),
    .INIT_05(256'h2AB04C3FF800200000600050000211C8000440FFC00011505400000F246610C9),
    .INIT_06(256'h036058026008C4028E780020006700760320008422FC00082300050420A38600),
    .INIT_07(256'h020130C800201F4C0410000003F400818300000004E800810D10280096242380),
    .INIT_08(256'h0305420411440601020C1E0000041CBA2EE96C0608504402F14CC41261104448),
    .INIT_09(256'h0206081E20260C8008242081410E420614803201522210160860460008083198),
    .INIT_0A(256'h004000000240004000040008000380000000000AD304004E0C00080884210000),
    .INIT_0B(256'h022010100510082044010201149E000040059022863F0F71C000103070004060),
    .INIT_0C(256'h0184011000200000014808000006100008054004403000000308420020100004),
    .INIT_0D(256'h86083C03820700440F50C1C000508200400A0053613254C1C305238583193544),
    .INIT_0E(256'h2008000000401060005010E0064800180B80112044B1082DBD01663047448200),
    .INIT_0F(256'h0040000102000000600038B80040000420020020282060004008010390041021),
    .INIT_10(256'h49A20C803001622A8191180002A8526F7C49A802000002000008400080000420),
    .INIT_11(256'h0091DFC9E0023883801C90021040B85A0081030A24704D04A4940648022427F3),
    .INIT_12(256'h994001807E000060030242F26463080838810411498E21A238840814C0869852),
    .INIT_13(256'hB71400C207491825F9D71F7E9911D02606400CA9BB64000A5100040D6DBABBA0),
    .INIT_14(256'h2CC50C05654002902618C304CA8050A059D04DD441C00012100410005A5414A4),
    .INIT_15(256'h64EB60645D609005739DC328011EB000201020FA0003A180D34D702D46601A90),
    .INIT_16(256'h0C88401F16F22334361D040000042000800000040000820810000010C2228531),
    .INIT_17(256'h0D8564288259AD200080D502302307100164A0014603469860E36261800B0154),
    .INIT_18(256'h08100A01002205071ACA00A68571A8504A34D146CA834DE010338D3C01471028),
    .INIT_19(256'h800000090001008997E26200818020040010180A040000008000000000000080),
    .INIT_1A(256'h101401BE10000001800E01FFFFFFFFE000000000008000802000000004001009),
    .INIT_1B(256'h00000405E0018000000000000000000000003C6E8000000000000042079FA145),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_011 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n723,open_n724,addra[13]}),
    .dia({open_n728,open_n729,open_n730,open_n731,open_n732,open_n733,open_n734,dia[11],open_n735}),
    .wea(wea[1]),
    .doa({open_n750,open_n751,open_n752,open_n753,open_n754,open_n755,open_n756,open_n757,inst_doa_i0_011}));
  // address_offset=0;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h1088000014004246202084000000000001001000000040440004050000200411),
    .INIT_01(256'h8241556808000A20000324101020000800482850406000000422000000420000),
    .INIT_02(256'h1822004000000088800C0001060200001480C0000280440400100142A6034120),
    .INIT_03(256'hC18A40008060C20200015A802806A21001010080020208A401C0304040001100),
    .INIT_04(256'h1000339D40004E6E318010100097380C16A69035A808FEA200502B50084C0080),
    .INIT_05(256'h200008004100C005008802844104604828440000004C3653540800100000050A),
    .INIT_06(256'h0502010080010000200001200301018085003912004440427C02800000046816),
    .INIT_07(256'h13A0408004020011081200100080000024404020010000000040000A4A420220),
    .INIT_08(256'h1020108488408021408910421208A240900AC044420210440590040682281420),
    .INIT_09(256'h01A80240C8404000142A39109030C08084026446092020904104202141022225),
    .INIT_0A(256'h000000000080040000400001248006002B50150804C80911805A081202B0C180),
    .INIT_0B(256'h02040100401476CA111BE80000208053086C4081E800080004810000001C4040),
    .INIT_0C(256'h10100000147BBB6E42D415AD6640010020001B28000002000820021009510008),
    .INIT_0D(256'h8826000008805480000400020120010100240A080A12A41C08664D0140010508),
    .INIT_0E(256'h220900A42000800461802800008500171000A768800759801420000240010001),
    .INIT_0F(256'h004000010D43708001D84103D800800C90C14A08182000408109882042049821),
    .INIT_10(256'h00C9A134019EF0322AB80B01346E002563EF4002000002400009000090000480),
    .INIT_11(256'h2022AA26B8A9144CF1237000CFBE253541B204EC26AB97A682D801B800280289),
    .INIT_12(256'h0458004000388881010C7C263810B7A4544CFBC496F51349591BE7933B794F37),
    .INIT_13(256'h22E401500809E108E915E22B881E211E245788AFEC10EC4FC022111082142C00),
    .INIT_14(256'h39400054DACE4844B72A0829B59D158236B39243A8B3E4A9154645AE2149BBBA),
    .INIT_15(256'h844F8853E213C848842214580839CB0081100000078440A0218F88C681164840),
    .INIT_16(256'h55C05849A370021D91E78A27C95222322D74C81C82771322C9F1F13B227108D8),
    .INIT_17(256'h37C8DC0024A6FAA2D902763357C9EB2200DC0012F2D80BD34851202003F78991),
    .INIT_18(256'h8A400BA4103E348A8937A69BC4A89A4D37937933B799E6E4045544D71522895E),
    .INIT_19(256'h308DF02A8F70823024020824107710078818CC7F02E0E074400B801E0E8C0105),
    .INIT_1A(256'h050000EC00000000000800600000000000000000000000000018180608A45090),
    .INIT_1B(256'h00000001E000800000000000000000007FFF8000000000002060638006719054),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_012 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n783,open_n784,addra[13]}),
    .dia({open_n788,open_n789,open_n790,open_n791,open_n792,open_n793,open_n794,dia[12],open_n795}),
    .wea(wea[1]),
    .doa({open_n810,open_n811,open_n812,open_n813,open_n814,open_n815,open_n816,open_n817,inst_doa_i0_012}));
  // address_offset=0;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000A3F5FA01800040000800FF1AE837B1DA4A1860F7167EE451E140181613C10),
    .INIT_01(256'hB291A9084D12291018B964021FA3FFE003480000981CEFFB278AF77780420804),
    .INIT_02(256'h1022404020C00098180800001B6080000380812003704C01001B000E9B05C13A),
    .INIT_03(256'hF572A1F0026582A49F819C80111529A8FD01008FF800060E80D31D7103FED130),
    .INIT_04(256'h89FC9D015804F40D20A02603FEE6A369115B50B9C9E651291F503393B2095922),
    .INIT_05(256'h0290A150043CB00000081A074D370D502B68C0FFFF6EA98D23717F403FFFF5C7),
    .INIT_06(256'h68E43900807A2B4196043A84D402F2808001B57A16477F564978D68C918E4C08),
    .INIT_07(256'h4120410004020291D80207907D030087A44F7D3869070087077C5B92485A0C20),
    .INIT_08(256'h0001800328120080040000020891A24980080101000840010000092C82E80836),
    .INIT_09(256'h5555147E40114973745810008010000180004001E81D90010004B18004400E24),
    .INIT_0A(256'h81C10862227932782C1A203C9203F8C0F1818894CCA0363B4FAC10381D0E8A03),
    .INIT_0B(256'hE800014050022980EE968101F63E0F77A43191A0B33FB01FF6211EF07F86981F),
    .INIT_0C(256'h4787D97256111102849600842047D420022A42091D91F5BF237E79C0C00ABF81),
    .INIT_0D(256'h3EAC3EC23710420121EBD1EEC08001A0FE10200FEA62581A27840561D3F48042),
    .INIT_0E(256'h6BB317500E8CA16658D23CF742FA292515B2BA09D4AA01B041A807F207158980),
    .INIT_0F(256'h3A060805068D4121665001F951D123A0E2816F0825627D02020420A7D3D9DECA),
    .INIT_10(256'h084820D03E65100229C0040904B002029F11C1D07041D0704741C4741C23A0E2),
    .INIT_11(256'h2062FC0568093809092580109142113C0532090400BA08A0894812C000481700),
    .INIT_12(256'h6C2058C07FC60924209010480FE728A4780914448D1E03C92114489242851158),
    .INIT_13(256'h62C10D0C2CC94100119903320894201286640CC81030D04080201330820C101A),
    .INIT_14(256'h022004284A86C94C90464050950E022012A13302A8B404F0054044F00109A946),
    .INIT_15(256'h80098801C203080984260C20244104061B0000FED804923012020500FEE6C948),
    .INIT_16(256'h4E00200826801002DE1A8A2809E002022780860841681022868E28B722310048),
    .INIT_17(256'h2849600422251E00990482205F022422096000210948240D02E00101FC288811),
    .INIT_18(256'h002000A0582C148F0168A09444F01E412892892428522D040C5F80AD01270121),
    .INIT_19(256'h308B1022F89110C60881591010680E18002F03043E011800406809E000080076),
    .INIT_1A(256'h401000CE00000005800805600000000000000003265318C63000040004A5E409),
    .INIT_1B(256'h00000001E0018000000000000000000000000000000000000000003FC54C9950),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_013 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n843,open_n844,addra[13]}),
    .dia({open_n848,open_n849,open_n850,open_n851,open_n852,open_n853,open_n854,dia[13],open_n855}),
    .wea(wea[1]),
    .doa({open_n870,open_n871,open_n872,open_n873,open_n874,open_n875,open_n876,open_n877,inst_doa_i0_013}));
  // address_offset=0;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h1088000104004084000094000010080001000410000044440084040001210410),
    .INIT_01(256'h820111088A002A800021241210200000004828501040080014000000004A08C4),
    .INIT_02(256'h10230040040000CC8008000142920000148080800240540400140042A2014524),
    .INIT_03(256'hC18200004060820A000118802206200001010880000008840068104240001180),
    .INIT_04(256'h8000159D4010566E318030040086A00C146280318804582000502310000C0004),
    .INIT_05(256'h200409044140A045408022805145404828410000004C21414400000000000542),
    .INIT_06(256'h0B05440A0202005020010328100B028001083112804400426D0080100004481C),
    .INIT_07(256'h01010001004802101830084001004120040000820C004120440040124A020202),
    .INIT_08(256'h0002400098480001000810420008A24094081004000000040580008400290120),
    .INIT_09(256'h01A02840C04044B2540894008010000084205005591400000004200000002224),
    .INIT_0A(256'h200000000002000000000000000000002310010004AC0811403800100020C880),
    .INIT_0B(256'h000000A028006DC00916800000208047402C01A0E80000000401000000044000),
    .INIT_0C(256'h101000001459994A429448842040000000048B28000000000020000000000000),
    .INIT_0D(256'h0C240000190040C00804000200200100000402080A32A81C0AA64D0140018040),
    .INIT_0E(256'h220100842000800440802C00000600071000AB68848B59800020400200018800),
    .INIT_0F(256'h0089000104815000005801035808000810814A0810280040010108A042009800),
    .INIT_10(256'h48C100D0068750202B49150120D25222E3A74004080004080010200102000810),
    .INIT_11(256'h206074277881284D4906A290D9E2182C41320D84041B1CA40948135140481509),
    .INIT_12(256'h0C3000C000D009207098744A3800BC84684D9E408F5A12C1701E6C8363C5556C),
    .INIT_13(256'h60C401100CC96108D199A3338096211E86668CCB7830F24AC0221330820C1800),
    .INIT_14(256'h12200428DACEC9CC92464051B59A022036B33300A83684D1154405D40961A976),
    .INIT_15(256'h840F8851E213C80984260C3000594600030000001A049011130E85868016C9C8),
    .INIT_16(256'h5A48A8090592924BD0C78A2D09A22A202EC0880880799202CEEEC88C00310858),
    .INIT_17(256'h3C41A8A4230796209906C2220F8B2E0209A8A02389482E0D12A129200D3A8901),
    .INIT_18(256'h02602BA4482F308D097CA41E40D096083C83C8363C5B2B240C0E84EF10250971),
    .INIT_19(256'h310F5022F390805008011814B0790E1A08B8471D02818044C00A0068089C0307),
    .INIT_1A(256'h1411015B10000005801A87E000000000000000000000000000888C2244A50010),
    .INIT_1B(256'h00000405E000000000000000000000007FFFFFFF800000000080800004E96501),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_014 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n903,open_n904,addra[13]}),
    .dia({open_n908,open_n909,open_n910,open_n911,open_n912,open_n913,open_n914,dia[14],open_n915}),
    .wea(wea[1]),
    .doa({open_n930,open_n931,open_n932,open_n933,open_n934,open_n935,open_n936,open_n937,inst_doa_i0_014}));
  // address_offset=0;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h908D80A1090490E24824C0A004415800434A44114004E866112606A80811B482),
    .INIT_01(256'h884C41492208628285023615F3780002882C162E276012AAC0540088224F4B7C),
    .INIT_02(256'h56A28D47481A358E2589A034A61058034C989A00D6C644D206B06080C66961E4),
    .INIT_03(256'h0B17440562F2AB5A4015BD852C2D77D20131D0A0018230E6194607D968029143),
    .INIT_04(256'h14028FF03C491FF8000888640896A80A3242257BDC00F977C2D2B7B8051AA450),
    .INIT_05(256'h28040908488FA0A8A1555F4BEFBD60243CC2020000DE702023BDE194800005A6),
    .INIT_06(256'h7D7C42A9446713E0402242501B533F8515947392605485F7D32D8400000458A0),
    .INIT_07(256'h2E54AAA2AA955E5AFC05502A8140AA4846A080457A90AA48848EE5FE6A822045),
    .INIT_08(256'hA85A294C8B414452B972AD10AFC8E7449E4210A8A5B5A9A2EE2A620544FD943A),
    .INIT_09(256'h233C1540D480F436D42C326AA851214CF18A49AB5CB44940B28F0C5202859226),
    .INIT_0A(256'h4C108411100C850240A58282494000142F7037481DA3833F202EB115B321EA30),
    .INIT_0B(256'h040A26511412E19508D6948400E0C07F107C65D76C800040043140080047FEC9),
    .INIT_0C(256'h3EC80C08957BBB6E62D51CA524100D9501557C6B26047F40882503A010C8604C),
    .INIT_0D(256'hECEF802CDC50BA289C0AA41220694710012D2BC00A5F584C92FFBE2B780851C1),
    .INIT_0E(256'hCA3809BE30E1840CD4D13E089E4A84173804BDCABA2FEF4819761007208961F4),
    .INIT_0F(256'h879BA2B14C21C4C0885475035424C87938A04A81102D0050278F3CA86720CE1C),
    .INIT_10(256'h507B470AC78BA96012200490209A541A6106043C9D1C3C9D10F2710F26887938),
    .INIT_11(256'hB2B324078491064B41400A829146282449D21B9C6D0FC91516ECA0055BACA101),
    .INIT_12(256'h1424204280F0891F70804C2A2810ACC44209965D9550A66BEC5440A2E603B54E),
    .INIT_13(256'h204811505BDA001205BAC005405E2501A0081239F05BB2291522933086143A04),
    .INIT_14(256'h2A056C209A6CF14CB542FA4134D85690269B5E6AA810A0025545520001249B2A),
    .INIT_15(256'hACFD4DE0114FC8498426150210B1C041051296010504C3F4045B902C8114F14F),
    .INIT_16(256'hD1C86C81005AA4EBD0410A2C49A0AA2BB6D0802804498ABB86EA0888001BB6F8),
    .INIT_17(256'h207802A8E30412A5F9090616C5E57BABF002ADD816FFC433DC2A6A540D57435D),
    .INIT_18(256'h7902C1376C4EBC88536095905D8533DA20D68A28203620B77764A9F69321C982),
    .INIT_19(256'hBA8A5022B7708AD80CC1103210CF2F2000A8435242CBA052840BA66E0E995606),
    .INIT_1A(256'h5444008D8000000000070060000000000000000DFBF94A5294F4F13D7C251C8B),
    .INIT_1B(256'h00000001E00000000000000000000000000000000000000000000040026E6E40),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_015 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n963,open_n964,addra[13]}),
    .dia({open_n968,open_n969,open_n970,open_n971,open_n972,open_n973,open_n974,dia[15],open_n975}),
    .wea(wea[1]),
    .doa({open_n990,open_n991,open_n992,open_n993,open_n994,open_n995,open_n996,open_n997,inst_doa_i0_015}));
  // address_offset=0;data_offset=16;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hF4BF7FFFB01D02A107C0503FFBD11C07BF4B565890FBEC66ED267C8BC1F5FCAE),
    .INIT_01(256'h8E4F4169B8D262B852E2240813F7FFE83848200BCDDA07FFAF19F77FDF7E3AEC),
    .INIT_02(256'h9D22DA5CB036A9DA3B6D60A8FEE8360A8EB6D522B6FD4DA315B7D102EED371E6),
    .INIT_03(256'hCB0677FBFBF2C35B3FA139902E2C621FFFD184DFFAA01824494C32CCCFFFF166),
    .INIT_04(256'h93FDCEE7BCB304507A31F9E7FF96E818B2420D739BE65C627FF42737F85AA685),
    .INIT_05(256'hB2B6B959553FB13132679E73CF3F7FC0FFECC1FFFFFEF8A63639DE14FFFFFD6F),
    .INIT_06(256'hFDFD7C28717FE0499F747EE4FE66FF061AE79FFA76DB3A55D170F28C95AEDE89),
    .INIT_07(256'h47863CFC33207ADCF99067833FFF0C87970F3D987CD70C872F3FFA166C3CAE01),
    .INIT_08(256'h47838E07AF560E832E246B578B59ABDFB262151B0898C71B5C4CAFBE613F483E),
    .INIT_09(256'hAB0A17FFE0D56D7FFE7A3882C196520DB182E20BFA8D92650CF6DF889C785E64),
    .INIT_0A(256'hD380000006FDBEF81F1EBA724913FFE2EF7BB79FFFA2C37F5FAAAA10A2B1E924),
    .INIT_0B(256'hF9536840907BE9A1A857A33BE0FFAE5EE665FBA2AC7FF0FFFEC53E0000756077),
    .INIT_0C(256'h785FEB72F7DDDD46D79E7FBDE6EFC56448707FFBBFFBFB7D2FFEFB00E01F4F0F),
    .INIT_0D(256'hFFF77EC1FFF0884F2FE37BFF890396C47E323FD7FA3FAFBA85F8CDCB77FE1D46),
    .INIT_0E(256'hDE78B7BCBFDCB97E56D67DFF827FB9A997B7EFF8E30FFF8264344FF3475FA15F),
    .INIT_0F(256'h77CF3C256C9DE1FB7E7067FF73A9F77C7FCACEB8780CFD068B2F7907BB1C8EF8),
    .INIT_10(256'h415B7A71397EEB2BBB7D7DA0AF0B5053BE3A93BE39E3BE39EEF8FEEF8EF77C7F),
    .INIT_11(256'hBBEB7506F49F2C5959F6FAB1DFFA19E5D3B2110C45CD8595F58CA37D5BDCA541),
    .INIT_12(256'h6582C841FFFE8858F2A290816FFFE8FC6CDB144D8D5B36DB5F9FEFBE43FB3586),
    .INIT_13(256'h4BCFA53E8A030E9C00053B6ABF919399E0231202019DE2A92020B11082048178),
    .INIT_14(256'h0A65852D1EAC7BCE914E4B5A3D59460A47ABF6A7ACF6A4C607C574D12124A9D6),
    .INIT_15(256'h1D10743FEF9E98C9846605AEE7E92EDE191A99FEC104FFF856D618ADFFFC7BC8),
    .INIT_16(256'hDBE3FD35792A90070FFAEA204008AA2A908CDF49E960AAA92225C12D3FD727C6),
    .INIT_17(256'h335A9EA423FE76E9D90A2602CDE169D3FA9EADE2FD9FE9AF4A1B6909F0F75109),
    .INIT_18(256'hDA2061A5481DBF89DB7295F94A9DB6ABF28B3BF137FAB2577C8C6DFE93E18B49),
    .INIT_19(256'hF30EB86966D1F977F02AE77210D62CFA89E7ED8ABED7F85AD1FB5DEA0B500BFF),
    .INIT_1A(256'h1505418F10000000001880600000001FFFE01E47EFF318C632FAFCBEFCE4BFDA),
    .INIT_1B(256'h00000606E000000000000000000000000000000000000000001FC00003B7C405),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_016 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1023,open_n1024,addra[13]}),
    .dia({open_n1028,open_n1029,open_n1030,open_n1031,open_n1032,open_n1033,open_n1034,dia[16],open_n1035}),
    .wea(wea[2]),
    .doa({open_n1050,open_n1051,open_n1052,open_n1053,open_n1054,open_n1055,open_n1056,open_n1057,inst_doa_i0_016}));
  // address_offset=0;data_offset=17;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h900D0061013C120C088054D000511C00034B56581000EC660126048800000200),
    .INIT_01(256'h8E4F45493A80AE002123361153F00000006C0408047A02ABE4100880107F9FB8),
    .INIT_02(256'h50A3A151400205CEE4282006E68B00006CC2828016C0C61600B40802C60B7160),
    .INIT_03(256'h0B064801EAF2834A00013980242C62100129D48001601864154402CCF00111C8),
    .INIT_04(256'h100197F502017FFFFFF03A040096E818324200739804FC6202D02730001AA400),
    .INIT_05(256'h28261909480FA03030061E03CF3C20003CE0000002DC70A202094019000005AE),
    .INIT_06(256'hF97D4038096707C808007601FA023F0038065992204005F5D120A0000424D880),
    .INIT_07(256'h82060C0003007F50FCE00000010800000C00020078380000240CE5FE4804A009),
    .INIT_08(256'h070A000C8B40040018304B508FC8EEC4AC63500800700002DC0CE69400FF973A),
    .INIT_09(256'h232A0240406A543EDE2FA0408010500481E081035834041010152C0860001224),
    .INIT_0A(256'h40000000000C840000000802490000002738230814A20111402AA2100231E820),
    .INIT_0B(256'h03E5D0B42D0AE1810857800000A0007E0072019AA00000000401000000756041),
    .INIT_0C(256'h1130100015FFFF6E53DC5DAD6620050030013FF800005E0008240300010E4008),
    .INIT_0D(256'hCFFE01063671D868180400020010022080203FA80AFFFFFE1FFFFFE3F00EE240),
    .INIT_0E(256'hDE7881BC2000808458802C00C00780019A40FFFFBC6DB9D88424000208212AA1),
    .INIT_0F(256'h078BC0012481C008007039017020007830804EA0382C0000030F7800033C8FFD),
    .INIT_10(256'h417BFA74868AB83E93653481BF9A5046C28C003C1E003C1E00F0600F07007830),
    .INIT_11(256'hB2FB644ECCB706CB79C27AB1F5D20BE4419A13AC0709933775DEE13D52DEE113),
    .INIT_12(256'h1474004080D88818E1AADC0808002DDC4E49B6DD857392FBCEDD72BEEB2397CE),
    .INIT_13(256'hCBEC03000BCFF17B87FFFB7F9FFF3DD9B6FFFFFB40DEF2291562B51082141200),
    .INIT_14(256'h2620246DAAE6CBDCB4C650DB55CB162E6AB9FEEFFCF6A4C255C576D02124AFFE),
    .INIT_15(256'h1CC016AB1518286A842205F60031E4C00112840005042C7D655B90288006CBDB),
    .INIT_16(256'h9B2BA409F97A905A4127AE22C40CAA3E908E880C80E0AAA93225402D155BB444),
    .INIT_17(256'h32529EA4213E5620CD0B36038CC8DBFB5A9EA9625DCD6D2F1A3929040DF5D1F4),
    .INIT_18(256'hD3280AB0085F9B89C937B779DF9C97FFF7FFABF9B2FEF2F65EECE4D996E0DBDD),
    .INIT_19(256'h3B8FFAEBF3F102203A1BFC2690FF3E7B8B809F5C02C3E052D00B046E0A590206),
    .INIT_1A(256'h454500CC10000004801D87E00000001FFFFFE067EFF318C632F2F0BCFC251CD4),
    .INIT_1B(256'h00000000E0000000000000000000000000000000000000001FC0000004187051),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_017 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1083,open_n1084,addra[13]}),
    .dia({open_n1088,open_n1089,open_n1090,open_n1091,open_n1092,open_n1093,open_n1094,dia[17],open_n1095}),
    .wea(wea[2]),
    .doa({open_n1110,open_n1111,open_n1112,open_n1113,open_n1114,open_n1115,open_n1116,open_n1117,inst_doa_i0_017}));
  // address_offset=0;data_offset=18;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h94BD006112052243102454F0007F9F7803EFF7DF9F00EFEE01BEC4CC01F5FEA0),
    .INIT_01(256'hBEDFE96D7FC163A88C1A6448BFF00008C308A20F47DEE2ABF88908881F7F9F7C),
    .INIT_02(256'h1A2A946B10E991CA228C9290A790EA290DA8C80A4FCAC542527CA90EF7A7F1FC),
    .INIT_03(256'h3FFE7E03F3F7CFFE8027FF917D3FE79F0145FD800202BEEEC3774FFFFC039555),
    .INIT_04(256'h3003AFF7B2533FFFFFC038BC0CF7FB7C77FFC7FFF80CFFE7E2D4FFF0099FFF9F),
    .INIT_05(256'hA0261904030FE30302619E53CF3D608F3CE4300002DC73F3433DFF1DC000253F),
    .INIT_06(256'h7D7F44E8616743C808B8F662FB673FA65FC7FB9268DC05F7FB29A4000424788E),
    .INIT_07(256'h0B9830B4F0219A7CFD91E00F01683C1807300081FCD03C18240FE5FEFE1EB210),
    .INIT_08(256'h881206448F4447110A4485578B48A356921A943A29510E3222422696603FD47B),
    .INIT_09(256'hFFFF17C0E444443EDEAE3888C91E2246F18AE2204EB60A3728644C10E8A99264),
    .INIT_0A(256'h4041086666FD86047F25820EDB13FF003FF07F0F1CEB373BC07EBB39FFBFEBB7),
    .INIT_0B(256'h0AB6B8F43D13F7E75FDFE62017E0817E407E63C7730008E004E181F27FFFFCE9),
    .INIT_0C(256'h37F8191097FFFF6ED7DE7FBDE6E03F827E4F7FFBA6207FFE0C7E03C8E5DEFF8E),
    .INIT_0D(256'hFFFF00087FF1FEEE0A1EA003C7E08BC13C2E3FF80EFFFFFE8DFFE3CBF018F2CC),
    .INIT_0E(256'hFFFF09FCF0C2988D73842C009D07905F9A44BFFFFE6FFFDACBAEC03248E9ABFF),
    .INIT_0F(256'h0FCBF0254F83F0C081F87F03F878C0FC3CC7FFFE3DEE0140870FF9A863FFDFFF),
    .INIT_10(256'h507BFB4C879EBA7E936576A7BF9B540FE1AE007E1F807E1F81F8781F87C0FC3C),
    .INIT_11(256'hBBF3644ECCB706DB69427A92FFFA0FE4D1DA13AC2F0BD33777FEE13D5BEEE113),
    .INIT_12(256'h8DFE86C080F9893FE1BEFCE77818ADDC4EDBB6DD8573B6FBCEDFFFBEEBF3B7CE),
    .INIT_13(256'hD86EA3729BCFF5FF87FAC01515FF3FC6BFFFFFD30430FE6D1522B7308E0CAC61),
    .INIT_14(256'h2E45A565BEEEF1DEB5CA5BCB7DDB56266FBB5E6AFE17E6CB57C7F7D221A48F42),
    .INIT_15(256'h19F79F31979FE88A84621D76C0B1C5D8670810013F844C74255B956F8116F1DB),
    .INIT_16(256'h9B2BA509B17AB1DFC1C7AE2FCDB6AA3FBEF6994DA8FF9BFB9FFFDF6F7FD36684),
    .INIT_17(256'h21521AA0A12C3668ED0B36378FECDBBBFA1AADD0BEFFE4BBFE3B6B040FF5DBF4),
    .INIT_18(256'hDB286BB5485FB9895337B739DF9533FF77FE9B79A5FEE2F776E4EDD99660DBDC),
    .INIT_19(256'hBB8FFAEBF7F1CB563A1BFC3690FF3E7B8BE07B5EBEF3E47ED18BC67E0FDD1F87),
    .INIT_1A(256'h1441110A00000005950C87E00000001FFFFFFF87EFF318C632FAFCBEFCA51CDE),
    .INIT_1B(256'h00000000E00000000000000000000000000000000000000000001C00012631C5),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_018 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1143,open_n1144,addra[13]}),
    .dia({open_n1148,open_n1149,open_n1150,open_n1151,open_n1152,open_n1153,open_n1154,dia[18],open_n1155}),
    .wea(wea[2]),
    .doa({open_n1170,open_n1171,open_n1172,open_n1173,open_n1174,open_n1175,open_n1176,open_n1177,inst_doa_i0_018}));
  // address_offset=0;data_offset=19;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h00080080013810AC0CC081000000000001000000000000000000040000000000),
    .INIT_01(256'h8000052800008C2025213211F00000001864060703A000000410000000420000),
    .INIT_02(256'hD5A32B54C0172C0CC569702E401B5602E0D69680B80546B405C0500080584100),
    .INIT_03(256'hC002000000608201000118800200200001B900C001E000001C0830000000118A),
    .INIT_04(256'hC80050084C80E001404987400082000080000811880200200050231040400000),
    .INIT_05(256'h1800000958008030300602204104124928402000004E235174000002000005C2),
    .INIT_06(256'h8C0400D01882844401C08243110702806721B51240C40042421050000004CA03),
    .INIT_07(256'h851E0CCCC301E7301961860C0F9430181C330E01882830181C0040126E3A0019),
    .INIT_08(256'h478808080800080230306E000480EFD2BE79C00000A08118FE0CC00401E84320),
    .INIT_09(256'h0000000040AA7032540990428098500AF06A410B1E820442149722081470C264),
    .INIT_0A(256'h00000000000000000000000000000000231001000780C0450008001000000000),
    .INIT_0B(256'h00000000000068000010000000000044000001B8AC0040000605000000240000),
    .INIT_0C(256'h0800000014000002000000000020004400108004000000000020000000010000),
    .INIT_0D(256'h08240107800400001400001208131424C21002000B6278C6650722C740000530),
    .INIT_0E(256'h02000084000080064CD03809424800001000A000809009291030000300010000),
    .INIT_0F(256'h0089000004004000181000011000000810884A00500000060921080002008800),
    .INIT_10(256'h086E2C844001410128180900064E021000416004080004080010200102000810),
    .INIT_11(256'h2037376D300B280E813CE000A106316D03228E5440DC0C80A81A5670000A55DA),
    .INIT_12(256'h14000150000008C052000008000032AE680C59579E9A026F31905097960DC927),
    .INIT_13(256'h27C001000C311039F8073FEEEA1151A00008003DF9DF8082A060111082141300),
    .INIT_14(256'h118008124006C04492328024800A11A510011310B9F000140540000D0159F9BF),
    .INIT_15(256'hEAC84244746028698426048803482A000112AC000024B3A9528408800006C040),
    .INIT_16(256'h40C0583434D0042050000A20000802000008C00800402000200140B080220D39),
    .INIT_17(256'h2CED380866ED92819144CA0064032632013800090008024000A00042000A0009),
    .INIT_18(256'h00400000022015CD01E880B645D0125168964966681129A4056680A601650122),
    .INIT_19(256'h200800000010028806C000081440000400980021020000000008000000000004),
    .INIT_1A(256'h10514018000000040408C67FFFFFFFE000000001221108421010100408240001),
    .INIT_1B(256'h00000404E0000000000000000000000000000000000000000000000306306904),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_019 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1203,open_n1204,addra[13]}),
    .dia({open_n1208,open_n1209,open_n1210,open_n1211,open_n1212,open_n1213,open_n1214,dia[19],open_n1215}),
    .wea(wea[2]),
    .doa({open_n1230,open_n1231,open_n1232,open_n1233,open_n1234,open_n1235,open_n1236,open_n1237,inst_doa_i0_019}));
  // address_offset=0;data_offset=20;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h5F4B006000220246806EA00E8013041101C95A4910504488008C840081201000),
    .INIT_01(256'hB31D359EE9225AE40289A0E01890001C02C1C000086044010000B2250C7E0CAA),
    .INIT_02(256'h3873B0C1400042EC061E04C00298614C00E1E0D30208760E98148201A08057B5),
    .INIT_03(256'hC04A01A26062C34180415A981440A000558339C00611280062A8C41B02585D88),
    .INIT_04(256'h20005C028240340CEE88380AB083018800960415A81300A011582B500048AE05),
    .INIT_05(256'h00E326809200C60000000200410590403970000002ECA0A3F81200002DB29552),
    .INIT_06(256'h0A06000000028040024803001002038001203F57B8642040594081F63E644FC4),
    .INIT_07(256'h0100000800001A1018E0000001840004040802000828000404004C1E4B22F000),
    .INIT_08(256'h0002002118080100000800430522A24EA2EC020410000000758D02C4012A5381),
    .INIT_09(256'h8808002C406A40B3578B900480180002E9FD40114F50000A0004B40400002A24),
    .INIT_0A(256'h80603000038110000010A008920002802B50051084D0007100484C5080D8ED40),
    .INIT_0B(256'h81C3C04010006B00509800001F0C017404011182A400061E8601000008642004),
    .INIT_0C(256'h2014C08316D111028E14300000201E000064C484891040002220000282A40001),
    .INIT_0D(256'h0C3700013300C00004D450020020010200001309AE671B38078DA70140005000),
    .INIT_0E(256'h834500844C00804464F83800690B0025D498F20882AA25890020201A02159400),
    .INIT_0F(256'h08ED004C8582E90000B000D1B041008E50C0CF1231F40102C10108A4B244CB18),
    .INIT_10(256'h9C4008880504FAC0A840F1008910271567F9E84728004728011CA011CA008E50),
    .INIT_11(256'h2D243846BC43009DFD35D139CFBA006C212A4DE4B81A3EF0282B53FDCD1B5610),
    .INIT_12(256'h2D35804800A01840693F50E7AD263FAD60CDFFE087F9B24158FBEFC77BF55F83),
    .INIT_13(256'h14E421008C7015B305F009C02A016CF317C06FD01130CC66BF225BB8E28C48C0),
    .INIT_14(256'h480B0003DBB64A44D9020607B768C845F6ED130DA93364D83D481594D5E589BA),
    .INIT_15(256'hDB905F85D0AC294DC73685CD801139B0091780001C14253B65AA18D4DE064A40),
    .INIT_16(256'h4207880467FB93DDBBB6BA668974524624B18848886F1962ABD9F7F2FA38D305),
    .INIT_17(256'hBF4DFEEE602FF6109526F27C0F1BAF1E29DEE28AE828AB88B6DA3920022FDE15),
    .INIT_18(256'hC7BC2FB890BDDDACD137F03FECCD12C177937D77B759EFF5A4C768D78862135E),
    .INIT_19(256'h211BE98AE0110A80080E2905926F86041093DA5E8210000D40484030012C0554),
    .INIT_1A(256'h041045BC10000001145940200000000000000001221738CE7010140409AC414C),
    .INIT_1B(256'h00000000E000000000000000000000000000000000000000202023C0030698E1),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_020 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1263,open_n1264,addra[13]}),
    .dia({open_n1268,open_n1269,open_n1270,open_n1271,open_n1272,open_n1273,open_n1274,dia[20],open_n1275}),
    .wea(wea[2]),
    .doa({open_n1290,open_n1291,open_n1292,open_n1293,open_n1294,open_n1295,open_n1296,open_n1297,inst_doa_i0_020}));
  // address_offset=0;data_offset=21;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h55640060002C02728037C00920120418008112691100448C0188800011200000),
    .INIT_01(256'h28183634C3824EA40A8F80C00C10001403C18040080065500000C3309C08128B),
    .INIT_02(256'h0019900100004006220606C4E098206C002060DB00405106D804000022003C15),
    .INIT_03(256'hC04A0143405C4188804052B894C0A0004840E0000603B844622C9613439008C4),
    .INIT_04(256'h200078400200711040083018C045018020960405281A00A008480A500062CC05),
    .INIT_05(256'hB8AF29011A02DA0000000200410580400960000002E8A0A3A038010016C31050),
    .INIT_06(256'h0A16800A000280401208030010020B90000004409864304959D002947CA03687),
    .INIT_07(256'h000100880000120010E0004001900086000C02000820008604104C1C00008000),
    .INIT_08(256'h02024001D168210800081F53870800082E0C100400204004710C320000049700),
    .INIT_09(256'h88082830026846834223840004004822546A1005459410020004980060000800),
    .INIT_0A(256'h004600222281000028028008920002000A50051003540C7080478C0094D80140),
    .INIT_0B(256'h40C0C14852005A02568C00001730012E00004123840004132220000008202002),
    .INIT_0C(256'h08160100020D1101C4840684206003003004620890106A022004008041450080),
    .INIT_0D(256'h40000003A3005400083040004000002002041B08C44C3B040918A20000004558),
    .INIT_0E(256'h21890084400080014F500401901D802490A05A184228A6085420001204100E19),
    .INIT_0F(256'h08E9000E8B83E88001F0C060F060808E104485D230F00102C30108A620804400),
    .INIT_10(256'h940E28D007055A86A9B08B818FBC250D7358604708004708011C2011C2008E10),
    .INIT_11(256'h0547CE61CD0A3044743F7BA85AE8015860684CA0B1F27CB1A94157BDC5415398),
    .INIT_12(256'h01EC000800E0150B4B175025AE4415293E44AA87026F918E29EEAD3529D446D3),
    .INIT_13(256'hB324001001AE15B1024816B0705550B30900121011004366F7828A006180A600),
    .INIT_14(256'h10A81008D3A00B2042150011A746112434E8085202C2049D5800C5EF18C13288),
    .INIT_15(256'hFA304928124B2155030188F8001122800213C0000C12A5B272EA0D74E8400B20),
    .INIT_16(256'h41845C0C6DFB921FFD20A04449BE9000A73A48040029D902E51ACEE0A88BF705),
    .INIT_17(256'h9D13DEEA0233A0303426D058F13B216C23DEE6A3A1408A8500BA3920062AD415),
    .INIT_18(256'h879C6BF052A58227D01531CE877D0C71953D53969D095BF0A8DAE811A3860857),
    .INIT_19(256'h92015B2AB80148C0E04C0B308229060416B9A84680210027F800801004FF8702),
    .INIT_1A(256'h015014B880000001C142C5600000000000000003A71738CE72525494AD8111C0),
    .INIT_1B(256'h00000000E0000000000000000000000000000000000000000000003FC58B5295),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_021 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1323,open_n1324,addra[13]}),
    .dia({open_n1328,open_n1329,open_n1330,open_n1331,open_n1332,open_n1333,open_n1334,dia[21],open_n1335}),
    .wea(wea[2]),
    .doa({open_n1350,open_n1351,open_n1352,open_n1353,open_n1354,open_n1355,open_n1356,open_n1357,inst_doa_i0_021}));
  // address_offset=0;data_offset=22;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h4616154BA8208252812DF001C0BE85A014B5BBCF1C0145C8059880640095D420),
    .INIT_01(256'h10100F3643007DF6489FE4E01E92AAB6232DC020A810977181441340856A0628),
    .INIT_02(256'h0033900908A0C04E2A0E04C5F0B8004C1420E0F3005059069805008B38002005),
    .INIT_03(256'hC0DE00024854A2988AC1D3D81443E0008141AD8AAE01386D608D9411432049F4),
    .INIT_04(256'h61544D43EE007191C87830AB006311A624B486BD38BA03E0004A1F5290454C07),
    .INIT_05(256'hA3A6BB40129B9A888100160A6925E848BB6200AAA7ECACF3A139200018E43170),
    .INIT_06(256'h58D4AA01044E2262960A270494076E89000110621C46365168C8EE9C3FB81E04),
    .INIT_07(256'h000002080894061292E01500A99302408482AB145A25024006284D5448908040),
    .INIT_08(256'h00428020A5580100040A10E32C09020E82049104840C2000712C30A000AC9734),
    .INIT_09(256'h9DC12C00804845A7762380202000000154EA00856194D1038004980292400200),
    .INIT_0A(256'h40C181511285002810A18A1ADB5004007E591D80045806018ADBCC04C8C85DC1),
    .INIT_0B(256'h0880C04812484EC2D1CA4088B7008B6EB4084183C62A9403C3130A02082C3200),
    .INIT_0C(256'h441001280200D102840400B4206546B0442C64D2A000AD81004429650086B040),
    .INIT_0D(256'h4FC42A4114E4E023A14600A620000000411017040DCF3BF8019CB78122A2E2D6),
    .INIT_0E(256'hA9ED14865085A10CE6D25452283B2026B1007816CE72A7CA8A28055200018E7E),
    .INIT_0F(256'h18E9002D8987F88125F84003F8D0818F10816F5536E055934103187040F677BC),
    .INIT_10(256'hDCD648D029BE3A81EA7D8F9189537738E3A720CF8800CF08033E2033C2018E10),
    .INIT_11(256'hAD6459448C1B2EC09D3DD1380510004961784944B1D3EAB1A9435EE88D435E51),
    .INIT_12(256'h647988C8557A902A5A1B7C43BF908A6D38C1550B0C8E32D70DF14AA450A508AF),
    .INIT_13(256'hF3E07419C83555F7135B36B2FFD56CF30D64DAD851306B64F5029102B2806ED4),
    .INIT_14(256'h1A990420D9EA8B28C3534241B3D05304367AA29282F1ACDF5940FD95189F38C8),
    .INIT_15(256'h6339DD081643214815A081959459F235191280AC5F903563416F80B6F192CB48),
    .INIT_16(256'h53EC7C044A61312BF0C7204B59BEB801EF7A84C09D7AD91EE518CC4316BAD304),
    .INIT_17(256'hAA1E744E205944B43C24A258F9F2A5FEAE7442A0494AA10D2362130157F1D40F),
    .INIT_18(256'hC7782F741ABBAFAB116A31E54B310EB2EA8E22E5224094C1AC99889183C5D82A),
    .INIT_19(256'h3A873B26CFF0DD7C86099C17F2748A0F9EB7611C96D1E8DC4C0348BE1B8CC501),
    .INIT_1A(256'h1114448190000005C057C7E00000000000000001621738CE701014041985D972),
    .INIT_1B(256'h00000606E00000000000000000000000000000000000000000C0C00006B93E4C),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_022 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1383,open_n1384,addra[13]}),
    .dia({open_n1388,open_n1389,open_n1390,open_n1391,open_n1392,open_n1393,open_n1394,dia[22],open_n1395}),
    .wea(wea[2]),
    .doa({open_n1410,open_n1411,open_n1412,open_n1413,open_n1414,open_n1415,open_n1416,open_n1417,inst_doa_i0_022}));
  // address_offset=0;data_offset=23;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h5F560C5A882082424324F0041196C7BA0DA5BBEF1D616788459892651125048A),
    .INIT_01(256'h30183526439A4EE208CB90601CE2667C2260C0608804F7D11144E4069C2816A9),
    .INIT_02(256'h081BC00128C04056300606C068D8A06C038061DB00685407D806808CB8807416),
    .INIT_03(256'hC1EB2033485CA38C99D0FFBC95C6B1882400A5099C01BA68608DC411400E0DF0),
    .INIT_04(256'h60CC4D43CA083191CE28300C22C3118624F6A40FF87B12B105481AF234664D45),
    .INIT_05(256'hA3A639981232B28001004200E38DED40F960C0998EF9A5F3A03801001F08D0F1),
    .INIT_06(256'h1A9DBA020402A0E2520E03801402CEC9020005709D443A41CDD4829D3CA1FE8E),
    .INIT_07(256'h200182080010121238E4004001918286400C02440A2182868600CC5604018044),
    .INIT_08(256'h2002C0039DCA214884020FD2841822492E0C908584286084748C298104249782),
    .INIT_09(256'h88812846C278C4C742238420244008275CFF180584DC1003800C994292042822),
    .INIT_0A(256'hC1D1A8222285A2187009E23EDA540640FAF19794435C140189DACC1084C84DC1),
    .INIT_0B(256'h20C0814852404ED2F7CA4118760A872EA608D3E1E52634881720860A88282C18),
    .INIT_0C(256'h5211417046001D0284000085A064D6304426E6D88181EC03212419A180062081),
    .INIT_0D(256'h468018E13784C8412009118E6000403083001302264E3A180595A7010273E002),
    .INIT_0E(256'hA3CD878E5A8CA52FCED35CC7DAFFA9A5B0125A188E2AA788806004D601048E78),
    .INIT_0F(256'h38E9082F8B8FF8A027F8401BF9E0A38E12070DDA39F44D8343810CF951E6FF3D),
    .INIT_10(256'hFE96C8D027EEBE90A27DBFB1D95F7FB0EBA1E1C70841C708473C2473C2238E12),
    .INIT_11(256'h8D6459408E3B2EC09E3FFBFD9552164DF05E4940B3D3EA3BA94B57FDED535E51),
    .INIT_12(256'h687F68884CF6902A6ADB781BB8132AE97EC9554B088FB2D70DF54A2652A409AF),
    .INIT_13(256'hF0AD557D09BF55F7135336A2AFD518F38D6CDA9C5D506F6075239110B0C85398),
    .INIT_14(256'h9AA90428DBA6CA6843574251B746532436E9B8D02A35E45F5802D57F198D93C8),
    .INIT_15(256'hFB39DB8C142F214001A2CDDF3459BFE71B128098DE9435225B6F07B68526CA48),
    .INIT_16(256'h13EDFD06CB7BFB29F09EAA6BC8FEBE16ABFA5EA5D13ED86A670F37E7BE8AD14C),
    .INIT_17(256'hCA5CFEFF40DD46F82F24A05979F285FCACFEF6A9494AB10D227A3FA13F75F485),
    .INIT_18(256'hC7786FF05AAD9FAAD06ABBF509AD1496CA0422C50A4096F5A88DE891C7C5D92B),
    .INIT_19(256'h9687BF3A7B93D8B0C6491B13F23E0E0E9E9F611CA4E1B8F7F82B81FA0EFF8763),
    .INIT_1A(256'h1415044480000000405D40600000000000000003E737BCEF7A535CDEAD815150),
    .INIT_1B(256'h00000000E0000000000000000000000000000000000000000000000007CBCA70),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_023 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1443,open_n1444,addra[13]}),
    .dia({open_n1448,open_n1449,open_n1450,open_n1451,open_n1452,open_n1453,open_n1454,dia[23],open_n1455}),
    .wea(wea[2]),
    .doa({open_n1470,open_n1471,open_n1472,open_n1473,open_n1474,open_n1475,open_n1476,open_n1477,inst_doa_i0_023}));
  // address_offset=0;data_offset=24;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h20087C25680C012040008009EA284204A01081040889501108C12A20080E014F),
    .INIT_01(256'h0000000080116C5042418F040021E1FE217A0020800110001144F77002C82B5C),
    .INIT_02(256'h0818D0692820C0181A0206459860A06417A0A13900380D03C8038C0288844102),
    .INIT_03(256'hD42421424800E21407C00908045010C8C8400217860384002000C00003B0EC24),
    .INIT_04(256'hE03C12BC0A000E6F39A801EBCC200222010A009202104C11082A0501B0018442),
    .INIT_05(256'h180010011A910A0080004500A088886802088187818408048000002027EF0830),
    .INIT_06(256'h02000809000C20A0C40800042000400900000000808002828100200068044A01),
    .INIT_07(256'h404080860094101020680000800B8040C0808140101180408230100608804040),
    .INIT_08(256'h020201011C0101C081081083009002472F040081802C208505801308000823B4),
    .INIT_09(256'h1048003040244030A109C220A05141068875008047410102024C004004002C02),
    .INIT_0A(256'h5204840100000A8208A2904049500020E509824408100A630785440418520440),
    .INIT_0B(256'h508080088220109000120081E0100E0482000202245E0413EC0120020020200A),
    .INIT_0C(256'h09863A00200001CC000000001C2C000103001920B41980001020802040400010),
    .INIT_0D(256'h388078030C0062028970C86E2008400201410504CE34A60002E2CA000602F285),
    .INIT_0E(256'h0200A008118D8004D00001C020000006B1A1E5F08E877B8BCBE003C204110466),
    .INIT_0F(256'h41380408A010CC1146340061321414030161000902003C20E000100640000800),
    .INIT_10(256'hE4CA38D019752C860180802086E37932F3B62201002201802826028060140301),
    .INIT_11(256'h8563EF21C60F100184700148841201F8B80C404090F22219E9415800A54153C9),
    .INIT_12(256'h01838008432E100090095442AFC4A2B9500041450194018B2BA142BE10251974),
    .INIT_13(256'h1C0861218065F0CEEFFDFFFFF07F030D3B97B76BE9205930200110102080ADC4),
    .INIT_14(256'h00180003D1EAC0E0C0010007A3D01003747B121CAF0100240D0000011008008C),
    .INIT_15(256'h45CFD973F590E908050284238011407101000086C5142051012A8094F8D280C0),
    .INIT_16(256'h0C04010C368160A9BCC5224200081600000890C91C224C002100C41B57C9ACB5),
    .INIT_17(256'hA20D005202284E5C072022486D108534A90052A44942A50D03C11600F2A96430),
    .INIT_18(256'h0094257400B3BDAE092299A10DE096D162B4AB4122428D00AC6B04B8C3420008),
    .INIT_19(256'h00892D00038222200CA3380102240895149467B9801440084C185014110C8108),
    .INIT_1A(256'h154005BB90000001C057C0600000001FFFE01E504024A42949282A4811040208),
    .INIT_1B(256'h00080202FFFC000000000000000000077FFFFFFF80000000001FC00002817F08),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_024 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1503,open_n1504,addra[13]}),
    .dia({open_n1508,open_n1509,open_n1510,open_n1511,open_n1512,open_n1513,open_n1514,dia[24],open_n1515}),
    .wea(wea[3]),
    .doa({open_n1530,open_n1531,open_n1532,open_n1533,open_n1534,open_n1535,open_n1536,open_n1537,inst_doa_i0_024}));
  // address_offset=0;data_offset=25;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h3248431C40000308400020063386C1C73CA4308206F24388AC3836219305028A),
    .INIT_01(256'h0022136B80127C524240B62C00201FFE20605020400015540200117702A807FE),
    .INIT_02(256'h1830D001202041101A0604C1186000C412A061B104309903980308812C820103),
    .INIT_03(256'hC001000AC8804200204000080468D000030102907E0900006040804000CC1820),
    .INIT_04(256'hE20018000A1920010628100801000812020060C28010200000BC292408100480),
    .INIT_05(256'h3422110416A032810110010880028460300C807F801500068100A19003EE3D70),
    .INIT_06(256'h17001600001820A196080C44070484010000400280033D00040C840128200640),
    .INIT_07(256'h6240008E0894041008680180B01B82C6848C315C063782C68BB0A80448804040),
    .INIT_08(256'h20024104988805418402000C6048A000130410048000200280A0130604003380),
    .INIT_09(256'h100382015064C0049509C4000050010608F7A0060AC040020044000200041024),
    .INIT_0A(256'h10000411000188004221D00E92404022202A06002010300410082C3808410143),
    .INIT_0B(256'h1A84800C023800810083200200810E04100190402441BC0C3491803000B42000),
    .INIT_0C(256'h0003C0082800010200088000102BC00100014050998200C208C00062301090C8),
    .INIT_0D(256'h868C46C11602004080A112002140421342380580142130201300820245E24001),
    .INIT_0E(256'h220101281190801C4004293624004444B432F0000AA000080020080640030460),
    .INIT_0F(256'h01380408C400E81A003400043008100201810008080880006200040048008801),
    .INIT_10(256'h3481011100040C8010020062A0008D2003003001102009002024020044101221),
    .INIT_11(256'h6F00201C060000380400064880060004C80C4018B402601806D9600325096807),
    .INIT_12(256'h8102A1483F061000A0019000CBE720810038000010100E400070400200090100),
    .INIT_13(256'h700E102240A0109502432486E10112A10F0C9E184160413064231000A0840140),
    .INIT_14(256'h109C035241A6C026E21B02848340058410699810AA300204A0440200190C8802),
    .INIT_15(256'h4A1044A4112C294801229002918100500100807EC014201000220010BEE40100),
    .INIT_16(256'h801083150004E100B000624004094E201004990124204C012020000000089504),
    .INIT_17(256'h80C00112A500004007200E5A05300006E40196D012D8D0610000C62800207400),
    .INIT_18(256'h4044207000E190A806209800008060000080000040800009E0040300C0200702),
    .INIT_19(256'h20890D400011028001920001226010001480208080100000441840000018400C),
    .INIT_1A(256'h400004C5800000004057C0600000001FFFFFE060042430884020040803241018),
    .INIT_1B(256'h00000202E000000000000000000000007FFFFFFF800000001FC0000000A977F7),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_025 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1563,open_n1564,addra[13]}),
    .dia({open_n1568,open_n1569,open_n1570,open_n1571,open_n1572,open_n1573,open_n1574,dia[25],open_n1575}),
    .wea(wea[3]),
    .doa({open_n1590,open_n1591,open_n1592,open_n1593,open_n1594,open_n1595,open_n1596,open_n1597,inst_doa_i0_025}));
  // address_offset=0;data_offset=26;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h300000010800005880098000083EC37880A4A1860F084B8820B88C0181050088),
    .INIT_01(256'h2000061D00017E46000392C01C23FFF4004580406006E0004004F777006A062A),
    .INIT_02(256'h0033902118C0C00C000A0CC00490A0440100A011040885068800880D00000041),
    .INIT_03(256'hCA0D000AC8A02000004020582468D00003008C00040100006320800200003980),
    .INIT_04(256'hE00108000A1020010028000801808000000202021014808000A8040008000440),
    .INIT_05(256'h42001100128102008010010022888340E08000FF800044008400000007EE0872),
    .INIT_06(256'h1009640104010002000800702100042804000010000000A00300800028044260),
    .INIT_07(256'h2041000808040012287000200010824040800000162082400880000648800004),
    .INIT_08(256'h2002600001480501810200442008004083040080800020848000088504200328),
    .INIT_09(256'h406212011020443494098200A050000690E00806088001028004000000241006),
    .INIT_0A(256'h1010841100748C024020DA020150402009202200243000014028040464400840),
    .INIT_0B(256'h12848008022020800042100001010EC4514190C004000480089180CA00B42400),
    .INIT_0C(256'h000020082000010200000000102000100005C0008008000080A0002100104000),
    .INIT_0D(256'h06A80021160000008800080000004012010001001E003000110000020002C041),
    .INIT_0E(256'h2000000211808414C20008000C000004B00150002A2000080020000600038460),
    .INIT_0F(256'h012804088600CC1000300005305010132101080920080010E20000004A008800),
    .INIT_10(256'h5580031400040E80000100328000513003003009902001102026020244100301),
    .INIT_11(256'h0D80008C068101100400000A01062820890C5014B002611812C160004589C023),
    .INIT_12(256'h8102810900001800A0039001C800600541180040841044400030408002090000),
    .INIT_13(256'hD00C00204168100002400780610100010F001200010041313120210022840144),
    .INIT_14(256'h2C49890541A6D030518B8B8A834955801068AAD02A1000002444000038083706),
    .INIT_15(256'h00004000100021088502840291810051011081000010600000620018800E4811),
    .INIT_16(256'h000801940002A320B000686000004020000498210420CC006000000000080004),
    .INIT_17(256'hA080008AA10010448728085805304004F40087940249C0632004684000207400),
    .INIT_18(256'h4800207100A1802023209810008222082000082060802001B0001180D0202200),
    .INIT_19(256'h00810F080003028010820000E220000014C0208082100000C51040000018008C),
    .INIT_1A(256'h0000059680000000405540600000001FFFFFFF824424A42D6800200801A01018),
    .INIT_1B(256'h00000000E000000000000000000000007FFFFFFF8000000000000C0005FC2AA8),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_026 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1623,open_n1624,addra[13]}),
    .dia({open_n1628,open_n1629,open_n1630,open_n1631,open_n1632,open_n1633,open_n1634,dia[26],open_n1635}),
    .wea(wea[3]),
    .doa({open_n1650,open_n1651,open_n1652,open_n1653,open_n1654,open_n1655,open_n1656,open_n1657,inst_doa_i0_026}));
  // address_offset=0;data_offset=27;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h200800000000800000008000083E837881A4A1864F084B8820B88E66530500A8),
    .INIT_01(256'h8000000000084E400003800410240014004010606002000000440000406A0628),
    .INIT_02(256'h083380090020C1040006044000102044008060130408950288200102A4804140),
    .INIT_03(256'hCA0C000AC0808000006168082C40100002400000040300002108800000003880),
    .INIT_04(256'hE00018000A0960010028200C0180200010022016801020400038040000000480),
    .INIT_05(256'h012611041281028001104400A2088260040001006C040402800000800011C570),
    .INIT_06(256'h0001420300001002000A04702304040004100000018000800300800028004260),
    .INIT_07(256'h20408088088400100874006000900200000080C0122002008000802408810200),
    .INIT_08(256'h2002010090480500890200442000224082165084800400000020001204280300),
    .INIT_09(256'h002200015020400014098000A040000290E2A00400004102000C000002001026),
    .INIT_0A(256'h5000000010000C0200809202410000202D280240349008050008040400410840),
    .INIT_0B(256'h1284800802200090085310000001204440200880240004000C10000000252000),
    .INIT_0C(256'h000020003400010200000000102000110000C0008008000000A0020010000000),
    .INIT_0D(256'h0E880001160100408800080200080000000901001E2030000300000040024001),
    .INIT_0E(256'h2200810A118180104280200008001454B001F0000AA000080020000220038460),
    .INIT_0F(256'h002A040AA400CC18003000053000100201430A2920000040E00294A048000020),
    .INIT_10(256'h0581033400040C8000000030A000111003003009902001002004420264100301),
    .INIT_11(256'h25A0200806810018150000A880020804C00E500CB402211814D3E0010DA94003),
    .INIT_12(256'h1102A14800001880800190018800400140101040900006000060008200010000),
    .INIT_13(256'h108C11304828100003C00780608100010F001200017041307400200020800140),
    .INIT_14(256'h2C48080041A41976F18B8000834955801068B8500A30200034000000190C3400),
    .INIT_15(256'h00004000100021488502800291210050201200000014600000320010800ED951),
    .INIT_16(256'h0000018500008220B0006260400068000000102104204C006000000000080004),
    .INIT_17(256'hA0C00022200002600628025A0510400E240003C402CAC0514100482000206400),
    .INIT_18(256'h4800207100A1802802801C10000032082080082040200005B4040100D0200302),
    .INIT_19(256'h20810D40001302800082000072E000001C80208082100000401840000008000C),
    .INIT_1A(256'h800004F810000001C057407FFFFFFFE000000002442420084000000011201018),
    .INIT_1B(256'h00000000E000000000000000000000007FFFFFFF800000000000000102020020),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_027 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1683,open_n1684,addra[13]}),
    .dia({open_n1688,open_n1689,open_n1690,open_n1691,open_n1692,open_n1693,open_n1694,dia[27],open_n1695}),
    .wea(wea[3]),
    .doa({open_n1710,open_n1711,open_n1712,open_n1713,open_n1714,open_n1715,open_n1716,open_n1717,inst_doa_i0_027}));
  // address_offset=0;data_offset=28;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h200800000000000040008000083E837881A4A1864F081B9920F98C44410500A8),
    .INIT_01(256'h80000160000044420000A40000200014006410202002000044000000406A0628),
    .INIT_02(256'h083380010000400C020E04C000102044008020110000840698208080A4804140),
    .INIT_03(256'h0005000AC020C2000061490C0440404003410080040100002000800000003880),
    .INIT_04(256'hE00018000A0060010028000C01824800000220168010000000BC292004000440),
    .INIT_05(256'h0002110012800208000041082000826034800000000404208000000000000D72),
    .INIT_06(256'h1300020004010022400A0160030404000400110280008000840400102C044240),
    .INIT_07(256'h0040000A000000020A6000608210024004000044162080008080202408810200),
    .INIT_08(256'h0042010009000500010200002008804002040080800400020000009504200328),
    .INIT_09(256'h000282015060C000000BA600800101029262A08400004002820C000202000024),
    .INIT_0A(256'h500000000000880000809000014000202D2802402490000100002C1020400040),
    .INIT_0B(256'h128480080228A090005310800001004440000880240004000C91000800242200),
    .INIT_0C(256'h000020003400000200000002102000010000C0008008000000A0020000000040),
    .INIT_0D(256'h0EAC0021160000000000080220004010010105001420300003000000400A4001),
    .INIT_0E(256'h2200800211C08414C280280008000004B001F0008AA000080060000620038460),
    .INIT_0F(256'h002804080400CC10003001053004100301C34A2900000040428210004A008820),
    .INIT_10(256'h4441051000040C80000010328000513003003001802009102024420244100201),
    .INIT_11(256'h0D80000C068100101400022A01040000818E5004B402211812DB680047894803),
    .INIT_12(256'h850280480000188000011001C8006085001810009000064000200080060A0100),
    .INIT_13(256'hD00C002008201000024004806181000109001E00011041317000200020800140),
    .INIT_14(256'h2C48080041A6D976F18B8000834955801069BAD0A21020003100000018083B04),
    .INIT_15(256'h00004000100021088502800290010050250280000014604000320018800ED951),
    .INIT_16(256'h0000811400028320B000604040006A00000010098020CC002000000000080004),
    .INIT_17(256'h8000008280040044C728065A05104004B00022C01648D01101004A4000206400),
    .INIT_18(256'h4800207100A190A003209C10400032000082080060902000B0000180D0200202),
    .INIT_19(256'h20810D000001028010920000D2E020001480208082100000441840000008000C),
    .INIT_1A(256'h000005E280000001405D406000000000000000000006308C6020200810041018),
    .INIT_1B(256'h00000202E000000000000000000000007FFFFFFF80000000202033C0020A0220),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_028 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1743,open_n1744,addra[13]}),
    .dia({open_n1748,open_n1749,open_n1750,open_n1751,open_n1752,open_n1753,open_n1754,dia[28],open_n1755}),
    .wea(wea[3]),
    .doa({open_n1770,open_n1771,open_n1772,open_n1773,open_n1774,open_n1775,open_n1776,open_n1777,inst_doa_i0_028}));
  // address_offset=0;data_offset=29;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h200800000800800000008000083EC37881A4A1864F081B9920F98E444111028A),
    .INIT_01(256'h80000169000044420000B6001020001E006400000002000000400000406A0628),
    .INIT_02(256'h183390490820C004020E04C00010204400806011040084068820000204004140),
    .INIT_03(256'h0001000AC8A0C200007169080440400003410080040100002000800000003884),
    .INIT_04(256'hE00018000A00600100280008018248001802001680100010003C290000000400),
    .INIT_05(256'h0000100012810280001004088208806034800000000400208000008000000D72),
    .INIT_06(256'h0308020104041082000804002A14040004101112800000000304000028044A40),
    .INIT_07(256'h0000820A00040410286000208210000044808280102002400000000640810240),
    .INIT_08(256'h0002000009010540010200002008A24082040080000420000020000604280300),
    .INIT_09(256'h000200014060C0349009A400A05101021062A804080041028204004202041024),
    .INIT_0A(256'h101084000004880000009A00010000202D2002002490080500082C1420401040),
    .INIT_0B(256'h128480080220A080005380800001004450000880240004000C81000800242200),
    .INIT_0C(256'h000020003400000200000002102000100100C0008008000080A0022010000040),
    .INIT_0D(256'h0EAC0001160000000000080200080002000101001E2030000300000040024001),
    .INIT_0E(256'h2200010811808014C2802800080000049001F0008AA000080060000620038460),
    .INIT_0F(256'h013A04080400C810003400053004100301C34A2900000040400000004A008820),
    .INIT_10(256'h0440003000040EA000001022A000114003003001802001002004020040101221),
    .INIT_11(256'h2720200C06000018050002A881060800890C5000940A201812CBE8004DA36003),
    .INIT_12(256'h8502804800001800200110008800600100181000901004000020000000000000),
    .INIT_13(256'h108C002001E0100003C00780200100010F001E000170C33175203110A2840140),
    .INIT_14(256'h2C48080041A6D976F18B8000834955801069AA9002202000304000001808BA02),
    .INIT_15(256'h00004000100029400120840281210051210200000014205000220030800ED951),
    .INIT_16(256'h000081150000A400B0006A6040006A000000102104204C002000000000080004),
    .INIT_17(256'hA0C000AA210400408628004A01100006E40026D0025280030000420000207500),
    .INIT_18(256'h4800207100A1802003209C10008020000000000000000004E4040180C0000300),
    .INIT_19(256'h20890F40001102800082000052E000001480208082100000441840000008000C),
    .INIT_1A(256'hA00005AA80000001C055C0600000000000000000000420084020200810241018),
    .INIT_1B(256'h00000000E000000000000000000000007FFFFFFF800000000000003FC202A28A),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_029 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1803,open_n1804,addra[13]}),
    .dia({open_n1808,open_n1809,open_n1810,open_n1811,open_n1812,open_n1813,open_n1814,dia[29],open_n1815}),
    .wea(wea[3]),
    .doa({open_n1830,open_n1831,open_n1832,open_n1833,open_n1834,open_n1835,open_n1836,open_n1837,inst_doa_i0_029}));
  // address_offset=0;data_offset=30;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h210800200804800000008000083EC37881A4A1864F081B9920F98E444115028A),
    .INIT_01(256'h80000169000844400020A40410200016004010202000000000000000506A1628),
    .INIT_02(256'h083380410800400E20060440A018004C00A0E0530408850698208000A0815140),
    .INIT_03(256'h0000000BC8A0C2000061480804401040034100800401104020048000000039C0),
    .INIT_04(256'hE00018B08A0862C14028000801824882000200168010000000BC290000000401),
    .INIT_05(256'h900010011A000208810041002080104024020000009440208080000000000D72),
    .INIT_06(256'h100942010404108200080400220504400500111280000000200400002805DA61),
    .INIT_07(256'h000000080890001208741000001082404480824402208240888080264A810240),
    .INIT_08(256'h20C221000901014080000110A008A242AA040000042400807000220600280328),
    .INIT_09(256'h8802000140684430140BA400801000029062A00408000002000C000000000022),
    .INIT_0A(256'h501084000004880200009202484000202D2802002690084500082C1020400040),
    .INIT_0B(256'h128480080228A080001310800001004440800880240004000C91000000242200),
    .INIT_0C(256'h000020083400000200000042102000110100C0008008000080A0020000000040),
    .INIT_0D(256'h4EAC0001160400000004080220204010000405001E2030000300000040024000),
    .INIT_0E(256'h2200800211818015C080280080008004B001F1208AA164080060000620038460),
    .INIT_0F(256'h012A04080400C810003000053000100201C74AB800040050400004004A008820),
    .INIT_10(256'h14575E1000040C80000520B08B01450803003009902009102024420244101221),
    .INIT_11(256'hA50501080681021815000809810622E4C1CE5014940A2118044944050719C042),
    .INIT_12(256'h0406A2480000180002211080880040814210000B041086170070402E02090100),
    .INIT_13(256'h10C80130082010020240148016010041090052000110C3B055229110A284C344),
    .INIT_14(256'h2C48080041A6D976F18B8000834955801068B850AA20200475000001790CBF06),
    .INIT_15(256'h000040001000294885228586802130D0011200000014204004221010800ED951),
    .INIT_16(256'h00290584580A2080B00068404008E000000A982984606C000000000000080004),
    .INIT_17(256'hA0C00202645C1260E7280A4A0510400622028388144980610008600000206400),
    .INIT_18(256'h0D8C243100A19028428018000B8430B2E02E02E060902014A0A02100D0204302),
    .INIT_19(256'h20890F4000110A80028A000652E000001580208082100002581840000049C50C),
    .INIT_1A(256'hD55551FD100000019508806000000000000000024426308C6222208890241058),
    .INIT_1B(256'h00000202E000000000000000000000007FFFFFFF8000000000C0C00007DFF55D),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_030 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1863,open_n1864,addra[13]}),
    .dia({open_n1868,open_n1869,open_n1870,open_n1871,open_n1872,open_n1873,open_n1874,dia[30],open_n1875}),
    .wea(wea[3]),
    .doa({open_n1890,open_n1891,open_n1892,open_n1893,open_n1894,open_n1895,open_n1896,open_n1897,inst_doa_i0_030}));
  // address_offset=0;data_offset=31;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h200800000800800000008800083EC37881A4A1864F081B9920F98E44410100AA),
    .INIT_01(256'h80000169000844420000B60410200014006410202002000000440000406A0628),
    .INIT_02(256'h183390490020C00C020E04C00010204C00A0E0130408050698208880A0804140),
    .INIT_03(256'h0001000AC820C200006148080440104003410080040100002000800000003984),
    .INIT_04(256'hE00018000A00600100280008018248020002201680100010003C290004000440),
    .INIT_05(256'h000010001281028881104508A208100034820000009440000080008000000D72),
    .INIT_06(256'h0000000404000022400A00100210000004101112808000808000000028044A60),
    .INIT_07(256'h0000000A00040010087010000010800004000204002080008080000648000004),
    .INIT_08(256'h20C2410009010140000000002008A24082000000000400000000000600280328),
    .INIT_09(256'h000200015060C434940BA400A05101029062A00408004002000C000202000226),
    .INIT_0A(256'h50108400000488000000920000000020290800002490080500082C1020400040),
    .INIT_0B(256'h1284800802282080005310800001004440000A80240004000C91000000242200),
    .INIT_0C(256'h000020083400000200000042102000110100C0008008000080A0022010000040),
    .INIT_0D(256'h0EAC0021160000008000080220084010010105001E2030000300000040024001),
    .INIT_0E(256'h220001081180801442812800080004009001F0008AA000080020000220038460),
    .INIT_0F(256'h002804080400C810003000053000101321C34A2820000040420210004A008820),
    .INIT_10(256'h0040000000000C00000000208000000000003001002001802006020060100301),
    .INIT_11(256'h2120200C068100181100000081062024C18E1004040801180008400001084002),
    .INIT_12(256'h0402A04000000840802000800000608440181040941006410050408202090100),
    .INIT_13(256'h10CC113048201000024004800001000109001200011082305520111082044144),
    .INIT_14(256'h2C4808000026D976F18B8000004955800009BAD0AA30200035400000790CBF06),
    .INIT_15(256'h00004000100028488422050280201050010200000004004004001000000ED951),
    .INIT_16(256'h000001840000000000006A2040006A000000982984400C000000000000080004),
    .INIT_17(256'h20C0000024041264C70802020400400220000080000880000400400000006000),
    .INIT_18(256'h480030110001908803A09C1040803200208208206090200424040180D0200302),
    .INIT_19(256'h20880E40001102800082000050C000000080208082100000001840000000000C),
    .INIT_1A(256'h8000002A000000000002002000000000000000024426308C6000000000241018),
    .INIT_1B(256'h00000000E000000000000000000000007FFFFFFF80000000000000000088080A),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_000000_031 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1923,open_n1924,addra[13]}),
    .dia({open_n1928,open_n1929,open_n1930,open_n1931,open_n1932,open_n1933,open_n1934,dia[31],open_n1935}),
    .wea(wea[3]),
    .doa({open_n1950,open_n1951,open_n1952,open_n1953,open_n1954,open_n1955,open_n1956,open_n1957,inst_doa_i0_031}));
  // address_offset=8192;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_000 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n1983,open_n1984,addra[13]}),
    .dia({open_n1988,open_n1989,open_n1990,open_n1991,open_n1992,open_n1993,open_n1994,dia[0],open_n1995}),
    .wea(wea[0]),
    .doa({open_n2010,open_n2011,open_n2012,open_n2013,open_n2014,open_n2015,open_n2016,open_n2017,inst_doa_i1_000}));
  // address_offset=8192;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_001 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2043,open_n2044,addra[13]}),
    .dia({open_n2048,open_n2049,open_n2050,open_n2051,open_n2052,open_n2053,open_n2054,dia[1],open_n2055}),
    .wea(wea[0]),
    .doa({open_n2070,open_n2071,open_n2072,open_n2073,open_n2074,open_n2075,open_n2076,open_n2077,inst_doa_i1_001}));
  // address_offset=8192;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_002 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2103,open_n2104,addra[13]}),
    .dia({open_n2108,open_n2109,open_n2110,open_n2111,open_n2112,open_n2113,open_n2114,dia[2],open_n2115}),
    .wea(wea[0]),
    .doa({open_n2130,open_n2131,open_n2132,open_n2133,open_n2134,open_n2135,open_n2136,open_n2137,inst_doa_i1_002}));
  // address_offset=8192;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_003 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2163,open_n2164,addra[13]}),
    .dia({open_n2168,open_n2169,open_n2170,open_n2171,open_n2172,open_n2173,open_n2174,dia[3],open_n2175}),
    .wea(wea[0]),
    .doa({open_n2190,open_n2191,open_n2192,open_n2193,open_n2194,open_n2195,open_n2196,open_n2197,inst_doa_i1_003}));
  // address_offset=8192;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_004 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2223,open_n2224,addra[13]}),
    .dia({open_n2228,open_n2229,open_n2230,open_n2231,open_n2232,open_n2233,open_n2234,dia[4],open_n2235}),
    .wea(wea[0]),
    .doa({open_n2250,open_n2251,open_n2252,open_n2253,open_n2254,open_n2255,open_n2256,open_n2257,inst_doa_i1_004}));
  // address_offset=8192;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_005 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2283,open_n2284,addra[13]}),
    .dia({open_n2288,open_n2289,open_n2290,open_n2291,open_n2292,open_n2293,open_n2294,dia[5],open_n2295}),
    .wea(wea[0]),
    .doa({open_n2310,open_n2311,open_n2312,open_n2313,open_n2314,open_n2315,open_n2316,open_n2317,inst_doa_i1_005}));
  // address_offset=8192;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_006 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2343,open_n2344,addra[13]}),
    .dia({open_n2348,open_n2349,open_n2350,open_n2351,open_n2352,open_n2353,open_n2354,dia[6],open_n2355}),
    .wea(wea[0]),
    .doa({open_n2370,open_n2371,open_n2372,open_n2373,open_n2374,open_n2375,open_n2376,open_n2377,inst_doa_i1_006}));
  // address_offset=8192;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_007 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2403,open_n2404,addra[13]}),
    .dia({open_n2408,open_n2409,open_n2410,open_n2411,open_n2412,open_n2413,open_n2414,dia[7],open_n2415}),
    .wea(wea[0]),
    .doa({open_n2430,open_n2431,open_n2432,open_n2433,open_n2434,open_n2435,open_n2436,open_n2437,inst_doa_i1_007}));
  // address_offset=8192;data_offset=8;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_008 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2463,open_n2464,addra[13]}),
    .dia({open_n2468,open_n2469,open_n2470,open_n2471,open_n2472,open_n2473,open_n2474,dia[8],open_n2475}),
    .wea(wea[1]),
    .doa({open_n2490,open_n2491,open_n2492,open_n2493,open_n2494,open_n2495,open_n2496,open_n2497,inst_doa_i1_008}));
  // address_offset=8192;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_009 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2523,open_n2524,addra[13]}),
    .dia({open_n2528,open_n2529,open_n2530,open_n2531,open_n2532,open_n2533,open_n2534,dia[9],open_n2535}),
    .wea(wea[1]),
    .doa({open_n2550,open_n2551,open_n2552,open_n2553,open_n2554,open_n2555,open_n2556,open_n2557,inst_doa_i1_009}));
  // address_offset=8192;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_010 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2583,open_n2584,addra[13]}),
    .dia({open_n2588,open_n2589,open_n2590,open_n2591,open_n2592,open_n2593,open_n2594,dia[10],open_n2595}),
    .wea(wea[1]),
    .doa({open_n2610,open_n2611,open_n2612,open_n2613,open_n2614,open_n2615,open_n2616,open_n2617,inst_doa_i1_010}));
  // address_offset=8192;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_011 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2643,open_n2644,addra[13]}),
    .dia({open_n2648,open_n2649,open_n2650,open_n2651,open_n2652,open_n2653,open_n2654,dia[11],open_n2655}),
    .wea(wea[1]),
    .doa({open_n2670,open_n2671,open_n2672,open_n2673,open_n2674,open_n2675,open_n2676,open_n2677,inst_doa_i1_011}));
  // address_offset=8192;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_012 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2703,open_n2704,addra[13]}),
    .dia({open_n2708,open_n2709,open_n2710,open_n2711,open_n2712,open_n2713,open_n2714,dia[12],open_n2715}),
    .wea(wea[1]),
    .doa({open_n2730,open_n2731,open_n2732,open_n2733,open_n2734,open_n2735,open_n2736,open_n2737,inst_doa_i1_012}));
  // address_offset=8192;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_013 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2763,open_n2764,addra[13]}),
    .dia({open_n2768,open_n2769,open_n2770,open_n2771,open_n2772,open_n2773,open_n2774,dia[13],open_n2775}),
    .wea(wea[1]),
    .doa({open_n2790,open_n2791,open_n2792,open_n2793,open_n2794,open_n2795,open_n2796,open_n2797,inst_doa_i1_013}));
  // address_offset=8192;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_014 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2823,open_n2824,addra[13]}),
    .dia({open_n2828,open_n2829,open_n2830,open_n2831,open_n2832,open_n2833,open_n2834,dia[14],open_n2835}),
    .wea(wea[1]),
    .doa({open_n2850,open_n2851,open_n2852,open_n2853,open_n2854,open_n2855,open_n2856,open_n2857,inst_doa_i1_014}));
  // address_offset=8192;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_015 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2883,open_n2884,addra[13]}),
    .dia({open_n2888,open_n2889,open_n2890,open_n2891,open_n2892,open_n2893,open_n2894,dia[15],open_n2895}),
    .wea(wea[1]),
    .doa({open_n2910,open_n2911,open_n2912,open_n2913,open_n2914,open_n2915,open_n2916,open_n2917,inst_doa_i1_015}));
  // address_offset=8192;data_offset=16;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_016 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n2943,open_n2944,addra[13]}),
    .dia({open_n2948,open_n2949,open_n2950,open_n2951,open_n2952,open_n2953,open_n2954,dia[16],open_n2955}),
    .wea(wea[2]),
    .doa({open_n2970,open_n2971,open_n2972,open_n2973,open_n2974,open_n2975,open_n2976,open_n2977,inst_doa_i1_016}));
  // address_offset=8192;data_offset=17;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_017 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3003,open_n3004,addra[13]}),
    .dia({open_n3008,open_n3009,open_n3010,open_n3011,open_n3012,open_n3013,open_n3014,dia[17],open_n3015}),
    .wea(wea[2]),
    .doa({open_n3030,open_n3031,open_n3032,open_n3033,open_n3034,open_n3035,open_n3036,open_n3037,inst_doa_i1_017}));
  // address_offset=8192;data_offset=18;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_018 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3063,open_n3064,addra[13]}),
    .dia({open_n3068,open_n3069,open_n3070,open_n3071,open_n3072,open_n3073,open_n3074,dia[18],open_n3075}),
    .wea(wea[2]),
    .doa({open_n3090,open_n3091,open_n3092,open_n3093,open_n3094,open_n3095,open_n3096,open_n3097,inst_doa_i1_018}));
  // address_offset=8192;data_offset=19;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_019 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3123,open_n3124,addra[13]}),
    .dia({open_n3128,open_n3129,open_n3130,open_n3131,open_n3132,open_n3133,open_n3134,dia[19],open_n3135}),
    .wea(wea[2]),
    .doa({open_n3150,open_n3151,open_n3152,open_n3153,open_n3154,open_n3155,open_n3156,open_n3157,inst_doa_i1_019}));
  // address_offset=8192;data_offset=20;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_020 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3183,open_n3184,addra[13]}),
    .dia({open_n3188,open_n3189,open_n3190,open_n3191,open_n3192,open_n3193,open_n3194,dia[20],open_n3195}),
    .wea(wea[2]),
    .doa({open_n3210,open_n3211,open_n3212,open_n3213,open_n3214,open_n3215,open_n3216,open_n3217,inst_doa_i1_020}));
  // address_offset=8192;data_offset=21;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_021 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3243,open_n3244,addra[13]}),
    .dia({open_n3248,open_n3249,open_n3250,open_n3251,open_n3252,open_n3253,open_n3254,dia[21],open_n3255}),
    .wea(wea[2]),
    .doa({open_n3270,open_n3271,open_n3272,open_n3273,open_n3274,open_n3275,open_n3276,open_n3277,inst_doa_i1_021}));
  // address_offset=8192;data_offset=22;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_022 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3303,open_n3304,addra[13]}),
    .dia({open_n3308,open_n3309,open_n3310,open_n3311,open_n3312,open_n3313,open_n3314,dia[22],open_n3315}),
    .wea(wea[2]),
    .doa({open_n3330,open_n3331,open_n3332,open_n3333,open_n3334,open_n3335,open_n3336,open_n3337,inst_doa_i1_022}));
  // address_offset=8192;data_offset=23;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_023 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3363,open_n3364,addra[13]}),
    .dia({open_n3368,open_n3369,open_n3370,open_n3371,open_n3372,open_n3373,open_n3374,dia[23],open_n3375}),
    .wea(wea[2]),
    .doa({open_n3390,open_n3391,open_n3392,open_n3393,open_n3394,open_n3395,open_n3396,open_n3397,inst_doa_i1_023}));
  // address_offset=8192;data_offset=24;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_024 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3423,open_n3424,addra[13]}),
    .dia({open_n3428,open_n3429,open_n3430,open_n3431,open_n3432,open_n3433,open_n3434,dia[24],open_n3435}),
    .wea(wea[3]),
    .doa({open_n3450,open_n3451,open_n3452,open_n3453,open_n3454,open_n3455,open_n3456,open_n3457,inst_doa_i1_024}));
  // address_offset=8192;data_offset=25;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_025 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3483,open_n3484,addra[13]}),
    .dia({open_n3488,open_n3489,open_n3490,open_n3491,open_n3492,open_n3493,open_n3494,dia[25],open_n3495}),
    .wea(wea[3]),
    .doa({open_n3510,open_n3511,open_n3512,open_n3513,open_n3514,open_n3515,open_n3516,open_n3517,inst_doa_i1_025}));
  // address_offset=8192;data_offset=26;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_026 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3543,open_n3544,addra[13]}),
    .dia({open_n3548,open_n3549,open_n3550,open_n3551,open_n3552,open_n3553,open_n3554,dia[26],open_n3555}),
    .wea(wea[3]),
    .doa({open_n3570,open_n3571,open_n3572,open_n3573,open_n3574,open_n3575,open_n3576,open_n3577,inst_doa_i1_026}));
  // address_offset=8192;data_offset=27;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_027 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3603,open_n3604,addra[13]}),
    .dia({open_n3608,open_n3609,open_n3610,open_n3611,open_n3612,open_n3613,open_n3614,dia[27],open_n3615}),
    .wea(wea[3]),
    .doa({open_n3630,open_n3631,open_n3632,open_n3633,open_n3634,open_n3635,open_n3636,open_n3637,inst_doa_i1_027}));
  // address_offset=8192;data_offset=28;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_028 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3663,open_n3664,addra[13]}),
    .dia({open_n3668,open_n3669,open_n3670,open_n3671,open_n3672,open_n3673,open_n3674,dia[28],open_n3675}),
    .wea(wea[3]),
    .doa({open_n3690,open_n3691,open_n3692,open_n3693,open_n3694,open_n3695,open_n3696,open_n3697,inst_doa_i1_028}));
  // address_offset=8192;data_offset=29;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_029 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3723,open_n3724,addra[13]}),
    .dia({open_n3728,open_n3729,open_n3730,open_n3731,open_n3732,open_n3733,open_n3734,dia[29],open_n3735}),
    .wea(wea[3]),
    .doa({open_n3750,open_n3751,open_n3752,open_n3753,open_n3754,open_n3755,open_n3756,open_n3757,inst_doa_i1_029}));
  // address_offset=8192;data_offset=30;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_030 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3783,open_n3784,addra[13]}),
    .dia({open_n3788,open_n3789,open_n3790,open_n3791,open_n3792,open_n3793,open_n3794,dia[30],open_n3795}),
    .wea(wea[3]),
    .doa({open_n3810,open_n3811,open_n3812,open_n3813,open_n3814,open_n3815,open_n3816,open_n3817,inst_doa_i1_030}));
  // address_offset=8192;data_offset=31;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;working_numbyte=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_16384x32_sub_008192_031 (
    .addra(addra[12:0]),
    .clka(clka),
    .csa({open_n3843,open_n3844,addra[13]}),
    .dia({open_n3848,open_n3849,open_n3850,open_n3851,open_n3852,open_n3853,open_n3854,dia[31],open_n3855}),
    .wea(wea[3]),
    .doa({open_n3870,open_n3871,open_n3872,open_n3873,open_n3874,open_n3875,open_n3876,open_n3877,inst_doa_i1_031}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_0  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i1_010),
    .sel(addra_piped),
    .o(doa[10]));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_0  (
    .i0(inst_doa_i0_011),
    .i1(inst_doa_i1_011),
    .sel(addra_piped),
    .o(doa[11]));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_0  (
    .i0(inst_doa_i0_012),
    .i1(inst_doa_i1_012),
    .sel(addra_piped),
    .o(doa[12]));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_0  (
    .i0(inst_doa_i0_013),
    .i1(inst_doa_i1_013),
    .sel(addra_piped),
    .o(doa[13]));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_0  (
    .i0(inst_doa_i0_014),
    .i1(inst_doa_i1_014),
    .sel(addra_piped),
    .o(doa[14]));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_0  (
    .i0(inst_doa_i0_015),
    .i1(inst_doa_i1_015),
    .sel(addra_piped),
    .o(doa[15]));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_0  (
    .i0(inst_doa_i0_016),
    .i1(inst_doa_i1_016),
    .sel(addra_piped),
    .o(doa[16]));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_0  (
    .i0(inst_doa_i0_017),
    .i1(inst_doa_i1_017),
    .sel(addra_piped),
    .o(doa[17]));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_0  (
    .i0(inst_doa_i0_018),
    .i1(inst_doa_i1_018),
    .sel(addra_piped),
    .o(doa[18]));
  AL_MUX \inst_doa_mux_b19/al_mux_b0_0_0  (
    .i0(inst_doa_i0_019),
    .i1(inst_doa_i1_019),
    .sel(addra_piped),
    .o(doa[19]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b20/al_mux_b0_0_0  (
    .i0(inst_doa_i0_020),
    .i1(inst_doa_i1_020),
    .sel(addra_piped),
    .o(doa[20]));
  AL_MUX \inst_doa_mux_b21/al_mux_b0_0_0  (
    .i0(inst_doa_i0_021),
    .i1(inst_doa_i1_021),
    .sel(addra_piped),
    .o(doa[21]));
  AL_MUX \inst_doa_mux_b22/al_mux_b0_0_0  (
    .i0(inst_doa_i0_022),
    .i1(inst_doa_i1_022),
    .sel(addra_piped),
    .o(doa[22]));
  AL_MUX \inst_doa_mux_b23/al_mux_b0_0_0  (
    .i0(inst_doa_i0_023),
    .i1(inst_doa_i1_023),
    .sel(addra_piped),
    .o(doa[23]));
  AL_MUX \inst_doa_mux_b24/al_mux_b0_0_0  (
    .i0(inst_doa_i0_024),
    .i1(inst_doa_i1_024),
    .sel(addra_piped),
    .o(doa[24]));
  AL_MUX \inst_doa_mux_b25/al_mux_b0_0_0  (
    .i0(inst_doa_i0_025),
    .i1(inst_doa_i1_025),
    .sel(addra_piped),
    .o(doa[25]));
  AL_MUX \inst_doa_mux_b26/al_mux_b0_0_0  (
    .i0(inst_doa_i0_026),
    .i1(inst_doa_i1_026),
    .sel(addra_piped),
    .o(doa[26]));
  AL_MUX \inst_doa_mux_b27/al_mux_b0_0_0  (
    .i0(inst_doa_i0_027),
    .i1(inst_doa_i1_027),
    .sel(addra_piped),
    .o(doa[27]));
  AL_MUX \inst_doa_mux_b28/al_mux_b0_0_0  (
    .i0(inst_doa_i0_028),
    .i1(inst_doa_i1_028),
    .sel(addra_piped),
    .o(doa[28]));
  AL_MUX \inst_doa_mux_b29/al_mux_b0_0_0  (
    .i0(inst_doa_i0_029),
    .i1(inst_doa_i1_029),
    .sel(addra_piped),
    .o(doa[29]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b30/al_mux_b0_0_0  (
    .i0(inst_doa_i0_030),
    .i1(inst_doa_i1_030),
    .sel(addra_piped),
    .o(doa[30]));
  AL_MUX \inst_doa_mux_b31/al_mux_b0_0_0  (
    .i0(inst_doa_i0_031),
    .i1(inst_doa_i1_031),
    .sel(addra_piped),
    .o(doa[31]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped),
    .o(doa[7]));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_0  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i1_008),
    .sel(addra_piped),
    .o(doa[8]));
  AL_MUX \inst_doa_mux_b9/al_mux_b0_0_0  (
    .i0(inst_doa_i0_009),
    .i1(inst_doa_i1_009),
    .sel(addra_piped),
    .o(doa[9]));

endmodule 

module AL_DFF_X
  (
  ar,
  as,
  clk,
  d,
  en,
  sr,
  ss,
  q
  );

  input ar;
  input as;
  input clk;
  input d;
  input en;
  input sr;
  input ss;
  output q;

  wire enout;
  wire srout;
  wire ssout;

  AL_MUX u_en (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset (
    .i0(ssout),
    .i1(1'b0),
    .sel(sr),
    .o(srout));
  AL_DFF u_seq (
    .clk(clk),
    .d(srout),
    .reset(ar),
    .set(as),
    .q(q));
  AL_MUX u_set (
    .i0(enout),
    .i1(1'b1),
    .sel(ss),
    .o(ssout));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  // synthesis translate_off
  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end
  // synthesis translate_on

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

